* NGSPICE file created from cbx_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

.subckt cbx_1__0_ bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
+ bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
+ bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_ bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
+ bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_ bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
+ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9]
+ chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13]
+ chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] pReset
+ prog_clk top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_ top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
+ top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_ vccd1 vssd1 vssd1_uq0 vccd1_uq0
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_501_ prog_clk mem_top_ipin_4.DFFR_3_.Q _037_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_4.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_432_ _070_ vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__inv_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_294_ mem_top_ipin_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__inv_2
X_363_ net14 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output56_A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__304__A mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__506__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_346_ net2 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_0_.out sky130_fd_sc_hd__inv_2
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_415_ _069_ vssd1 vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__inv_2
XFILLER_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_277_ mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _135_ sky130_fd_sc_hd__inv_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_630__95 vssd1 vssd1 vccd1 vccd1 net95 _630__95/LO sky130_fd_sc_hd__conb_1
XANTENNA__529__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_329_ mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _091_ sky130_fd_sc_hd__inv_2
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_680_ mux_top_ipin_0.INVTX1_5_.out _174_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__402__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__312__A mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_663_ mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out _157_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XANTENNA_input18_A chanx_left_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_594_ mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out _088_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output86_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__307__A mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 chanx_left_out[12] sky130_fd_sc_hd__buf_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 chanx_right_out[8] sky130_fd_sc_hd__buf_2
X_646_ mux_bottom_ipin_0.INVTX1_2_.out _140_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_577_ net6 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_500_ prog_clk mem_top_ipin_4.DFFR_4_.Q _036_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_4.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_431_ _070_ vssd1 vssd1 vccd1 vccd1 _035_ sky130_fd_sc_hd__inv_2
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_362_ net33 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_293_ mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _125_ sky130_fd_sc_hd__inv_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__410__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_629_ mux_top_ipin_2.INVTX1_7_.out _123_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_output49_A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__320__A mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_414_ _066_ vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__buf_4
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_276_ mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _136_ sky130_fd_sc_hd__inv_2
X_345_ net30 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XANTENNA__405__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__497__D mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__315__A mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_606__93 vssd1 vssd1 vccd1 vccd1 net93 _606__93/LO sky130_fd_sc_hd__conb_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_259_ mem_top_ipin_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _156_ sky130_fd_sc_hd__inv_2
X_328_ mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__inv_2
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__519__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_662_ mux_bottom_ipin_0.INVTX1_0_.out _156_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_593_ mux_bottom_ipin_1.INVTX1_7_.out _087_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__413__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output79_A net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__323__A mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__491__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 chanx_right_out[9] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 chanx_right_out[16] sky130_fd_sc_hd__buf_2
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 chanx_left_out[6] sky130_fd_sc_hd__buf_2
XFILLER_56_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_645_ mux_top_ipin_2.INVTX1_3_.out _139_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_input30_A chanx_right_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__408__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_576_ net7 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_430_ _070_ vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__inv_2
X_292_ mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _126_ sky130_fd_sc_hd__inv_2
XFILLER_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__228__A mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_361_ net20 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_628_ mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out _122_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_559_ net24 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_413_ _068_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__inv_2
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_275_ mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _142_ sky130_fd_sc_hd__inv_2
XFILLER_41_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_344_ mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net89 sky130_fd_sc_hd__inv_2
XANTENNA__421__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__331__A mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__241__A mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_258_ mem_top_ipin_4.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _153_ sky130_fd_sc_hd__inv_2
XANTENNA__416__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_327_ mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _095_ sky130_fd_sc_hd__inv_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_661_ mux_bottom_ipin_0.INVTX1_3_.out _155_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_592_ net92 _086_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_
+ sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 chanx_left_out[7] sky130_fd_sc_hd__buf_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 chanx_right_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_575_ net8 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_644_ mux_bottom_ipin_0.INVTX1_5_.out _138_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_input23_A chanx_right_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__509__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__424__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_291_ mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _131_ sky130_fd_sc_hd__inv_2
X_360_ net39 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__481__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_627_ mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out _121_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XANTENNA__419__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_558_ net25 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
X_489_ prog_clk mem_top_ipin_2.DFFR_3_.Q _025_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_2.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__329__A mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__239__A mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_412_ _068_ vssd1 vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__inv_2
XFILLER_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_274_ mem_top_ipin_3.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _134_ sky130_fd_sc_hd__inv_2
X_343_ net11 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_326_ mem_bottom_ipin_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _085_ sky130_fd_sc_hd__inv_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_257_ mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _161_ sky130_fd_sc_hd__inv_2
XANTENNA__432__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__342__A net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__252__A mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_309_ mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _103_ sky130_fd_sc_hd__inv_2
XANTENNA__427__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__337__A mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_591_ mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out _085_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_660_ mux_bottom_ipin_1.INVTX1_6_.out _154_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__247__A mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 chanx_right_out[18] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_574_ net9 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A chanx_left_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_643_ mux_bottom_ipin_0.INVTX1_4_.out _137_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__440__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__615__A mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A chanx_left_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__500__D mem_top_ipin_4.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__350__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_290_ mem_top_ipin_2.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__inv_2
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__260__A mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_488_ prog_clk mem_top_ipin_2.DFFR_4_.Q _024_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_2.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_626_ mux_top_ipin_0.INVTX1_2_.out _120_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_557_ net26 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XANTENNA__435__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_642__96 vssd1 vssd1 vccd1 vccd1 net96 _642__96/LO sky130_fd_sc_hd__conb_1
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__345__A net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_411_ _068_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__inv_2
XFILLER_37_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_342_ net24 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_273_ mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _139_ sky130_fd_sc_hd__inv_2
XANTENNA__255__A mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_609_ mux_bottom_ipin_2.INVTX1_3_.out _103_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__471__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_325_ mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__inv_2
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_256_ mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _162_ sky130_fd_sc_hd__inv_2
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__494__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__443__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_308_ mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__inv_2
X_239_ mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _178_ sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__353__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_590_ mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out _084_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__438__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__348__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 chanx_left_out[9] sky130_fd_sc_hd__buf_2
X_642_ net96 _136_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__258__A mem_top_ipin_4.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_573_ net10 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__541__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_625_ mux_top_ipin_1.INVTX1_3_.out _119_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_487_ prog_clk mem_top_ipin_0.DFFR_5_.Q _023_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_1.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_556_ net27 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_618__94 vssd1 vssd1 vccd1 vccd1 net94 _618__94/LO sky130_fd_sc_hd__conb_1
XANTENNA__361__A net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ _068_ vssd1 vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__inv_2
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_341_ mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__inv_2
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_272_ mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _140_ sky130_fd_sc_hd__inv_2
XANTENNA__271__A mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__446__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_608_ mux_top_ipin_0.INVTX1_5_.out _102_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__266__A mem_top_ipin_4.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_324_ mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _087_ sky130_fd_sc_hd__inv_2
X_255_ mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _167_ sky130_fd_sc_hd__inv_2
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chanx_right_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_307_ mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _108_ sky130_fd_sc_hd__inv_2
X_238_ mem_top_ipin_6.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _170_ sky130_fd_sc_hd__inv_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__484__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__364__A net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_641_ mux_bottom_ipin_0.INVTX1_7_.out _135_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_572_ net11 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__509__D mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input21_A chanx_right_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_624_ mux_top_ipin_1.INVTX1_6_.out _118_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_555_ net28 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_2
X_486_ prog_clk mem_top_ipin_1.DFFR_0_.Q _022_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_1.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__522__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_340_ mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _074_ sky130_fd_sc_hd__inv_2
X_271_ mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _144_ sky130_fd_sc_hd__inv_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_607_ mux_top_ipin_0.INVTX1_4_.out _101_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_469_ prog_clk net1 _005_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_0.DFFR_0_.Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__372__A mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__522__D mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__547__A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_254_ mem_top_ipin_5.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _157_ sky130_fd_sc_hd__inv_2
X_323_ mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__inv_2
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__277__A mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_306_ mem_top_ipin_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__inv_2
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_237_ mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _175_ sky130_fd_sc_hd__inv_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__560__A net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__380__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_640_ mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out _134_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
X_571_ net21 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__555__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__525__D mem_bottom_ipin_2.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__375__A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__474__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A chanx_left_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_623_ mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out _117_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
X_485_ prog_clk mem_top_ipin_1.DFFR_1_.Q _021_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_1.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__285__A mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_554_ net29 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output82_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__497__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A chanx_left_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_270_ mem_top_ipin_3.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _141_ sky130_fd_sc_hd__inv_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_468_ prog_clk mem_bottom_ipin_0.DFFR_0_.Q _004_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_0.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_606_ net93 _100_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_399_ _067_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__inv_2
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__653__A mux_bottom_ipin_1.INVTX1_7_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__512__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ mem_bottom_ipin_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__inv_2
X_253_ mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _159_ sky130_fd_sc_hd__inv_2
XANTENNA__563__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__383__A net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_305_ mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__inv_2
XFILLER_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__293__A mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_236_ mem_top_ipin_6.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _176_ sky130_fd_sc_hd__inv_2
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__288__A mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_219_ mem_bottom_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _200_ sky130_fd_sc_hd__inv_2
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_56_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_570_ net31 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__571__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_654__97 vssd1 vssd1 vccd1 vccd1 net97 _654__97/LO sky130_fd_sc_hd__conb_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_699_ mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out _193_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out sky130_fd_sc_hd__ebufn_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_622_ mux_top_ipin_1.INVTX1_2_.out _116_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_484_ prog_clk mem_top_ipin_1.DFFR_2_.Q _020_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_1.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_553_ net30 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__296__A mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_605_ mux_top_ipin_0.INVTX1_7_.out _099_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_398_ _067_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__inv_2
X_467_ prog_clk mem_bottom_ipin_0.DFFR_1_.Q _003_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_0.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__464__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_252_ mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _160_ sky130_fd_sc_hd__inv_2
X_321_ mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _089_ sky130_fd_sc_hd__inv_2
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__487__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_519_ prog_clk mem_top_ipin_7.DFFR_3_.Q _055_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_7.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__574__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_235_ mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _180_ sky130_fd_sc_hd__inv_2
X_304_ mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__inv_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__502__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__394__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input37_A chanx_right_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_218_ mem_bottom_ipin_2.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _193_ sky130_fd_sc_hd__inv_2
XANTENNA__525__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__389__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_698_ mux_top_ipin_0.INVTX1_2_.out _192_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_621_ mux_top_ipin_0.INVTX1_3_.out _115_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_552_ net2 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_483_ prog_clk mem_top_ipin_1.DFFR_3_.Q _019_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_1.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_604_ mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out _098_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XANTENNA__577__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_466_ prog_clk mem_bottom_ipin_0.DFFR_2_.Q _002_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_0.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_397_ _067_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__inv_2
XFILLER_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__397__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _166_ sky130_fd_sc_hd__inv_2
X_320_ mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__inv_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_518_ prog_clk mem_top_ipin_7.DFFR_4_.Q _054_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__dfrtp_4
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_449_ _072_ vssd1 vssd1 vccd1 vccd1 _051_ sky130_fd_sc_hd__inv_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_303_ mem_top_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__inv_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_234_ mem_top_ipin_6.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _177_ sky130_fd_sc_hd__inv_2
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__477__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_217_ mem_bottom_ipin_2.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _194_ sky130_fd_sc_hd__inv_2
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_697_ mux_top_ipin_0.INVTX1_5_.out _191_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__515__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_620_ mux_top_ipin_1.INVTX1_5_.out _114_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_551_ net12 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_482_ prog_clk mem_top_ipin_1.DFFR_4_.Q _018_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_1.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_603_ mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out _097_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_465_ prog_clk mem_bottom_ipin_0.DFFR_3_.Q _001_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_0.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__593__A mux_bottom_ipin_1.INVTX1_7_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A chanx_left_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_396_ _067_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__inv_2
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output80_A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A chanx_left_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_250_ mem_top_ipin_5.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _158_ sky130_fd_sc_hd__inv_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_517_ prog_clk mem_top_ipin_5.DFFR_5_.Q _053_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_6.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_448_ _072_ vssd1 vssd1 vccd1 vccd1 _050_ sky130_fd_sc_hd__inv_2
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__473__D mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_379_ mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net46 sky130_fd_sc_hd__inv_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_302_ mem_top_ipin_1.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _109_ sky130_fd_sc_hd__inv_2
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_233_ mem_top_ipin_7.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _185_ sky130_fd_sc_hd__inv_2
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__468__D mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_216_ mem_bottom_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _197_ sky130_fd_sc_hd__inv_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_696_ mux_top_ipin_1.INVTX1_6_.out _190_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__467__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_481_ prog_clk mem_bottom_ipin_2.DFFR_5_.Q _017_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_0.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_550_ net13 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__520__RESET_B _056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__476__D mem_top_ipin_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_679_ mux_top_ipin_0.INVTX1_4_.out _173_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_602_ mux_bottom_ipin_0.INVTX1_0_.out _096_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_464_ prog_clk mem_bottom_ipin_0.DFFR_4_.Q _000_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_0.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_395_ _067_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__inv_2
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__505__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__528__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_447_ net40 vssd1 vssd1 vccd1 vccd1 _072_ sky130_fd_sc_hd__buf_4
X_516_ prog_clk mem_top_ipin_6.DFFR_0_.Q _052_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_6.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_378_ mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net45 sky130_fd_sc_hd__inv_2
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_301_ mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__inv_2
XFILLER_42_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_232_ mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _186_ sky130_fd_sc_hd__inv_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__484__D mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_666__98 vssd1 vssd1 vccd1 vccd1 net98 _666__98/LO sky130_fd_sc_hd__conb_1
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_215_ mem_bottom_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _198_ sky130_fd_sc_hd__inv_2
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__479__D mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input35_A chanx_right_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_695_ mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out _189_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_480_ prog_clk mem_top_ipin_0.DFFR_0_.Q _016_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_0.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__400__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__492__D mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_678_ net99 _172_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_601_ mux_bottom_ipin_1.INVTX1_3_.out _095_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_463_ _066_ vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__inv_2
X_394_ _067_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__inv_2
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__305__A mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_515_ prog_clk mem_top_ipin_6.DFFR_1_.Q _051_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_6.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_446_ _071_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__inv_2
X_377_ mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net44 sky130_fd_sc_hd__inv_2
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_300_ mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__inv_2
X_231_ mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _191_ sky130_fd_sc_hd__inv_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_429_ _070_ vssd1 vssd1 vccd1 vccd1 _033_ sky130_fd_sc_hd__inv_2
Xinput1 ccff_head vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__518__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_214_ mem_bottom_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _201_ sky130_fd_sc_hd__inv_2
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__313__A mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__223__A mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A chanx_right_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__490__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_694_ mux_top_ipin_0.INVTX1_4_.out _188_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__308__A mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_677_ mux_top_ipin_0.INVTX1_7_.out _171_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_600_ mux_bottom_ipin_1.INVTX1_6_.out _094_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_462_ _066_ vssd1 vssd1 vccd1 vccd1 _064_ sky130_fd_sc_hd__inv_2
X_393_ _067_ vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__inv_2
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output59_A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__411__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__321__A mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__231__A mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A chanx_left_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_514_ prog_clk mem_top_ipin_6.DFFR_2_.Q _050_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_6.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_445_ _071_ vssd1 vssd1 vccd1 vccd1 _048_ sky130_fd_sc_hd__inv_2
XANTENNA__406__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_376_ net29 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__498__D mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__316__A mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A chanx_left_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_230_ mem_top_ipin_7.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _181_ sky130_fd_sc_hd__inv_2
XANTENNA__226__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_428_ _070_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__inv_2
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_359_ net8 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 chanx_left_in[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_213_ mem_bottom_ipin_2.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _199_ sky130_fd_sc_hd__inv_2
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_693_ mux_top_ipin_0.INVTX1_3_.out _187_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__508__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__324__A mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__640__TE_B _134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input40_A pReset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_676_ mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out _170_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__409__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__319__A mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__480__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_461_ _066_ vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__inv_2
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_392_ _066_ vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__buf_4
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_659_ mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out _153_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_444_ _071_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__inv_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_513_ prog_clk mem_top_ipin_6.DFFR_3_.Q _049_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_6.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_375_ net16 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__422__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_358_ mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net41 sky130_fd_sc_hd__inv_2
X_427_ _070_ vssd1 vssd1 vccd1 vccd1 _031_ sky130_fd_sc_hd__inv_2
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__417__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_289_ mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput3 chanx_left_in[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__327__A mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__237__A mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_692_ mux_top_ipin_1.INVTX1_5_.out _186_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__430__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__340__A mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A chanx_right_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_675_ mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out _169_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__335__A mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_391_ net40 vssd1 vssd1 vccd1 vccd1 _066_ sky130_fd_sc_hd__clkbuf_4
X_460_ _066_ vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__inv_2
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__245__A mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_658_ mux_bottom_ipin_0.INVTX1_2_.out _152_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_589_ mux_bottom_ipin_0.INVTX1_6_.out _083_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_512_ prog_clk mem_top_ipin_6.DFFR_4_.Q _048_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_6.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_443_ _071_ vssd1 vssd1 vccd1 vccd1 _046_ sky130_fd_sc_hd__inv_2
XFILLER_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_374_ net35 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__470__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output64_A net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_678__99 vssd1 vssd1 vccd1 vccd1 net99 _678__99/LO sky130_fd_sc_hd__conb_1
XANTENNA__613__A mux_top_ipin_0.INVTX1_3_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__493__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_426_ _070_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__inv_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_357_ net25 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XANTENNA__433__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_288_ mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _124_ sky130_fd_sc_hd__inv_2
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 chanx_left_in[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__343__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__253__A mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__428__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_409_ _068_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__inv_2
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__338__A mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_691_ mux_top_ipin_1.INVTX1_4_.out _185_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__248__A mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput40 pReset vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__621__A mux_top_ipin_0.INVTX1_3_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_674_ mux_bottom_ipin_1.INVTX1_2_.out _168_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_input26_A chanx_right_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__441__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__501__D mem_top_ipin_4.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_390_ net23 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_657_ mux_bottom_ipin_0.INVTX1_1_.out _151_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_588_ mux_bottom_ipin_0.INVTX1_3_.out _082_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_511_ prog_clk mem_top_ipin_4.DFFR_5_.Q _047_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_5.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_700__101 vssd1 vssd1 vccd1 vccd1 net101 _700__101/LO sky130_fd_sc_hd__conb_1
X_442_ _071_ vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__inv_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_373_ net10 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.INVTX1_6_.out sky130_fd_sc_hd__clkinv_2
XANTENNA__256__A mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output57_A net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_425_ _066_ vssd1 vssd1 vccd1 vccd1 _070_ sky130_fd_sc_hd__buf_4
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_287_ mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _130_ sky130_fd_sc_hd__inv_2
X_356_ net12 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 chanx_left_in[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_408_ _068_ vssd1 vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__inv_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__444__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_339_ mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__inv_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__483__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_690_ net100 _184_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
X_583__91 vssd1 vssd1 vccd1 vccd1 net91 _583__91/LO sky130_fd_sc_hd__conb_1
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__264__A mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__439__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 chanx_right_in[18] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__349__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_673_ mux_bottom_ipin_1.INVTX1_5_.out _167_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_input19_A chanx_left_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output87_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__521__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__542__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_587_ mux_bottom_ipin_0.INVTX1_0_.out _081_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_656_ mux_bottom_ipin_1.INVTX1_5_.out _150_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__362__A net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_441_ _071_ vssd1 vssd1 vccd1 vccd1 _044_ sky130_fd_sc_hd__inv_2
X_510_ prog_clk mem_top_ipin_5.DFFR_0_.Q _046_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_5.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_372_ mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net43 sky130_fd_sc_hd__inv_2
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__272__A mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_639_ mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out _133_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_8_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_424_ _069_ vssd1 vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__inv_2
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_286_ mem_top_ipin_2.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__inv_2
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_355_ net31 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 chanx_left_in[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__550__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_407_ _068_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__inv_2
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_338_ mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _076_ sky130_fd_sc_hd__inv_2
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_269_ mem_top_ipin_4.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _149_ sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_592__92 vssd1 vssd1 vccd1 vccd1 net92 _592__92/LO sky130_fd_sc_hd__conb_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__520__D mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__370__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__280__A mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 chanx_left_in[9] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 chanx_right_in[1] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_2
XANTENNA__365__A mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__515__D mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_672_ mux_top_ipin_5.INVTX1_6_.out _166_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__275__A mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__473__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__496__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input31_A chanx_right_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_655_ mux_bottom_ipin_1.INVTX1_4_.out _149_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_586_ mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out _080_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_440_ _071_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__inv_2
X_371_ net28 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__553__A net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__511__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_707_ mux_bottom_ipin_1.INVTX1_2_.out _201_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_638_ mux_top_ipin_1.INVTX1_2_.out _132_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_569_ net32 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__373__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__548__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_423_ _069_ vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__inv_2
X_354_ net18 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__283__A mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_285_ mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _127_ sky130_fd_sc_hd__inv_2
Xinput7 chanx_left_in[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__368__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_406_ _068_ vssd1 vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__inv_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_337_ mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__inv_2
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_268_ mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _150_ sky130_fd_sc_hd__inv_2
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 chanx_right_in[0] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 chanx_left_in[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_2
Xinput32 chanx_right_in[2] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__381__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_671_ mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out _165_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__556__A net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__291__A mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__376__A net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_654_ net97 _148_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input24_A chanx_right_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_585_ mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out _079_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_370_ net15 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_706_ mux_bottom_ipin_2.INVTX1_3_.out _200_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_637_ mux_top_ipin_2.INVTX1_3_.out _131_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_499_ prog_clk mem_top_ipin_2.DFFR_5_.Q _035_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_3.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_568_ net33 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__486__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_422_ _069_ vssd1 vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__inv_2
XANTENNA__564__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_353_ net37 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
X_284_ mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _128_ sky130_fd_sc_hd__inv_2
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 chanx_left_in[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__384__A mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__501__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__559__A net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_405_ _068_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__inv_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_267_ mem_top_ipin_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _155_ sky130_fd_sc_hd__inv_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_336_ mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _078_ sky130_fd_sc_hd__inv_2
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__524__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__289__A mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_319_ mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__inv_2
Xinput33 chanx_right_in[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 chanx_right_in[10] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_left_in[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_670_ mux_bottom_ipin_1.INVTX1_4_.out _164_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__572__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A chanx_left_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_653_ mux_bottom_ipin_1.INVTX1_7_.out _147_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_584_ mux_bottom_ipin_0.INVTX1_7_.out _078_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__387__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A chanx_left_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_705_ mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out _199_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out sky130_fd_sc_hd__ebufn_2
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__297__A mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_636_ mux_top_ipin_2.INVTX1_6_.out _130_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_567_ net34 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
X_498_ prog_clk mem_top_ipin_3.DFFR_0_.Q _034_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_3.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_421_ _069_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__inv_2
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_283_ mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _132_ sky130_fd_sc_hd__inv_2
X_352_ net6 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 chanx_left_in[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_2
X_619_ mux_top_ipin_1.INVTX1_4_.out _113_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_404_ _068_ vssd1 vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__inv_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_266_ mem_top_ipin_4.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _145_ sky130_fd_sc_hd__inv_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_335_ mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__inv_2
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__476__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__395__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__499__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_249_ mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _163_ sky130_fd_sc_hd__inv_2
Xinput34 chanx_right_in[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dlymetal6s2s_1
X_318_ mem_bottom_ipin_1.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _093_ sky130_fd_sc_hd__inv_2
Xinput12 chanx_left_in[1] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 chanx_right_in[11] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__514__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_652_ mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_2_out _146_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_583_ net91 _077_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_704_ mux_bottom_ipin_2.INVTX1_2_.out _198_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__578__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_635_ mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out _129_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
X_566_ net35 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_497_ prog_clk mem_top_ipin_3.DFFR_1_.Q _033_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_3.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__398__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_420_ _069_ vssd1 vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__inv_2
X_351_ mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net90 sky130_fd_sc_hd__inv_2
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_282_ mem_top_ipin_2.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _129_ sky130_fd_sc_hd__inv_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_618_ net94 _112_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_549_ net14 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_403_ _066_ vssd1 vssd1 vccd1 vccd1 _068_ sky130_fd_sc_hd__buf_4
X_334_ mem_bottom_ipin_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__inv_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_265_ mem_top_ipin_4.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _147_ sky130_fd_sc_hd__inv_2
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 chanx_left_in[2] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__dlymetal6s2s_1
X_317_ mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__inv_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput35 chanx_right_in[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__dlymetal6s2s_1
X_248_ mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _164_ sky130_fd_sc_hd__inv_2
Xinput24 chanx_right_in[12] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__466__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__466__D mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__489__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_651_ mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_1_out _145_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_4.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_582_ mux_bottom_ipin_0.INVTX1_4_.out _076_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__504__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_634_ mux_top_ipin_2.INVTX1_2_.out _128_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_703_ mux_bottom_ipin_1.INVTX1_3_.out _197_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input22_A chanx_right_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_496_ prog_clk mem_top_ipin_3.DFFR_2_.Q _032_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_3.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_565_ net36 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__527__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_350_ net5 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_281_ mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _137_ sky130_fd_sc_hd__inv_2
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_617_ mux_top_ipin_1.INVTX1_7_.out _111_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_479_ prog_clk mem_top_ipin_0.DFFR_1_.Q _015_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_0.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__474__D mem_bottom_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_548_ net15 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_402_ _067_ vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__inv_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_264_ mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _148_ sky130_fd_sc_hd__inv_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_333_ mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _082_ sky130_fd_sc_hd__inv_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__469__D net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 chanx_left_in[3] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
Xinput36 chanx_right_in[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_316_ mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__inv_2
X_247_ mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _168_ sky130_fd_sc_hd__inv_2
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput25 chanx_right_in[13] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__300__A mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_650_ mux_top_ipin_2.INVTX1_2_.out _144_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
X_581_ mux_bottom_ipin_0.INVTX1_5_.out _075_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input15_A chanx_left_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_702_ mux_bottom_ipin_2.INVTX1_5_.out _196_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_633_ mux_top_ipin_1.INVTX1_3_.out _127_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_495_ prog_clk mem_top_ipin_3.DFFR_3_.Q _031_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_3.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_564_ net37 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__479__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A chanx_left_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_280_ mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _138_ sky130_fd_sc_hd__inv_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_616_ mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_2_out _110_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_547_ net16 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_1
XANTENNA__490__D mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_478_ prog_clk mem_top_ipin_0.DFFR_2_.Q _014_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_0.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_401_ _067_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__inv_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_332_ mem_bottom_ipin_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _080_ sky130_fd_sc_hd__inv_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_263_ mem_top_ipin_4.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _154_ sky130_fd_sc_hd__inv_2
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__517__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__485__D mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__213__A mem_bottom_ipin_2.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_246_ mem_top_ipin_5.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _165_ sky130_fd_sc_hd__inv_2
Xinput15 chanx_left_in[4] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_2
X_315_ mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__inv_2
Xinput37 chanx_right_in[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_2
Xinput26 chanx_right_in[14] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_229_ mem_top_ipin_7.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _183_ sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_580_ mux_bottom_ipin_0.INVTX1_1_.out _074_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__401__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__311__A mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_632_ mux_bottom_ipin_2.INVTX1_5_.out _126_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_701_ mux_bottom_ipin_2.INVTX1_4_.out _195_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_563_ net38 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
X_494_ prog_clk mem_top_ipin_3.DFFR_4_.Q _030_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_3.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_615_ mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out _109_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_546_ net17 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
X_477_ prog_clk mem_top_ipin_0.DFFR_3_.Q _013_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_0.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__469__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_331_ mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__inv_2
X_400_ _067_ vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__inv_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_262_ mem_top_ipin_4.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _146_ sky130_fd_sc_hd__inv_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_529_ prog_clk mem_bottom_ipin_1.DFFR_5_.Q _065_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_2.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_314_ mem_top_ipin_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__inv_2
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 chanx_left_in[5] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_2
XANTENNA__404__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_245_ mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _173_ sky130_fd_sc_hd__inv_2
Xinput38 chanx_right_in[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput27 chanx_right_in[15] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__496__D mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__314__A mem_top_ipin_0.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__507__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__224__A mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input38_A chanx_right_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_228_ mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _184_ sky130_fd_sc_hd__inv_2
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__309__A mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_700_ net101 _194_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_493_ prog_clk mem_top_ipin_1.DFFR_5_.Q _029_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_2.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_631_ mux_bottom_ipin_2.INVTX1_4_.out _125_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_562_ net39 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__412__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__232__A mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A chanx_left_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_476_ prog_clk mem_top_ipin_0.DFFR_4_.Q _012_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_0.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_614_ mux_bottom_ipin_2.INVTX1_2_.out _108_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__407__A _068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_545_ net18 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__317__A mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__227__A mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_330_ mem_bottom_ipin_0.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__inv_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_261_ mem_top_ipin_4.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _151_ sky130_fd_sc_hd__inv_2
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_459_ _066_ vssd1 vssd1 vccd1 vccd1 _061_ sky130_fd_sc_hd__inv_2
X_528_ prog_clk mem_bottom_ipin_2.DFFR_0_.Q _064_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_2.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_244_ mem_top_ipin_6.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _174_ sky130_fd_sc_hd__inv_2
X_313_ mem_top_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__inv_2
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 chanx_left_in[6] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_2
Xinput28 chanx_right_in[16] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_2
Xinput39 chanx_right_in[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__420__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_227_ mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _190_ sky130_fd_sc_hd__inv_2
XANTENNA__415__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__325__A mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__235__A mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_630_ net95 _124_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_492_ prog_clk mem_top_ipin_2.DFFR_0_.Q _028_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_2.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_561_ net22 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A chanx_left_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_613_ mux_top_ipin_0.INVTX1_3_.out _107_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_475_ prog_clk mem_bottom_ipin_0.DFFR_5_.Q _011_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_1.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_544_ net19 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_2
XANTENNA__423__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__492__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__333__A mem_bottom_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_A chanx_left_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_260_ mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _152_ sky130_fd_sc_hd__inv_2
XFILLER_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__243__A mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_527_ prog_clk mem_bottom_ipin_2.DFFR_1_.Q _063_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_2.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__418__A _069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_458_ _066_ vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__inv_2
X_389_ net13 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__328__A mem_bottom_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 chanx_left_in[7] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__dlymetal6s2s_1
X_312_ mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__inv_2
X_243_ mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _179_ sky130_fd_sc_hd__inv_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 chanx_right_in[17] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_226_ net49 vssd1 vssd1 vccd1 vccd1 _182_ sky130_fd_sc_hd__inv_2
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__431__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__341__A mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__251__A mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__426__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__336__A mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_560_ net23 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_491_ prog_clk mem_top_ipin_2.DFFR_1_.Q _027_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_2.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_689_ mux_top_ipin_1.INVTX1_7_.out _183_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_612_ mux_top_ipin_0.INVTX1_6_.out _106_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_543_ net20 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_2
X_474_ prog_clk mem_bottom_ipin_1.DFFR_0_.Q _010_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_1.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output74_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_526_ prog_clk mem_bottom_ipin_2.DFFR_2_.Q _062_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_2.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_457_ _072_ vssd1 vssd1 vccd1 vccd1 _059_ sky130_fd_sc_hd__inv_2
X_388_ net32 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XANTENNA__434__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__344__A mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__482__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 chanx_left_in[8] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_2
X_311_ mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__inv_2
X_242_ mem_top_ipin_6.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _169_ sky130_fd_sc_hd__inv_2
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__429__A _070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_509_ prog_clk mem_top_ipin_5.DFFR_1_.Q _045_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_5.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__339__A mem_bottom_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__249__A mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_225_ mem_top_ipin_7.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _187_ sky130_fd_sc_hd__inv_2
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__520__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input36_A chanx_right_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__442__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__352__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__502__D mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_490_ prog_clk mem_top_ipin_2.DFFR_2_.Q _026_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_2.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__437__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_688_ mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_2_out _182_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__347__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_542_ net3 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_611_ mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out _105_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_473_ prog_clk mem_bottom_ipin_1.DFFR_1_.Q _009_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_1.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__257__A mem_top_ipin_5.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_525_ prog_clk mem_bottom_ipin_2.DFFR_3_.Q _061_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_2.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_456_ _072_ vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__inv_2
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_387_ net4 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_2.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__360__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__510__D mem_top_ipin_5.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_310_ mem_top_ipin_0.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__inv_2
XFILLER_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_241_ mem_top_ipin_6.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _171_ sky130_fd_sc_hd__inv_2
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_508_ prog_clk mem_top_ipin_5.DFFR_2_.Q _044_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_5.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_439_ _071_ vssd1 vssd1 vccd1 vccd1 _042_ sky130_fd_sc_hd__inv_2
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__445__A _071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__355__A net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_224_ mem_top_ipin_7.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _188_ sky130_fd_sc_hd__inv_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__525__RESET_B _061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__472__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input29_A chanx_right_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__495__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__543__A net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_687_ mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_1_out _181_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__510__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__363__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_610_ mux_top_ipin_0.INVTX1_2_.out _104_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_472_ prog_clk mem_bottom_ipin_1.DFFR_2_.Q _008_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_1.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_541_ net4 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__273__A mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__508__D mem_top_ipin_5.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__268__A mem_top_ipin_4.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input11_A chanx_left_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_386_ mux_bottom_ipin_2.mux_2level_tapbuf_basis_input3_mem3_2_out vssd1 vssd1 vccd1
+ vccd1 net88 sky130_fd_sc_hd__inv_2
X_524_ prog_clk mem_bottom_ipin_2.DFFR_4_.Q _060_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_2.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_455_ _072_ vssd1 vssd1 vccd1 vccd1 _057_ sky130_fd_sc_hd__inv_2
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_
+ sky130_fd_sc_hd__buf_2
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input3_A chanx_left_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_240_ mem_top_ipin_6.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _172_ sky130_fd_sc_hd__inv_2
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_507_ prog_clk mem_top_ipin_5.DFFR_3_.Q _043_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_5.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
X_438_ _071_ vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__inv_2
X_369_ net34 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__371__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_223_ mem_top_ipin_7.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _192_ sky130_fd_sc_hd__inv_2
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__546__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__281__A mem_top_ipin_3.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__366__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__516__D mem_top_ipin_6.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__276__A mem_top_ipin_3.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_686_ mux_bottom_ipin_2.INVTX1_2_.out _180_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_471_ prog_clk mem_bottom_ipin_1.DFFR_3_.Q _007_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_1.DFFR_4_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__485__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__554__A net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_669_ mux_bottom_ipin_1.INVTX1_3_.out _163_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_523_ prog_clk mem_top_ipin_6.DFFR_5_.Q _059_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_7.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__549__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_454_ _072_ vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__inv_2
XANTENNA__284__A mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_385_ mux_top_ipin_7.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net48 sky130_fd_sc_hd__inv_2
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__500__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__523__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__279__A mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_506_ prog_clk mem_top_ipin_5.DFFR_4_.Q _042_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_5.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_299_ mem_top_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__inv_2
X_368_ net3 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.INVTX1_4_.out sky130_fd_sc_hd__inv_2
X_437_ _071_ vssd1 vssd1 vccd1 vccd1 _040_ sky130_fd_sc_hd__inv_2
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_222_ mem_top_ipin_7.DFFR_3_.Q vssd1 vssd1 vccd1 vccd1 _189_ sky130_fd_sc_hd__inv_2
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__562__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__557__A net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__292__A mem_top_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__377__A mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input34_A chanx_right_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__287__A mem_top_ipin_2.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_685_ mux_top_ipin_5.INVTX1_5_.out _179_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_470_ prog_clk mem_bottom_ipin_1.DFFR_4_.Q _006_ vssd1 vssd1 vccd1 vccd1 mem_bottom_ipin_1.DFFR_5_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__570__A net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_599_ mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out _093_ vssd1 vssd1
+ vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
X_668_ mux_top_ipin_5.INVTX1_5_.out _162_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__390__A net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_453_ _072_ vssd1 vssd1 vccd1 vccd1 _055_ sky130_fd_sc_hd__inv_2
X_522_ prog_clk mem_top_ipin_7.DFFR_0_.Q _058_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_7.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__565__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_384_ mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net47 sky130_fd_sc_hd__inv_2
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 chanx_right_out[10] sky130_fd_sc_hd__buf_2
XFILLER_63_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 chanx_right_out[3] sky130_fd_sc_hd__buf_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__475__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_436_ net40 vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__buf_4
X_505_ prog_clk mem_top_ipin_3.DFFR_5_.Q _041_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_4.DFFR_0_.Q
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_298_ mem_top_ipin_1.DFFR_5_.Q vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__inv_2
XANTENNA__498__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_367_ net22 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_221_ mem_bottom_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _195_ sky130_fd_sc_hd__inv_2
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_419_ _069_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__inv_2
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__513__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__573__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__393__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__568__A net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_684_ mux_top_ipin_0.INVTX1_6_.out _178_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_input27_A chanx_right_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_667_ mux_top_ipin_5.INVTX1_4_.out _161_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
X_598_ mux_bottom_ipin_1.INVTX1_4_.out _092_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__671__A mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_0_out vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_452_ _072_ vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__inv_2
X_521_ prog_clk mem_top_ipin_7.DFFR_1_.Q _057_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_7.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_383_ net26 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 chanx_right_out[11] sky130_fd_sc_hd__buf_2
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 chanx_right_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_output58_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__576__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_366_ net9 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_1.INVTX1_6_.out sky130_fd_sc_hd__inv_2
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_504_ prog_clk mem_top_ipin_4.DFFR_0_.Q _040_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_4.DFFR_1_.Q
+ sky130_fd_sc_hd__dfrtp_2
X_435_ _070_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__inv_2
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_297_ mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__inv_2
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__396__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ccff_head vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_220_ mem_bottom_ipin_2.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _196_ sky130_fd_sc_hd__inv_2
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_418_ _069_ vssd1 vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__inv_2
X_349_ net36 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_3_.out sky130_fd_sc_hd__inv_2
XANTENNA__465__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__488__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_690__100 vssd1 vssd1 vccd1 vccd1 net100 _690__100/LO sky130_fd_sc_hd__conb_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_683_ mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out _177_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__503__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__526__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_666_ net98 _160_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_597_ mux_bottom_ipin_1.INVTX1_5_.out _091_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__399__A _067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_520_ prog_clk mem_top_ipin_7.DFFR_2_.Q _056_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_7.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_451_ _072_ vssd1 vssd1 vccd1 vccd1 _053_ sky130_fd_sc_hd__inv_2
X_382_ net19 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.INVTX1_4_.out sky130_fd_sc_hd__inv_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_649_ mux_bottom_ipin_0.INVTX1_3_.out _143_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_1_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_503_ prog_clk mem_top_ipin_4.DFFR_1_.Q _039_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_4.DFFR_2_.Q
+ sky130_fd_sc_hd__dfrtp_4
X_365_ mux_top_ipin_1.mux_2level_tapbuf_basis_input3_mem3_3_out vssd1 vssd1 vccd1
+ vccd1 net42 sky130_fd_sc_hd__inv_2
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_296_ mem_top_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__inv_2
X_434_ _070_ vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__inv_2
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_417_ _069_ vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__inv_2
X_348_ net17 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_2_.out sky130_fd_sc_hd__inv_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__472__D mem_bottom_ipin_1.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_279_ mem_top_ipin_3.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _143_ sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__467__D mem_bottom_ipin_0.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_682_ mux_top_ipin_5.INVTX1_4_.out _176_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__478__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_665_ mux_top_ipin_5.INVTX1_7_.out _159_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_input32_A chanx_right_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_596_ mux_bottom_ipin_0.INVTX1_1_.out _090_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__480__D mem_top_ipin_0.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_450_ _072_ vssd1 vssd1 vccd1 vccd1 _052_ sky130_fd_sc_hd__inv_2
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_381_ net38 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.INVTX1_5_.out sky130_fd_sc_hd__inv_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 chanx_right_out[6] sky130_fd_sc_hd__buf_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_648_ mux_bottom_ipin_0.INVTX1_6_.out _142_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_2_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_579_ mux_bottom_ipin_0.INVTX1_2_.out _073_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__516__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_502_ prog_clk mem_top_ipin_4.DFFR_2_.Q _038_ vssd1 vssd1 vccd1 vccd1 mem_top_ipin_4.DFFR_3_.Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_433_ _070_ vssd1 vssd1 vccd1 vccd1 _037_ sky130_fd_sc_hd__inv_2
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_295_ mem_top_ipin_1.DFFR_0_.Q vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__inv_2
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_364_ net27 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_0.INVTX1_7_.out sky130_fd_sc_hd__inv_2
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__693__A mux_top_ipin_0.INVTX1_3_.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_416_ _069_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__inv_2
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_278_ mem_top_ipin_3.DFFR_4_.Q vssd1 vssd1 vccd1 vccd1 _133_ sky130_fd_sc_hd__inv_2
X_347_ net21 vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_0.INVTX1_1_.out sky130_fd_sc_hd__inv_2
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__301__A mem_top_ipin_1.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_681_ mux_bottom_ipin_2.INVTX1_3_.out _175_ vssd1 vssd1 vccd1 vccd1 mux_top_ipin_6.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__478__D mem_top_ipin_0.DFFR_2_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_664_ mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_2_out _158_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_5.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_2
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_595_ mux_bottom_ipin_1.INVTX1_2_.out _089_ vssd1 vssd1 vccd1 vccd1 mux_bottom_ipin_1.mux_2level_tapbuf_basis_input3_mem3_0_out
+ sky130_fd_sc_hd__ebufn_2
XFILLER_28_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input25_A chanx_right_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_380_ net7 vssd1 vssd1 vccd1 vccd1 mux_top_ipin_5.INVTX1_6_.out sky130_fd_sc_hd__clkinv_2
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__buf_2
XFILLER_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__468__CLK prog_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_647_ mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_0_out _141_ vssd1 vssd1
+ vccd1 vccd1 mux_top_ipin_3.mux_2level_tapbuf_basis_input3_mem3_3_out sky130_fd_sc_hd__ebufn_4
X_578_ net5 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__491__D mem_top_ipin_2.DFFR_1_.Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

