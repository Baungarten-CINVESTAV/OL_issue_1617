magic
tech sky130A
magscale 1 2
timestamp 1674174269
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 38824 37732
<< metal2 >>
rect 18 39200 74 39800
rect 1950 39200 2006 39800
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18694 39200 18750 39800
rect 20626 39200 20682 39800
rect 21914 39200 21970 39800
rect 23846 39200 23902 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 35438 39200 35494 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 4526 200 4582 800
rect 6458 200 6514 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 23202 200 23258 800
rect 25134 200 25190 800
rect 26422 200 26478 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36726 200 36782 800
rect 38014 200 38070 800
<< obsm2 >>
rect 130 39144 1894 39250
rect 2062 39144 3826 39250
rect 3994 39144 5114 39250
rect 5282 39144 7046 39250
rect 7214 39144 8334 39250
rect 8502 39144 10266 39250
rect 10434 39144 12198 39250
rect 12366 39144 13486 39250
rect 13654 39144 15418 39250
rect 15586 39144 16706 39250
rect 16874 39144 18638 39250
rect 18806 39144 20570 39250
rect 20738 39144 21858 39250
rect 22026 39144 23790 39250
rect 23958 39144 25078 39250
rect 25246 39144 27010 39250
rect 27178 39144 28942 39250
rect 29110 39144 30230 39250
rect 30398 39144 32162 39250
rect 32330 39144 33450 39250
rect 33618 39144 35382 39250
rect 35550 39144 37314 39250
rect 37482 39144 38602 39250
rect 20 856 38712 39144
rect 130 144 1250 856
rect 1418 144 3182 856
rect 3350 144 4470 856
rect 4638 144 6402 856
rect 6570 144 8334 856
rect 8502 144 9622 856
rect 9790 144 11554 856
rect 11722 144 12842 856
rect 13010 144 14774 856
rect 14942 144 16706 856
rect 16874 144 17994 856
rect 18162 144 19926 856
rect 20094 144 21214 856
rect 21382 144 23146 856
rect 23314 144 25078 856
rect 25246 144 26366 856
rect 26534 144 28298 856
rect 28466 144 29586 856
rect 29754 144 31518 856
rect 31686 144 33450 856
rect 33618 144 34738 856
rect 34906 144 36670 856
rect 36838 144 37958 856
rect 38126 144 38712 856
rect 20 31 38712 144
<< metal3 >>
rect 200 38768 800 38888
rect 39200 38768 39800 38888
rect 39200 37408 39800 37528
rect 200 36728 800 36848
rect 200 35368 800 35488
rect 39200 35368 39800 35488
rect 200 33328 800 33448
rect 39200 33328 39800 33448
rect 39200 31968 39800 32088
rect 200 31288 800 31408
rect 200 29928 800 30048
rect 39200 29928 39800 30048
rect 39200 28568 39800 28688
rect 200 27888 800 28008
rect 200 26528 800 26648
rect 39200 26528 39800 26648
rect 200 24488 800 24608
rect 39200 24488 39800 24608
rect 39200 23128 39800 23248
rect 200 22448 800 22568
rect 200 21088 800 21208
rect 39200 21088 39800 21208
rect 39200 19728 39800 19848
rect 200 19048 800 19168
rect 200 17688 800 17808
rect 39200 17688 39800 17808
rect 200 15648 800 15768
rect 39200 15648 39800 15768
rect 39200 14288 39800 14408
rect 200 13608 800 13728
rect 200 12248 800 12368
rect 39200 12248 39800 12368
rect 39200 10888 39800 11008
rect 200 10208 800 10328
rect 200 8848 800 8968
rect 39200 8848 39800 8968
rect 200 6808 800 6928
rect 39200 6808 39800 6928
rect 39200 5448 39800 5568
rect 200 4768 800 4888
rect 200 3408 800 3528
rect 39200 3408 39800 3528
rect 39200 2048 39800 2168
rect 200 1368 800 1488
rect 39200 8 39800 128
<< obsm3 >>
rect 880 38688 39120 38861
rect 800 37608 39200 38688
rect 800 37328 39120 37608
rect 800 36928 39200 37328
rect 880 36648 39200 36928
rect 800 35568 39200 36648
rect 880 35288 39120 35568
rect 800 33528 39200 35288
rect 880 33248 39120 33528
rect 800 32168 39200 33248
rect 800 31888 39120 32168
rect 800 31488 39200 31888
rect 880 31208 39200 31488
rect 800 30128 39200 31208
rect 880 29848 39120 30128
rect 800 28768 39200 29848
rect 800 28488 39120 28768
rect 800 28088 39200 28488
rect 880 27808 39200 28088
rect 800 26728 39200 27808
rect 880 26448 39120 26728
rect 800 24688 39200 26448
rect 880 24408 39120 24688
rect 800 23328 39200 24408
rect 800 23048 39120 23328
rect 800 22648 39200 23048
rect 880 22368 39200 22648
rect 800 21288 39200 22368
rect 880 21008 39120 21288
rect 800 19928 39200 21008
rect 800 19648 39120 19928
rect 800 19248 39200 19648
rect 880 18968 39200 19248
rect 800 17888 39200 18968
rect 880 17608 39120 17888
rect 800 15848 39200 17608
rect 880 15568 39120 15848
rect 800 14488 39200 15568
rect 800 14208 39120 14488
rect 800 13808 39200 14208
rect 880 13528 39200 13808
rect 800 12448 39200 13528
rect 880 12168 39120 12448
rect 800 11088 39200 12168
rect 800 10808 39120 11088
rect 800 10408 39200 10808
rect 880 10128 39200 10408
rect 800 9048 39200 10128
rect 880 8768 39120 9048
rect 800 7008 39200 8768
rect 880 6728 39120 7008
rect 800 5648 39200 6728
rect 800 5368 39120 5648
rect 800 4968 39200 5368
rect 880 4688 39200 4968
rect 800 3608 39200 4688
rect 880 3328 39120 3608
rect 800 2248 39200 3328
rect 800 1968 39120 2248
rect 800 1568 39200 1968
rect 880 1288 39200 1568
rect 800 208 39200 1288
rect 800 35 39120 208
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 1715 2619 4128 37229
rect 4608 2619 19445 37229
<< labels >>
rlabel metal3 s 39200 26528 39800 26648 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 39200 37408 39800 37528 6 ccff_tail
port 2 nsew signal output
rlabel metal2 s 38658 39200 38714 39800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 38014 200 38070 800 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal3 s 39200 19728 39800 19848 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal2 s 35438 39200 35494 39800 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal3 s 200 3408 800 3528 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal3 s 200 19048 800 19168 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 31574 200 31630 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal3 s 39200 12248 39800 12368 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal2 s 20626 39200 20682 39800 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal2 s 1950 39200 2006 39800 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal2 s 36726 200 36782 800 6 chany_bottom_in[1]
port 13 nsew signal input
rlabel metal2 s 14830 200 14886 800 6 chany_bottom_in[2]
port 14 nsew signal input
rlabel metal3 s 200 4768 800 4888 6 chany_bottom_in[3]
port 15 nsew signal input
rlabel metal3 s 39200 33328 39800 33448 6 chany_bottom_in[4]
port 16 nsew signal input
rlabel metal2 s 13542 39200 13598 39800 6 chany_bottom_in[5]
port 17 nsew signal input
rlabel metal3 s 200 38768 800 38888 6 chany_bottom_in[6]
port 18 nsew signal input
rlabel metal3 s 200 33328 800 33448 6 chany_bottom_in[7]
port 19 nsew signal input
rlabel metal3 s 39200 5448 39800 5568 6 chany_bottom_in[8]
port 20 nsew signal input
rlabel metal2 s 9678 200 9734 800 6 chany_bottom_in[9]
port 21 nsew signal input
rlabel metal3 s 39200 28568 39800 28688 6 chany_bottom_out[0]
port 22 nsew signal output
rlabel metal2 s 16762 39200 16818 39800 6 chany_bottom_out[10]
port 23 nsew signal output
rlabel metal3 s 39200 31968 39800 32088 6 chany_bottom_out[11]
port 24 nsew signal output
rlabel metal3 s 200 27888 800 28008 6 chany_bottom_out[12]
port 25 nsew signal output
rlabel metal2 s 23846 39200 23902 39800 6 chany_bottom_out[13]
port 26 nsew signal output
rlabel metal3 s 39200 29928 39800 30048 6 chany_bottom_out[14]
port 27 nsew signal output
rlabel metal2 s 18 39200 74 39800 6 chany_bottom_out[15]
port 28 nsew signal output
rlabel metal3 s 200 1368 800 1488 6 chany_bottom_out[16]
port 29 nsew signal output
rlabel metal3 s 200 15648 800 15768 6 chany_bottom_out[17]
port 30 nsew signal output
rlabel metal2 s 8390 200 8446 800 6 chany_bottom_out[18]
port 31 nsew signal output
rlabel metal2 s 18694 39200 18750 39800 6 chany_bottom_out[1]
port 32 nsew signal output
rlabel metal2 s 15474 39200 15530 39800 6 chany_bottom_out[2]
port 33 nsew signal output
rlabel metal3 s 39200 8848 39800 8968 6 chany_bottom_out[3]
port 34 nsew signal output
rlabel metal2 s 25134 39200 25190 39800 6 chany_bottom_out[4]
port 35 nsew signal output
rlabel metal2 s 27066 39200 27122 39800 6 chany_bottom_out[5]
port 36 nsew signal output
rlabel metal2 s 34794 200 34850 800 6 chany_bottom_out[6]
port 37 nsew signal output
rlabel metal3 s 200 17688 800 17808 6 chany_bottom_out[7]
port 38 nsew signal output
rlabel metal3 s 39200 35368 39800 35488 6 chany_bottom_out[8]
port 39 nsew signal output
rlabel metal2 s 25134 200 25190 800 6 chany_bottom_out[9]
port 40 nsew signal output
rlabel metal3 s 200 21088 800 21208 6 chany_top_in[0]
port 41 nsew signal input
rlabel metal3 s 39200 2048 39800 2168 6 chany_top_in[10]
port 42 nsew signal input
rlabel metal3 s 39200 15648 39800 15768 6 chany_top_in[11]
port 43 nsew signal input
rlabel metal2 s 4526 200 4582 800 6 chany_top_in[12]
port 44 nsew signal input
rlabel metal3 s 200 13608 800 13728 6 chany_top_in[13]
port 45 nsew signal input
rlabel metal3 s 200 31288 800 31408 6 chany_top_in[14]
port 46 nsew signal input
rlabel metal2 s 28354 200 28410 800 6 chany_top_in[15]
port 47 nsew signal input
rlabel metal3 s 200 29928 800 30048 6 chany_top_in[16]
port 48 nsew signal input
rlabel metal2 s 7102 39200 7158 39800 6 chany_top_in[17]
port 49 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 chany_top_in[18]
port 50 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 chany_top_in[1]
port 51 nsew signal input
rlabel metal2 s 33506 200 33562 800 6 chany_top_in[2]
port 52 nsew signal input
rlabel metal3 s 39200 14288 39800 14408 6 chany_top_in[3]
port 53 nsew signal input
rlabel metal3 s 39200 6808 39800 6928 6 chany_top_in[4]
port 54 nsew signal input
rlabel metal3 s 200 6808 800 6928 6 chany_top_in[5]
port 55 nsew signal input
rlabel metal3 s 200 36728 800 36848 6 chany_top_in[6]
port 56 nsew signal input
rlabel metal3 s 39200 8 39800 128 6 chany_top_in[7]
port 57 nsew signal input
rlabel metal3 s 200 8848 800 8968 6 chany_top_in[8]
port 58 nsew signal input
rlabel metal3 s 39200 10888 39800 11008 6 chany_top_in[9]
port 59 nsew signal input
rlabel metal3 s 200 24488 800 24608 6 chany_top_out[0]
port 60 nsew signal output
rlabel metal2 s 29642 200 29698 800 6 chany_top_out[10]
port 61 nsew signal output
rlabel metal3 s 39200 24488 39800 24608 6 chany_top_out[11]
port 62 nsew signal output
rlabel metal2 s 10322 39200 10378 39800 6 chany_top_out[12]
port 63 nsew signal output
rlabel metal2 s 5170 39200 5226 39800 6 chany_top_out[13]
port 64 nsew signal output
rlabel metal2 s 18050 200 18106 800 6 chany_top_out[14]
port 65 nsew signal output
rlabel metal2 s 18 200 74 800 6 chany_top_out[15]
port 66 nsew signal output
rlabel metal2 s 23202 200 23258 800 6 chany_top_out[16]
port 67 nsew signal output
rlabel metal2 s 12254 39200 12310 39800 6 chany_top_out[17]
port 68 nsew signal output
rlabel metal2 s 21914 39200 21970 39800 6 chany_top_out[18]
port 69 nsew signal output
rlabel metal2 s 33506 39200 33562 39800 6 chany_top_out[1]
port 70 nsew signal output
rlabel metal3 s 200 26528 800 26648 6 chany_top_out[2]
port 71 nsew signal output
rlabel metal3 s 200 22448 800 22568 6 chany_top_out[3]
port 72 nsew signal output
rlabel metal2 s 1306 200 1362 800 6 chany_top_out[4]
port 73 nsew signal output
rlabel metal2 s 37370 39200 37426 39800 6 chany_top_out[5]
port 74 nsew signal output
rlabel metal2 s 28998 39200 29054 39800 6 chany_top_out[6]
port 75 nsew signal output
rlabel metal2 s 16762 200 16818 800 6 chany_top_out[7]
port 76 nsew signal output
rlabel metal3 s 39200 38768 39800 38888 6 chany_top_out[8]
port 77 nsew signal output
rlabel metal3 s 39200 3408 39800 3528 6 chany_top_out[9]
port 78 nsew signal output
rlabel metal3 s 200 10208 800 10328 6 left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
port 79 nsew signal output
rlabel metal3 s 39200 21088 39800 21208 6 left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
port 80 nsew signal output
rlabel metal2 s 6458 200 6514 800 6 left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
port 81 nsew signal output
rlabel metal2 s 12898 200 12954 800 6 left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
port 82 nsew signal output
rlabel metal2 s 19982 200 20038 800 6 left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_
port 83 nsew signal output
rlabel metal3 s 39200 23128 39800 23248 6 left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_
port 84 nsew signal output
rlabel metal2 s 21270 200 21326 800 6 left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_
port 85 nsew signal output
rlabel metal2 s 32218 39200 32274 39800 6 left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_
port 86 nsew signal output
rlabel metal2 s 30286 39200 30342 39800 6 pReset
port 87 nsew signal input
rlabel metal2 s 3882 39200 3938 39800 6 prog_clk
port 88 nsew signal input
rlabel metal2 s 8390 39200 8446 39800 6 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 89 nsew signal output
rlabel metal2 s 26422 200 26478 800 6 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 90 nsew signal output
rlabel metal3 s 200 12248 800 12368 6 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 91 nsew signal output
rlabel metal3 s 200 35368 800 35488 6 vccd1
port 92 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 92 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 92 nsew signal bidirectional
rlabel metal3 s 39200 17688 39800 17808 6 vssd1
port 93 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 93 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1885372
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/cby_0__1_/runs/23_01_19_18_23/results/signoff/cby_0__1_.magic.gds
string GDS_START 139574
<< end >>

