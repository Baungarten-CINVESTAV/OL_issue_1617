// This is the unpowered netlist.
module sb_0__4_ (bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
    bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_,
    bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_,
    ccff_head,
    ccff_tail,
    pReset,
    prog_clk,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_,
    right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_,
    right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
    right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
    vccd1,
    vssd1,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out);
 input bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
 input bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_;
 input bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_;
 input ccff_head;
 output ccff_tail;
 input pReset;
 input prog_clk;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_;
 input right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_;
 input right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
 input right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
 inout vccd1;
 inout vssd1;
 input [0:18] chanx_right_in;
 output [0:18] chanx_right_out;
 input [0:18] chany_bottom_in;
 output [0:18] chany_bottom_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire \mem_bottom_track_1.DFFR_0_.D ;
 wire \mem_bottom_track_1.DFFR_0_.Q ;
 wire \mem_bottom_track_1.DFFR_1_.Q ;
 wire \mem_bottom_track_11.DFFR_0_.D ;
 wire \mem_bottom_track_11.DFFR_0_.Q ;
 wire \mem_bottom_track_11.DFFR_1_.Q ;
 wire \mem_bottom_track_13.DFFR_0_.Q ;
 wire \mem_bottom_track_13.DFFR_1_.Q ;
 wire \mem_bottom_track_15.DFFR_0_.Q ;
 wire \mem_bottom_track_15.DFFR_1_.Q ;
 wire \mem_bottom_track_17.DFFR_0_.Q ;
 wire \mem_bottom_track_17.DFFR_1_.Q ;
 wire \mem_bottom_track_19.DFFR_0_.Q ;
 wire \mem_bottom_track_19.DFFR_1_.Q ;
 wire \mem_bottom_track_23.DFFR_0_.Q ;
 wire \mem_bottom_track_23.DFFR_1_.Q ;
 wire \mem_bottom_track_25.DFFR_0_.Q ;
 wire \mem_bottom_track_25.DFFR_1_.Q ;
 wire \mem_bottom_track_27.DFFR_0_.Q ;
 wire \mem_bottom_track_27.DFFR_1_.Q ;
 wire \mem_bottom_track_29.DFFR_0_.Q ;
 wire \mem_bottom_track_29.DFFR_1_.Q ;
 wire \mem_bottom_track_3.DFFR_0_.Q ;
 wire \mem_bottom_track_3.DFFR_1_.Q ;
 wire \mem_bottom_track_31.DFFR_0_.Q ;
 wire \mem_bottom_track_31.DFFR_1_.Q ;
 wire \mem_bottom_track_33.DFFR_0_.Q ;
 wire \mem_bottom_track_33.DFFR_1_.Q ;
 wire \mem_bottom_track_35.DFFR_0_.Q ;
 wire \mem_bottom_track_35.DFFR_1_.Q ;
 wire \mem_bottom_track_37.DFFR_0_.Q ;
 wire \mem_bottom_track_5.DFFR_0_.Q ;
 wire \mem_bottom_track_5.DFFR_1_.Q ;
 wire \mem_bottom_track_7.DFFR_0_.Q ;
 wire \mem_bottom_track_7.DFFR_1_.Q ;
 wire \mem_bottom_track_9.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_0_.Q ;
 wire \mem_right_track_0.DFFR_1_.Q ;
 wire \mem_right_track_10.DFFR_0_.D ;
 wire \mem_right_track_10.DFFR_0_.Q ;
 wire \mem_right_track_10.DFFR_1_.Q ;
 wire \mem_right_track_12.DFFR_0_.Q ;
 wire \mem_right_track_12.DFFR_1_.Q ;
 wire \mem_right_track_14.DFFR_0_.Q ;
 wire \mem_right_track_14.DFFR_1_.Q ;
 wire \mem_right_track_16.DFFR_0_.Q ;
 wire \mem_right_track_16.DFFR_1_.Q ;
 wire \mem_right_track_18.DFFR_0_.Q ;
 wire \mem_right_track_18.DFFR_1_.Q ;
 wire \mem_right_track_2.DFFR_0_.Q ;
 wire \mem_right_track_2.DFFR_1_.Q ;
 wire \mem_right_track_20.DFFR_0_.Q ;
 wire \mem_right_track_20.DFFR_1_.Q ;
 wire \mem_right_track_22.DFFR_0_.Q ;
 wire \mem_right_track_22.DFFR_1_.Q ;
 wire \mem_right_track_24.DFFR_0_.Q ;
 wire \mem_right_track_24.DFFR_1_.Q ;
 wire \mem_right_track_26.DFFR_0_.Q ;
 wire \mem_right_track_26.DFFR_1_.Q ;
 wire \mem_right_track_28.DFFR_0_.Q ;
 wire \mem_right_track_28.DFFR_1_.Q ;
 wire \mem_right_track_30.DFFR_0_.Q ;
 wire \mem_right_track_30.DFFR_1_.Q ;
 wire \mem_right_track_32.DFFR_0_.Q ;
 wire \mem_right_track_32.DFFR_1_.Q ;
 wire \mem_right_track_34.DFFR_0_.Q ;
 wire \mem_right_track_34.DFFR_1_.Q ;
 wire \mem_right_track_36.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_0_.Q ;
 wire \mem_right_track_4.DFFR_1_.Q ;
 wire \mem_right_track_6.DFFR_0_.Q ;
 wire \mem_right_track_6.DFFR_1_.Q ;
 wire \mem_right_track_8.DFFR_0_.Q ;
 wire \mux_bottom_track_1.INVTX1_0_.out ;
 wire \mux_bottom_track_1.INVTX1_1_.out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_1.out ;
 wire \mux_bottom_track_11.INVTX1_0_.out ;
 wire \mux_bottom_track_11.INVTX1_1_.out ;
 wire \mux_bottom_track_11.INVTX1_2_.out ;
 wire \mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_11.out ;
 wire \mux_bottom_track_13.INVTX1_0_.out ;
 wire \mux_bottom_track_13.INVTX1_2_.out ;
 wire \mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_13.out ;
 wire \mux_bottom_track_15.INVTX1_0_.out ;
 wire \mux_bottom_track_15.INVTX1_2_.out ;
 wire \mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_15.out ;
 wire \mux_bottom_track_17.INVTX1_0_.out ;
 wire \mux_bottom_track_17.INVTX1_2_.out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_17.out ;
 wire \mux_bottom_track_19.INVTX1_0_.out ;
 wire \mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_19.out ;
 wire \mux_bottom_track_23.INVTX1_0_.out ;
 wire \mux_bottom_track_23.INVTX1_1_.out ;
 wire \mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_23.out ;
 wire \mux_bottom_track_25.INVTX1_0_.out ;
 wire \mux_bottom_track_25.INVTX1_1_.out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_25.out ;
 wire \mux_bottom_track_27.INVTX1_0_.out ;
 wire \mux_bottom_track_27.INVTX1_1_.out ;
 wire \mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_27.out ;
 wire \mux_bottom_track_29.INVTX1_0_.out ;
 wire \mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_29.out ;
 wire \mux_bottom_track_3.INVTX1_0_.out ;
 wire \mux_bottom_track_3.INVTX1_1_.out ;
 wire \mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_3.out ;
 wire \mux_bottom_track_31.INVTX1_0_.out ;
 wire \mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_31.out ;
 wire \mux_bottom_track_33.INVTX1_0_.out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_33.out ;
 wire \mux_bottom_track_35.INVTX1_0_.out ;
 wire \mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_35.out ;
 wire \mux_bottom_track_37.INVTX1_0_.out ;
 wire \mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_37.out ;
 wire \mux_bottom_track_5.INVTX1_0_.out ;
 wire \mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_5.out ;
 wire \mux_bottom_track_7.INVTX1_0_.out ;
 wire \mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_7.out ;
 wire \mux_bottom_track_9.INVTX1_0_.out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_bottom_track_9.out ;
 wire \mux_right_track_0.INVTX1_0_.out ;
 wire \mux_right_track_0.INVTX1_1_.out ;
 wire \mux_right_track_0.INVTX1_2_.out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_0.out ;
 wire \mux_right_track_10.INVTX1_0_.out ;
 wire \mux_right_track_10.INVTX1_1_.out ;
 wire \mux_right_track_10.INVTX1_2_.out ;
 wire \mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_10.out ;
 wire \mux_right_track_12.INVTX1_1_.out ;
 wire \mux_right_track_12.INVTX1_2_.out ;
 wire \mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_12.out ;
 wire \mux_right_track_14.INVTX1_1_.out ;
 wire \mux_right_track_14.INVTX1_2_.out ;
 wire \mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_14.out ;
 wire \mux_right_track_16.INVTX1_1_.out ;
 wire \mux_right_track_16.INVTX1_2_.out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_16.out ;
 wire \mux_right_track_18.INVTX1_2_.out ;
 wire \mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_18.out ;
 wire \mux_right_track_2.INVTX1_1_.out ;
 wire \mux_right_track_2.INVTX1_2_.out ;
 wire \mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_2.out ;
 wire \mux_right_track_20.INVTX1_1_.out ;
 wire \mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_20.out ;
 wire \mux_right_track_22.INVTX1_1_.out ;
 wire \mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_22.out ;
 wire \mux_right_track_24.INVTX1_0_.out ;
 wire \mux_right_track_24.INVTX1_1_.out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_24.out ;
 wire \mux_right_track_26.INVTX1_0_.out ;
 wire \mux_right_track_26.INVTX1_1_.out ;
 wire \mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_26.out ;
 wire \mux_right_track_28.INVTX1_1_.out ;
 wire \mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_28.out ;
 wire \mux_right_track_30.INVTX1_1_.out ;
 wire \mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_30.out ;
 wire \mux_right_track_32.INVTX1_1_.out ;
 wire \mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_32.out ;
 wire \mux_right_track_34.INVTX1_1_.out ;
 wire \mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_34.out ;
 wire \mux_right_track_36.INVTX1_2_.out ;
 wire \mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_36.out ;
 wire \mux_right_track_4.INVTX1_2_.out ;
 wire \mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_4.out ;
 wire \mux_right_track_6.INVTX1_2_.out ;
 wire \mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_6.out ;
 wire \mux_right_track_8.INVTX1_2_.out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ;
 wire \mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ;
 wire \mux_right_track_8.out ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;

 sky130_fd_sc_hd__inv_2 _0404_ (.A(\mem_bottom_track_35.DFFR_1_.Q ),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _0405_ (.A(\mem_bottom_track_35.DFFR_0_.Q ),
    .Y(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0406_ (.A(\mem_bottom_track_35.DFFR_0_.Q ),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_1 _0407_ (.A(_0074_),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _0408_ (.A(\mem_bottom_track_35.DFFR_1_.Q ),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_1 _0409_ (.A(_0075_),
    .X(_0363_));
 sky130_fd_sc_hd__inv_2 _0410_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_2 _0411_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .Y(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0412_ (.A(\mem_bottom_track_33.DFFR_0_.Q ),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_1 _0413_ (.A(_0076_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _0414_ (.A(\mem_bottom_track_33.DFFR_1_.Q ),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_1 _0415_ (.A(_0077_),
    .X(_0359_));
 sky130_fd_sc_hd__inv_2 _0416_ (.A(\mem_bottom_track_31.DFFR_1_.Q ),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _0417_ (.A(\mem_bottom_track_31.DFFR_0_.Q ),
    .Y(_0358_));
 sky130_fd_sc_hd__clkbuf_1 _0418_ (.A(\mem_bottom_track_31.DFFR_0_.Q ),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _0419_ (.A(_0078_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0420_ (.A(\mem_bottom_track_31.DFFR_1_.Q ),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _0421_ (.A(_0079_),
    .X(_0355_));
 sky130_fd_sc_hd__inv_2 _0422_ (.A(\mem_bottom_track_29.DFFR_1_.Q ),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_2 _0423_ (.A(\mem_bottom_track_29.DFFR_0_.Q ),
    .Y(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0424_ (.A(\mem_bottom_track_29.DFFR_0_.Q ),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _0425_ (.A(_0080_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _0426_ (.A(\mem_bottom_track_29.DFFR_1_.Q ),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _0427_ (.A(_0081_),
    .X(_0351_));
 sky130_fd_sc_hd__inv_2 _0428_ (.A(\mem_bottom_track_27.DFFR_1_.Q ),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_2 _0429_ (.A(\mem_bottom_track_27.DFFR_0_.Q ),
    .Y(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _0430_ (.A(\mem_bottom_track_27.DFFR_0_.Q ),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _0431_ (.A(_0082_),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _0432_ (.A(\mem_bottom_track_27.DFFR_1_.Q ),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_1 _0433_ (.A(_0083_),
    .X(_0347_));
 sky130_fd_sc_hd__inv_2 _0434_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_2 _0435_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .Y(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _0436_ (.A(\mem_bottom_track_25.DFFR_0_.Q ),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_1 _0437_ (.A(_0084_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0438_ (.A(\mem_bottom_track_25.DFFR_1_.Q ),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0439_ (.A(_0085_),
    .X(_0343_));
 sky130_fd_sc_hd__inv_2 _0440_ (.A(\mem_bottom_track_23.DFFR_1_.Q ),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _0441_ (.A(\mem_bottom_track_23.DFFR_0_.Q ),
    .Y(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _0442_ (.A(\mem_bottom_track_23.DFFR_0_.Q ),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _0443_ (.A(_0086_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0444_ (.A(\mem_bottom_track_23.DFFR_1_.Q ),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_1 _0445_ (.A(_0087_),
    .X(_0339_));
 sky130_fd_sc_hd__inv_2 _0446_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _0447_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .Y(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _0448_ (.A(\mem_bottom_track_1.DFFR_0_.Q ),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0449_ (.A(_0088_),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_1 _0450_ (.A(\mem_bottom_track_1.DFFR_1_.Q ),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_1 _0451_ (.A(_0089_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_1 _0452_ (.A(\mem_right_track_0.DFFR_1_.Q ),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _0453_ (.A(_0090_),
    .X(_0177_));
 sky130_fd_sc_hd__inv_2 _0454_ (.A(\mem_right_track_34.DFFR_1_.Q ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_2 _0455_ (.A(\mem_right_track_34.DFFR_0_.Q ),
    .Y(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _0456_ (.A(\mem_right_track_34.DFFR_0_.Q ),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _0457_ (.A(_0091_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0458_ (.A(\mem_right_track_34.DFFR_1_.Q ),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _0459_ (.A(_0092_),
    .X(_0331_));
 sky130_fd_sc_hd__inv_2 _0460_ (.A(\mem_right_track_32.DFFR_1_.Q ),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_2 _0461_ (.A(\mem_right_track_32.DFFR_0_.Q ),
    .Y(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0462_ (.A(\mem_right_track_32.DFFR_0_.Q ),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_1 _0463_ (.A(_0093_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0464_ (.A(\mem_right_track_32.DFFR_1_.Q ),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _0465_ (.A(_0094_),
    .X(_0327_));
 sky130_fd_sc_hd__inv_2 _0466_ (.A(\mem_right_track_30.DFFR_1_.Q ),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_2 _0467_ (.A(\mem_right_track_30.DFFR_0_.Q ),
    .Y(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _0468_ (.A(\mem_right_track_30.DFFR_0_.Q ),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _0469_ (.A(_0095_),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _0470_ (.A(\mem_right_track_30.DFFR_1_.Q ),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _0471_ (.A(_0096_),
    .X(_0323_));
 sky130_fd_sc_hd__inv_2 _0472_ (.A(\mem_right_track_28.DFFR_1_.Q ),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _0473_ (.A(\mem_right_track_28.DFFR_0_.Q ),
    .Y(_0322_));
 sky130_fd_sc_hd__clkbuf_1 _0474_ (.A(\mem_right_track_28.DFFR_0_.Q ),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_1 _0475_ (.A(_0097_),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _0476_ (.A(\mem_right_track_28.DFFR_1_.Q ),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0477_ (.A(_0098_),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(\mem_right_track_26.DFFR_1_.Q ),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\mem_right_track_26.DFFR_0_.Q ),
    .Y(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _0480_ (.A(\mem_right_track_26.DFFR_0_.Q ),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_1 _0481_ (.A(_0099_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _0482_ (.A(\mem_right_track_26.DFFR_1_.Q ),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0483_ (.A(_0100_),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _0484_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .Y(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _0486_ (.A(\mem_right_track_24.DFFR_0_.Q ),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_1 _0487_ (.A(_0101_),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _0488_ (.A(\mem_right_track_24.DFFR_1_.Q ),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _0489_ (.A(_0102_),
    .X(_0311_));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(\mem_right_track_22.DFFR_1_.Q ),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_2 _0491_ (.A(\mem_right_track_22.DFFR_0_.Q ),
    .Y(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _0492_ (.A(\mem_right_track_22.DFFR_0_.Q ),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_1 _0493_ (.A(_0103_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _0494_ (.A(\mem_right_track_22.DFFR_1_.Q ),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0495_ (.A(_0104_),
    .X(_0307_));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\mem_right_track_20.DFFR_1_.Q ),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_2 _0497_ (.A(\mem_right_track_20.DFFR_0_.Q ),
    .Y(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _0498_ (.A(\mem_right_track_20.DFFR_0_.Q ),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_1 _0499_ (.A(_0105_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0500_ (.A(\mem_right_track_20.DFFR_1_.Q ),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0501_ (.A(_0106_),
    .X(_0303_));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(net61),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\mem_bottom_track_37.DFFR_0_.Q ),
    .Y(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _0504_ (.A(\mem_bottom_track_37.DFFR_0_.Q ),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0505_ (.A(_0107_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0506_ (.A(net61),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0507_ (.A(_0108_),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(\mem_bottom_track_37.DFFR_0_.Q ),
    .Y(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0509_ (.A(\mem_bottom_track_37.DFFR_0_.Q ),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0510_ (.A(_0109_),
    .X(_0298_));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(\mem_bottom_track_19.DFFR_1_.Q ),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(\mem_bottom_track_19.DFFR_0_.Q ),
    .Y(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _0513_ (.A(\mem_bottom_track_19.DFFR_0_.Q ),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0514_ (.A(_0110_),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _0515_ (.A(\mem_bottom_track_19.DFFR_1_.Q ),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _0516_ (.A(_0111_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(\mem_bottom_track_19.DFFR_0_.Q ),
    .Y(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _0518_ (.A(\mem_bottom_track_19.DFFR_0_.Q ),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0519_ (.A(_0112_),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _0522_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _0523_ (.A(_0113_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _0524_ (.A(\mem_bottom_track_17.DFFR_1_.Q ),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _0525_ (.A(_0114_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .Y(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _0527_ (.A(\mem_bottom_track_17.DFFR_0_.Q ),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_1 _0528_ (.A(_0115_),
    .X(_0286_));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(\mem_bottom_track_15.DFFR_1_.Q ),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(\mem_bottom_track_15.DFFR_0_.Q ),
    .Y(_0284_));
 sky130_fd_sc_hd__clkbuf_1 _0531_ (.A(\mem_bottom_track_15.DFFR_0_.Q ),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0532_ (.A(_0116_),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_1 _0533_ (.A(\mem_bottom_track_15.DFFR_1_.Q ),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _0534_ (.A(_0117_),
    .X(_0279_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(\mem_bottom_track_15.DFFR_0_.Q ),
    .Y(_0283_));
 sky130_fd_sc_hd__clkbuf_1 _0536_ (.A(\mem_bottom_track_15.DFFR_0_.Q ),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _0537_ (.A(_0118_),
    .X(_0280_));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(\mem_bottom_track_13.DFFR_1_.Q ),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(\mem_bottom_track_13.DFFR_0_.Q ),
    .Y(_0278_));
 sky130_fd_sc_hd__clkbuf_1 _0540_ (.A(\mem_bottom_track_13.DFFR_0_.Q ),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _0541_ (.A(_0119_),
    .X(_0275_));
 sky130_fd_sc_hd__clkbuf_1 _0542_ (.A(\mem_bottom_track_13.DFFR_1_.Q ),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0543_ (.A(_0120_),
    .X(_0273_));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(\mem_bottom_track_13.DFFR_0_.Q ),
    .Y(_0277_));
 sky130_fd_sc_hd__clkbuf_1 _0545_ (.A(\mem_bottom_track_13.DFFR_0_.Q ),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_1 _0546_ (.A(_0121_),
    .X(_0274_));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(\mem_bottom_track_11.DFFR_1_.Q ),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(\mem_bottom_track_11.DFFR_0_.Q ),
    .Y(_0272_));
 sky130_fd_sc_hd__clkbuf_1 _0549_ (.A(\mem_bottom_track_11.DFFR_0_.Q ),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _0550_ (.A(_0122_),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_1 _0551_ (.A(\mem_bottom_track_11.DFFR_1_.Q ),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_1 _0552_ (.A(_0123_),
    .X(_0267_));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(\mem_bottom_track_11.DFFR_0_.Q ),
    .Y(_0271_));
 sky130_fd_sc_hd__clkbuf_1 _0554_ (.A(\mem_bottom_track_11.DFFR_0_.Q ),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0555_ (.A(_0124_),
    .X(_0268_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(\mem_bottom_track_11.DFFR_0_.D ),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0266_));
 sky130_fd_sc_hd__clkbuf_1 _0558_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_1 _0559_ (.A(_0125_),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_1 _0560_ (.A(\mem_bottom_track_11.DFFR_0_.D ),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(_0126_),
    .X(_0261_));
 sky130_fd_sc_hd__inv_2 _0562_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .Y(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _0563_ (.A(\mem_bottom_track_9.DFFR_0_.Q ),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _0564_ (.A(_0127_),
    .X(_0262_));
 sky130_fd_sc_hd__inv_2 _0565_ (.A(\mem_bottom_track_7.DFFR_1_.Q ),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(\mem_bottom_track_7.DFFR_0_.Q ),
    .Y(_0260_));
 sky130_fd_sc_hd__clkbuf_1 _0567_ (.A(\mem_bottom_track_7.DFFR_0_.Q ),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _0568_ (.A(_0128_),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_1 _0569_ (.A(\mem_bottom_track_7.DFFR_1_.Q ),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _0570_ (.A(_0129_),
    .X(_0255_));
 sky130_fd_sc_hd__inv_2 _0571_ (.A(\mem_bottom_track_7.DFFR_0_.Q ),
    .Y(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _0572_ (.A(\mem_bottom_track_7.DFFR_0_.Q ),
    .X(_0130_));
 sky130_fd_sc_hd__clkbuf_1 _0573_ (.A(_0130_),
    .X(_0256_));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(\mem_bottom_track_5.DFFR_1_.Q ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(\mem_bottom_track_5.DFFR_0_.Q ),
    .Y(_0254_));
 sky130_fd_sc_hd__clkbuf_1 _0576_ (.A(\mem_bottom_track_5.DFFR_0_.Q ),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _0577_ (.A(_0131_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_1 _0578_ (.A(\mem_bottom_track_5.DFFR_1_.Q ),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(_0132_),
    .X(_0249_));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(\mem_bottom_track_5.DFFR_0_.Q ),
    .Y(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _0581_ (.A(\mem_bottom_track_5.DFFR_0_.Q ),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _0582_ (.A(_0133_),
    .X(_0250_));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(\mem_bottom_track_3.DFFR_1_.Q ),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _0584_ (.A(\mem_bottom_track_3.DFFR_0_.Q ),
    .Y(_0248_));
 sky130_fd_sc_hd__clkbuf_1 _0585_ (.A(\mem_bottom_track_3.DFFR_0_.Q ),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _0586_ (.A(_0134_),
    .X(_0245_));
 sky130_fd_sc_hd__clkbuf_1 _0587_ (.A(\mem_bottom_track_3.DFFR_1_.Q ),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _0588_ (.A(_0135_),
    .X(_0243_));
 sky130_fd_sc_hd__inv_2 _0589_ (.A(\mem_bottom_track_3.DFFR_0_.Q ),
    .Y(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _0590_ (.A(\mem_bottom_track_3.DFFR_0_.Q ),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _0591_ (.A(_0136_),
    .X(_0244_));
 sky130_fd_sc_hd__inv_2 _0592_ (.A(\mem_bottom_track_1.DFFR_0_.D ),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _0593_ (.A(\mem_right_track_36.DFFR_0_.Q ),
    .Y(_0242_));
 sky130_fd_sc_hd__clkbuf_1 _0594_ (.A(\mem_right_track_36.DFFR_0_.Q ),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0595_ (.A(_0137_),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_1 _0596_ (.A(\mem_bottom_track_1.DFFR_0_.D ),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0138_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(\mem_right_track_36.DFFR_0_.Q ),
    .Y(_0241_));
 sky130_fd_sc_hd__clkbuf_1 _0599_ (.A(\mem_right_track_36.DFFR_0_.Q ),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _0600_ (.A(_0139_),
    .X(_0238_));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\mem_right_track_18.DFFR_1_.Q ),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .Y(_0236_));
 sky130_fd_sc_hd__clkbuf_1 _0603_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .X(_0140_));
 sky130_fd_sc_hd__clkbuf_1 _0604_ (.A(_0140_),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_1 _0605_ (.A(\mem_right_track_18.DFFR_1_.Q ),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _0606_ (.A(_0141_),
    .X(_0231_));
 sky130_fd_sc_hd__inv_2 _0607_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .Y(_0235_));
 sky130_fd_sc_hd__clkbuf_1 _0608_ (.A(\mem_right_track_18.DFFR_0_.Q ),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_1 _0609_ (.A(_0142_),
    .X(_0232_));
 sky130_fd_sc_hd__inv_2 _0610_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _0611_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .Y(_0230_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_1 _0613_ (.A(_0143_),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_1 _0614_ (.A(\mem_right_track_16.DFFR_1_.Q ),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_1 _0615_ (.A(_0144_),
    .X(_0225_));
 sky130_fd_sc_hd__inv_2 _0616_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .Y(_0229_));
 sky130_fd_sc_hd__clkbuf_1 _0617_ (.A(\mem_right_track_16.DFFR_0_.Q ),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _0618_ (.A(_0145_),
    .X(_0226_));
 sky130_fd_sc_hd__inv_2 _0619_ (.A(\mem_right_track_14.DFFR_1_.Q ),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _0620_ (.A(\mem_right_track_14.DFFR_0_.Q ),
    .Y(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _0621_ (.A(\mem_right_track_14.DFFR_0_.Q ),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0622_ (.A(_0146_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _0623_ (.A(\mem_right_track_14.DFFR_1_.Q ),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(_0147_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _0625_ (.A(\mem_right_track_14.DFFR_0_.Q ),
    .Y(_0223_));
 sky130_fd_sc_hd__clkbuf_1 _0626_ (.A(\mem_right_track_14.DFFR_0_.Q ),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0627_ (.A(_0148_),
    .X(_0220_));
 sky130_fd_sc_hd__inv_2 _0628_ (.A(\mem_right_track_12.DFFR_1_.Q ),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _0629_ (.A(\mem_right_track_12.DFFR_0_.Q ),
    .Y(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _0630_ (.A(\mem_right_track_12.DFFR_0_.Q ),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _0631_ (.A(_0149_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(\mem_right_track_12.DFFR_1_.Q ),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_1 _0633_ (.A(_0150_),
    .X(_0213_));
 sky130_fd_sc_hd__inv_2 _0634_ (.A(\mem_right_track_12.DFFR_0_.Q ),
    .Y(_0217_));
 sky130_fd_sc_hd__clkbuf_1 _0635_ (.A(\mem_right_track_12.DFFR_0_.Q ),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _0636_ (.A(_0151_),
    .X(_0214_));
 sky130_fd_sc_hd__inv_2 _0637_ (.A(\mem_right_track_10.DFFR_1_.Q ),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .Y(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _0639_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_1 _0640_ (.A(_0152_),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_1 _0641_ (.A(\mem_right_track_10.DFFR_1_.Q ),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_1 _0642_ (.A(_0153_),
    .X(_0207_));
 sky130_fd_sc_hd__inv_2 _0643_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .Y(_0211_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(\mem_right_track_10.DFFR_0_.Q ),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_1 _0645_ (.A(_0154_),
    .X(_0208_));
 sky130_fd_sc_hd__inv_2 _0646_ (.A(\mem_right_track_10.DFFR_0_.D ),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _0647_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0649_ (.A(_0155_),
    .X(_0203_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(\mem_right_track_10.DFFR_0_.D ),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _0651_ (.A(_0156_),
    .X(_0201_));
 sky130_fd_sc_hd__inv_2 _0652_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .Y(_0205_));
 sky130_fd_sc_hd__clkbuf_1 _0653_ (.A(\mem_right_track_8.DFFR_0_.Q ),
    .X(_0157_));
 sky130_fd_sc_hd__clkbuf_1 _0654_ (.A(_0157_),
    .X(_0202_));
 sky130_fd_sc_hd__inv_2 _0655_ (.A(\mem_right_track_6.DFFR_1_.Q ),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _0656_ (.A(\mem_right_track_6.DFFR_0_.Q ),
    .Y(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _0657_ (.A(\mem_right_track_6.DFFR_0_.Q ),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0658_ (.A(_0158_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _0659_ (.A(\mem_right_track_6.DFFR_1_.Q ),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0159_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _0661_ (.A(\mem_right_track_6.DFFR_0_.Q ),
    .Y(_0199_));
 sky130_fd_sc_hd__clkbuf_1 _0662_ (.A(\mem_right_track_6.DFFR_0_.Q ),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_1 _0663_ (.A(_0160_),
    .X(_0196_));
 sky130_fd_sc_hd__inv_2 _0664_ (.A(\mem_right_track_4.DFFR_1_.Q ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _0665_ (.A(\mem_right_track_4.DFFR_0_.Q ),
    .Y(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(\mem_right_track_4.DFFR_0_.Q ),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_1 _0667_ (.A(_0161_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _0668_ (.A(\mem_right_track_4.DFFR_1_.Q ),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_1 _0669_ (.A(_0162_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _0670_ (.A(\mem_right_track_4.DFFR_0_.Q ),
    .Y(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _0671_ (.A(\mem_right_track_4.DFFR_0_.Q ),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(_0163_),
    .X(_0190_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(\mem_right_track_2.DFFR_1_.Q ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(\mem_right_track_2.DFFR_0_.Q ),
    .Y(_0188_));
 sky130_fd_sc_hd__clkbuf_1 _0675_ (.A(\mem_right_track_2.DFFR_1_.Q ),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0676_ (.A(_0164_),
    .X(_0185_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(\mem_right_track_2.DFFR_0_.Q ),
    .Y(_0187_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(\mem_right_track_2.DFFR_0_.Q ),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_1 _0679_ (.A(_0165_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(\mem_right_track_2.DFFR_0_.Q ),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_1 _0681_ (.A(_0166_),
    .X(_0183_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(\mem_right_track_0.DFFR_1_.Q ),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .Y(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0685_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _0686_ (.A(_0167_),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0687_ (.A(\mem_right_track_0.DFFR_0_.Q ),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0168_),
    .X(_0178_));
 sky130_fd_sc_hd__inv_2 _0689_ (.A(net53),
    .Y(\mux_right_track_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(net54),
    .Y(\mux_right_track_0.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_0.out ));
 sky130_fd_sc_hd__inv_2 _0692_ (.A(net39),
    .Y(\mux_right_track_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0693_ (.A(net55),
    .Y(\mux_right_track_2.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_2.out ));
 sky130_fd_sc_hd__inv_2 _0695_ (.A(net38),
    .Y(\mux_right_track_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0696_ (.A(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_4.out ));
 sky130_fd_sc_hd__inv_2 _0697_ (.A(net37),
    .Y(\mux_right_track_4.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0698_ (.A(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_6.out ));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(net36),
    .Y(\mux_right_track_6.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_8.out ));
 sky130_fd_sc_hd__inv_2 _0701_ (.A(net35),
    .Y(\mux_right_track_8.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_10.out ));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(net59),
    .Y(\mux_right_track_10.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0704_ (.A(net58),
    .Y(\mux_right_track_10.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0705_ (.A(net34),
    .Y(\mux_right_track_10.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_12.out ));
 sky130_fd_sc_hd__clkinv_2 _0707_ (.A(net60),
    .Y(\mux_right_track_12.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0708_ (.A(net33),
    .Y(\mux_right_track_12.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0709_ (.A(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_14.out ));
 sky130_fd_sc_hd__inv_2 _0710_ (.A(net51),
    .Y(\mux_right_track_14.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0711_ (.A(net32),
    .Y(\mux_right_track_14.INVTX1_2_.out ));
 sky130_fd_sc_hd__clkinv_2 _0712_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_16.out ));
 sky130_fd_sc_hd__inv_2 _0713_ (.A(net52),
    .Y(\mux_right_track_16.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkinv_2 _0714_ (.A(net49),
    .Y(\mux_right_track_16.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0715_ (.A(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_18.out ));
 sky130_fd_sc_hd__inv_2 _0716_ (.A(net48),
    .Y(\mux_right_track_18.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0717_ (.A(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_right_track_36.out ));
 sky130_fd_sc_hd__inv_2 _0718_ (.A(net40),
    .Y(\mux_right_track_36.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0719_ (.A(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_3.out ));
 sky130_fd_sc_hd__inv_2 _0720_ (.A(net10),
    .Y(\mux_bottom_track_3.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0721_ (.A(net19),
    .Y(\mux_bottom_track_3.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0722_ (.A(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_5.out ));
 sky130_fd_sc_hd__inv_2 _0723_ (.A(net18),
    .Y(\mux_bottom_track_5.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 _0724_ (.A(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_7.out ));
 sky130_fd_sc_hd__clkinv_2 _0725_ (.A(net17),
    .Y(\mux_bottom_track_7.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0726_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_9.out ));
 sky130_fd_sc_hd__inv_2 _0727_ (.A(net16),
    .Y(\mux_bottom_track_9.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_11.out ));
 sky130_fd_sc_hd__inv_2 _0729_ (.A(net4),
    .Y(\mux_bottom_track_11.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0730_ (.A(net15),
    .Y(\mux_bottom_track_11.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0731_ (.A(net5),
    .Y(\mux_bottom_track_11.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0732_ (.A(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_13.out ));
 sky130_fd_sc_hd__clkinv_2 _0733_ (.A(net14),
    .Y(\mux_bottom_track_13.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0734_ (.A(net6),
    .Y(\mux_bottom_track_13.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0735_ (.A(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_15.out ));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(net13),
    .Y(\mux_bottom_track_15.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(net7),
    .Y(\mux_bottom_track_15.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0738_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_17.out ));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(net30),
    .Y(\mux_bottom_track_17.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkinv_2 _0740_ (.A(net8),
    .Y(\mux_bottom_track_17.INVTX1_2_.out ));
 sky130_fd_sc_hd__inv_2 _0741_ (.A(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_19.out ));
 sky130_fd_sc_hd__inv_2 _0742_ (.A(net29),
    .Y(\mux_bottom_track_19.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ),
    .Y(\mux_bottom_track_37.out ));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(net21),
    .Y(\mux_bottom_track_37.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0745_ (.A(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_20.out ));
 sky130_fd_sc_hd__inv_2 _0746_ (.A(net47),
    .Y(\mux_right_track_20.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_22.out ));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(net46),
    .Y(\mux_right_track_22.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_24.out ));
 sky130_fd_sc_hd__inv_2 _0750_ (.A(net56),
    .Y(\mux_right_track_24.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0751_ (.A(net45),
    .Y(\mux_right_track_24.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0752_ (.A(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_26.out ));
 sky130_fd_sc_hd__inv_2 _0753_ (.A(net57),
    .Y(\mux_right_track_26.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0754_ (.A(net44),
    .Y(\mux_right_track_26.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0755_ (.A(\mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_28.out ));
 sky130_fd_sc_hd__inv_2 _0756_ (.A(net43),
    .Y(\mux_right_track_28.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0757_ (.A(\mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_30.out ));
 sky130_fd_sc_hd__inv_2 _0758_ (.A(net42),
    .Y(\mux_right_track_30.INVTX1_1_.out ));
 sky130_fd_sc_hd__clkinv_2 _0759_ (.A(\mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_32.out ));
 sky130_fd_sc_hd__clkinv_2 _0760_ (.A(net41),
    .Y(\mux_right_track_32.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0761_ (.A(\mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_right_track_34.out ));
 sky130_fd_sc_hd__clkinv_2 _0762_ (.A(net31),
    .Y(\mux_right_track_34.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0763_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_1.out ));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(net20),
    .Y(\mux_bottom_track_1.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(net9),
    .Y(\mux_bottom_track_1.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0766_ (.A(\mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_23.out ));
 sky130_fd_sc_hd__inv_2 _0767_ (.A(net27),
    .Y(\mux_bottom_track_23.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(net1),
    .Y(\mux_bottom_track_23.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0769_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_25.out ));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(net26),
    .Y(\mux_bottom_track_25.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(net2),
    .Y(\mux_bottom_track_25.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0772_ (.A(\mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_27.out ));
 sky130_fd_sc_hd__inv_2 _0773_ (.A(net25),
    .Y(\mux_bottom_track_27.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0774_ (.A(net3),
    .Y(\mux_bottom_track_27.INVTX1_1_.out ));
 sky130_fd_sc_hd__inv_2 _0775_ (.A(\mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_29.out ));
 sky130_fd_sc_hd__inv_2 _0776_ (.A(net24),
    .Y(\mux_bottom_track_29.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0777_ (.A(\mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_31.out ));
 sky130_fd_sc_hd__inv_2 _0778_ (.A(net23),
    .Y(\mux_bottom_track_31.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0779_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_33.out ));
 sky130_fd_sc_hd__clkinv_2 _0780_ (.A(net22),
    .Y(\mux_bottom_track_33.INVTX1_0_.out ));
 sky130_fd_sc_hd__inv_2 _0781_ (.A(\mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .Y(\mux_bottom_track_35.out ));
 sky130_fd_sc_hd__inv_2 _0782_ (.A(net12),
    .Y(\mux_bottom_track_35.INVTX1_0_.out ));
 sky130_fd_sc_hd__clkbuf_4 _0783_ (.A(net50),
    .X(_0169_));
 sky130_fd_sc_hd__buf_4 _0784_ (.A(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__inv_2 _0785_ (.A(_0170_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _0786_ (.A(_0170_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _0787_ (.A(_0170_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _0788_ (.A(_0170_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _0789_ (.A(_0170_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _0790_ (.A(_0170_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _0791_ (.A(_0170_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _0792_ (.A(_0170_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _0793_ (.A(_0170_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _0794_ (.A(_0170_),
    .Y(_0051_));
 sky130_fd_sc_hd__buf_4 _0795_ (.A(_0169_),
    .X(_0171_));
 sky130_fd_sc_hd__inv_2 _0796_ (.A(_0171_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _0797_ (.A(_0171_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(_0171_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(_0171_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(_0171_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _0801_ (.A(_0171_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _0802_ (.A(_0171_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _0803_ (.A(_0171_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(_0171_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(_0171_),
    .Y(_0061_));
 sky130_fd_sc_hd__buf_4 _0806_ (.A(_0169_),
    .X(_0172_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(_0172_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _0808_ (.A(_0172_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _0809_ (.A(_0172_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _0810_ (.A(_0172_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _0811_ (.A(_0172_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _0812_ (.A(_0172_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _0813_ (.A(_0172_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(_0172_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _0815_ (.A(_0172_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _0816_ (.A(_0172_),
    .Y(_0071_));
 sky130_fd_sc_hd__buf_4 _0817_ (.A(_0169_),
    .X(_0173_));
 sky130_fd_sc_hd__inv_2 _0818_ (.A(_0173_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _0819_ (.A(_0173_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _0820_ (.A(_0173_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(_0173_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0822_ (.A(_0173_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(_0173_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0824_ (.A(_0173_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0825_ (.A(_0173_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0826_ (.A(_0173_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(_0173_),
    .Y(_0007_));
 sky130_fd_sc_hd__buf_4 _0828_ (.A(_0169_),
    .X(_0174_));
 sky130_fd_sc_hd__inv_2 _0829_ (.A(_0174_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0830_ (.A(_0174_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0831_ (.A(_0174_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0832_ (.A(_0174_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0833_ (.A(_0174_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0834_ (.A(_0174_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _0835_ (.A(_0174_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(_0174_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _0837_ (.A(_0174_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _0838_ (.A(_0174_),
    .Y(_0017_));
 sky130_fd_sc_hd__buf_4 _0839_ (.A(_0169_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _0840_ (.A(_0175_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0175_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _0842_ (.A(_0175_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(_0175_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(_0175_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _0845_ (.A(_0175_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _0846_ (.A(_0175_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _0847_ (.A(_0175_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _0848_ (.A(_0175_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _0849_ (.A(_0175_),
    .Y(_0027_));
 sky130_fd_sc_hd__buf_4 _0850_ (.A(net50),
    .X(_0176_));
 sky130_fd_sc_hd__inv_2 _0851_ (.A(_0176_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _0852_ (.A(_0176_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _0853_ (.A(_0176_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _0854_ (.A(_0176_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _0855_ (.A(_0176_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _0856_ (.A(_0176_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _0857_ (.A(_0176_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _0858_ (.A(_0176_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _0859_ (.A(_0176_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _0860_ (.A(_0176_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _0861_ (.A(_0169_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0862_ (.A(_0169_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _0863_ (.A(_0169_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _0864_ (.A(_0169_),
    .Y(_0041_));
 sky130_fd_sc_hd__dfrtp_2 _0865_ (.CLK(prog_clk),
    .D(\mem_right_track_0.DFFR_0_.Q ),
    .RESET_B(_0042_),
    .Q(\mem_right_track_0.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0866_ (.CLK(prog_clk),
    .D(net11),
    .RESET_B(_0043_),
    .Q(\mem_right_track_0.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0867_ (.CLK(prog_clk),
    .D(\mem_right_track_2.DFFR_0_.Q ),
    .RESET_B(_0044_),
    .Q(\mem_right_track_2.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0868_ (.CLK(prog_clk),
    .D(\mem_right_track_0.DFFR_1_.Q ),
    .RESET_B(_0045_),
    .Q(\mem_right_track_2.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0869_ (.CLK(prog_clk),
    .D(\mem_right_track_4.DFFR_0_.Q ),
    .RESET_B(_0046_),
    .Q(\mem_right_track_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0870_ (.CLK(prog_clk),
    .D(\mem_right_track_2.DFFR_1_.Q ),
    .RESET_B(_0047_),
    .Q(\mem_right_track_4.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0871_ (.CLK(prog_clk),
    .D(\mem_right_track_6.DFFR_0_.Q ),
    .RESET_B(_0048_),
    .Q(\mem_right_track_6.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0872_ (.CLK(prog_clk),
    .D(\mem_right_track_4.DFFR_1_.Q ),
    .RESET_B(_0049_),
    .Q(\mem_right_track_6.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0873_ (.CLK(prog_clk),
    .D(\mem_right_track_8.DFFR_0_.Q ),
    .RESET_B(_0050_),
    .Q(\mem_right_track_10.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0874_ (.CLK(prog_clk),
    .D(\mem_right_track_6.DFFR_1_.Q ),
    .RESET_B(_0051_),
    .Q(\mem_right_track_8.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0875_ (.CLK(prog_clk),
    .D(\mem_right_track_10.DFFR_0_.Q ),
    .RESET_B(_0052_),
    .Q(\mem_right_track_10.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0876_ (.CLK(prog_clk),
    .D(\mem_right_track_10.DFFR_0_.D ),
    .RESET_B(_0053_),
    .Q(\mem_right_track_10.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0877_ (.CLK(prog_clk),
    .D(\mem_right_track_12.DFFR_0_.Q ),
    .RESET_B(_0054_),
    .Q(\mem_right_track_12.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0878_ (.CLK(prog_clk),
    .D(\mem_right_track_10.DFFR_1_.Q ),
    .RESET_B(_0055_),
    .Q(\mem_right_track_12.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0879_ (.CLK(prog_clk),
    .D(\mem_right_track_14.DFFR_0_.Q ),
    .RESET_B(_0056_),
    .Q(\mem_right_track_14.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0880_ (.CLK(prog_clk),
    .D(\mem_right_track_12.DFFR_1_.Q ),
    .RESET_B(_0057_),
    .Q(\mem_right_track_14.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0881_ (.CLK(prog_clk),
    .D(\mem_right_track_16.DFFR_0_.Q ),
    .RESET_B(_0058_),
    .Q(\mem_right_track_16.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0882_ (.CLK(prog_clk),
    .D(\mem_right_track_14.DFFR_1_.Q ),
    .RESET_B(_0059_),
    .Q(\mem_right_track_16.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0883_ (.CLK(prog_clk),
    .D(\mem_right_track_18.DFFR_0_.Q ),
    .RESET_B(_0060_),
    .Q(\mem_right_track_18.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0884_ (.CLK(prog_clk),
    .D(\mem_right_track_16.DFFR_1_.Q ),
    .RESET_B(_0061_),
    .Q(\mem_right_track_18.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0885_ (.CLK(prog_clk),
    .D(\mem_right_track_36.DFFR_0_.Q ),
    .RESET_B(_0062_),
    .Q(\mem_bottom_track_1.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0886_ (.CLK(prog_clk),
    .D(\mem_right_track_34.DFFR_1_.Q ),
    .RESET_B(_0063_),
    .Q(\mem_right_track_36.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0887_ (.CLK(prog_clk),
    .D(\mem_bottom_track_3.DFFR_0_.Q ),
    .RESET_B(_0064_),
    .Q(\mem_bottom_track_3.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0888_ (.CLK(prog_clk),
    .D(\mem_bottom_track_1.DFFR_1_.Q ),
    .RESET_B(_0065_),
    .Q(\mem_bottom_track_3.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0889_ (.CLK(prog_clk),
    .D(\mem_bottom_track_5.DFFR_0_.Q ),
    .RESET_B(_0066_),
    .Q(\mem_bottom_track_5.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0890_ (.CLK(prog_clk),
    .D(\mem_bottom_track_3.DFFR_1_.Q ),
    .RESET_B(_0067_),
    .Q(\mem_bottom_track_5.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0891_ (.CLK(prog_clk),
    .D(\mem_bottom_track_7.DFFR_0_.Q ),
    .RESET_B(_0068_),
    .Q(\mem_bottom_track_7.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0892_ (.CLK(prog_clk),
    .D(\mem_bottom_track_5.DFFR_1_.Q ),
    .RESET_B(_0069_),
    .Q(\mem_bottom_track_7.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0893_ (.CLK(prog_clk),
    .D(\mem_bottom_track_9.DFFR_0_.Q ),
    .RESET_B(_0070_),
    .Q(\mem_bottom_track_11.DFFR_0_.D ));
 sky130_fd_sc_hd__dfrtp_4 _0894_ (.CLK(prog_clk),
    .D(\mem_bottom_track_7.DFFR_1_.Q ),
    .RESET_B(_0071_),
    .Q(\mem_bottom_track_9.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0895_ (.CLK(prog_clk),
    .D(\mem_bottom_track_11.DFFR_0_.Q ),
    .RESET_B(_0072_),
    .Q(\mem_bottom_track_11.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0896_ (.CLK(prog_clk),
    .D(\mem_bottom_track_11.DFFR_0_.D ),
    .RESET_B(_0073_),
    .Q(\mem_bottom_track_11.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0897_ (.CLK(prog_clk),
    .D(\mem_bottom_track_13.DFFR_0_.Q ),
    .RESET_B(_0000_),
    .Q(\mem_bottom_track_13.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0898_ (.CLK(prog_clk),
    .D(\mem_bottom_track_11.DFFR_1_.Q ),
    .RESET_B(_0001_),
    .Q(\mem_bottom_track_13.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0899_ (.CLK(prog_clk),
    .D(\mem_bottom_track_15.DFFR_0_.Q ),
    .RESET_B(_0002_),
    .Q(\mem_bottom_track_15.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0900_ (.CLK(prog_clk),
    .D(\mem_bottom_track_13.DFFR_1_.Q ),
    .RESET_B(_0003_),
    .Q(\mem_bottom_track_15.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0901_ (.CLK(prog_clk),
    .D(\mem_bottom_track_17.DFFR_0_.Q ),
    .RESET_B(_0004_),
    .Q(\mem_bottom_track_17.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0902_ (.CLK(prog_clk),
    .D(\mem_bottom_track_15.DFFR_1_.Q ),
    .RESET_B(_0005_),
    .Q(\mem_bottom_track_17.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0903_ (.CLK(prog_clk),
    .D(\mem_bottom_track_19.DFFR_0_.Q ),
    .RESET_B(_0006_),
    .Q(\mem_bottom_track_19.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0904_ (.CLK(prog_clk),
    .D(\mem_bottom_track_17.DFFR_1_.Q ),
    .RESET_B(_0007_),
    .Q(\mem_bottom_track_19.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0905_ (.CLK(prog_clk),
    .D(\mem_bottom_track_37.DFFR_0_.Q ),
    .RESET_B(_0008_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_4 _0906_ (.CLK(prog_clk),
    .D(\mem_bottom_track_35.DFFR_1_.Q ),
    .RESET_B(_0009_),
    .Q(\mem_bottom_track_37.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0907_ (.CLK(prog_clk),
    .D(\mem_right_track_20.DFFR_0_.Q ),
    .RESET_B(_0010_),
    .Q(\mem_right_track_20.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0908_ (.CLK(prog_clk),
    .D(\mem_right_track_18.DFFR_1_.Q ),
    .RESET_B(_0011_),
    .Q(\mem_right_track_20.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0909_ (.CLK(prog_clk),
    .D(\mem_right_track_22.DFFR_0_.Q ),
    .RESET_B(_0012_),
    .Q(\mem_right_track_22.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0910_ (.CLK(prog_clk),
    .D(\mem_right_track_20.DFFR_1_.Q ),
    .RESET_B(_0013_),
    .Q(\mem_right_track_22.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0911_ (.CLK(prog_clk),
    .D(\mem_right_track_24.DFFR_0_.Q ),
    .RESET_B(_0014_),
    .Q(\mem_right_track_24.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0912_ (.CLK(prog_clk),
    .D(\mem_right_track_22.DFFR_1_.Q ),
    .RESET_B(_0015_),
    .Q(\mem_right_track_24.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_4 _0913_ (.CLK(prog_clk),
    .D(\mem_right_track_26.DFFR_0_.Q ),
    .RESET_B(_0016_),
    .Q(\mem_right_track_26.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0914_ (.CLK(prog_clk),
    .D(\mem_right_track_24.DFFR_1_.Q ),
    .RESET_B(_0017_),
    .Q(\mem_right_track_26.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0915_ (.CLK(prog_clk),
    .D(\mem_right_track_28.DFFR_0_.Q ),
    .RESET_B(_0018_),
    .Q(\mem_right_track_28.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0916_ (.CLK(prog_clk),
    .D(\mem_right_track_26.DFFR_1_.Q ),
    .RESET_B(_0019_),
    .Q(\mem_right_track_28.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0917_ (.CLK(prog_clk),
    .D(\mem_right_track_30.DFFR_0_.Q ),
    .RESET_B(_0020_),
    .Q(\mem_right_track_30.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0918_ (.CLK(prog_clk),
    .D(\mem_right_track_28.DFFR_1_.Q ),
    .RESET_B(_0021_),
    .Q(\mem_right_track_30.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0919_ (.CLK(prog_clk),
    .D(\mem_right_track_32.DFFR_0_.Q ),
    .RESET_B(_0022_),
    .Q(\mem_right_track_32.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0920_ (.CLK(prog_clk),
    .D(\mem_right_track_30.DFFR_1_.Q ),
    .RESET_B(_0023_),
    .Q(\mem_right_track_32.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0921_ (.CLK(prog_clk),
    .D(\mem_right_track_34.DFFR_0_.Q ),
    .RESET_B(_0024_),
    .Q(\mem_right_track_34.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0922_ (.CLK(prog_clk),
    .D(\mem_right_track_32.DFFR_1_.Q ),
    .RESET_B(_0025_),
    .Q(\mem_right_track_34.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0923_ (.CLK(prog_clk),
    .D(\mem_bottom_track_1.DFFR_0_.Q ),
    .RESET_B(_0026_),
    .Q(\mem_bottom_track_1.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0924_ (.CLK(prog_clk),
    .D(\mem_bottom_track_1.DFFR_0_.D ),
    .RESET_B(_0027_),
    .Q(\mem_bottom_track_1.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0925_ (.CLK(prog_clk),
    .D(\mem_bottom_track_23.DFFR_0_.Q ),
    .RESET_B(_0028_),
    .Q(\mem_bottom_track_23.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0926_ (.CLK(prog_clk),
    .D(\mem_bottom_track_19.DFFR_1_.Q ),
    .RESET_B(_0029_),
    .Q(\mem_bottom_track_23.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0927_ (.CLK(prog_clk),
    .D(\mem_bottom_track_25.DFFR_0_.Q ),
    .RESET_B(_0030_),
    .Q(\mem_bottom_track_25.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0928_ (.CLK(prog_clk),
    .D(\mem_bottom_track_23.DFFR_1_.Q ),
    .RESET_B(_0031_),
    .Q(\mem_bottom_track_25.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0929_ (.CLK(prog_clk),
    .D(\mem_bottom_track_27.DFFR_0_.Q ),
    .RESET_B(_0032_),
    .Q(\mem_bottom_track_27.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0930_ (.CLK(prog_clk),
    .D(\mem_bottom_track_25.DFFR_1_.Q ),
    .RESET_B(_0033_),
    .Q(\mem_bottom_track_27.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0931_ (.CLK(prog_clk),
    .D(\mem_bottom_track_29.DFFR_0_.Q ),
    .RESET_B(_0034_),
    .Q(\mem_bottom_track_29.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0932_ (.CLK(prog_clk),
    .D(\mem_bottom_track_27.DFFR_1_.Q ),
    .RESET_B(_0035_),
    .Q(\mem_bottom_track_29.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0933_ (.CLK(prog_clk),
    .D(\mem_bottom_track_31.DFFR_0_.Q ),
    .RESET_B(_0036_),
    .Q(\mem_bottom_track_31.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0934_ (.CLK(prog_clk),
    .D(\mem_bottom_track_29.DFFR_1_.Q ),
    .RESET_B(_0037_),
    .Q(\mem_bottom_track_31.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0935_ (.CLK(prog_clk),
    .D(\mem_bottom_track_33.DFFR_0_.Q ),
    .RESET_B(_0038_),
    .Q(\mem_bottom_track_33.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_1 _0936_ (.CLK(prog_clk),
    .D(\mem_bottom_track_31.DFFR_1_.Q ),
    .RESET_B(_0039_),
    .Q(\mem_bottom_track_33.DFFR_0_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0937_ (.CLK(prog_clk),
    .D(\mem_bottom_track_35.DFFR_0_.Q ),
    .RESET_B(_0040_),
    .Q(\mem_bottom_track_35.DFFR_1_.Q ));
 sky130_fd_sc_hd__dfrtp_2 _0938_ (.CLK(prog_clk),
    .D(\mem_bottom_track_33.DFFR_1_.Q ),
    .RESET_B(_0041_),
    .Q(\mem_bottom_track_35.DFFR_0_.Q ));
 sky130_fd_sc_hd__conb_1 _1021__101 (.HI(net101));
 sky130_fd_sc_hd__conb_1 _1027__102 (.HI(net102));
 sky130_fd_sc_hd__conb_1 _1033__103 (.HI(net103));
 sky130_fd_sc_hd__conb_1 _1039__104 (.HI(net104));
 sky130_fd_sc_hd__conb_1 _1045__105 (.HI(net105));
 sky130_fd_sc_hd__conb_1 _1051__106 (.HI(net106));
 sky130_fd_sc_hd__conb_1 _1057__107 (.HI(net107));
 sky130_fd_sc_hd__conb_1 _1063__108 (.HI(net108));
 sky130_fd_sc_hd__conb_1 _1069__109 (.HI(net109));
 sky130_fd_sc_hd__conb_1 _1075__110 (.HI(net110));
 sky130_fd_sc_hd__conb_1 _1081__111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 _1087__112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 _1093__113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 _1099__114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 _1105__115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 _1111__116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 _1117__117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 _1123__118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 _1129__119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 _1135__120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 _1140__121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 _1144__122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 _1148__123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 _1152__124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 _1156__125 (.HI(net125));
 sky130_fd_sc_hd__conb_1 _1160__126 (.HI(net126));
 sky130_fd_sc_hd__conb_1 _1164__127 (.HI(net127));
 sky130_fd_sc_hd__conb_1 _1168__128 (.HI(net128));
 sky130_fd_sc_hd__conb_1 _1172__129 (.HI(net129));
 sky130_fd_sc_hd__conb_1 _1176__130 (.HI(net130));
 sky130_fd_sc_hd__conb_1 _1180__131 (.HI(net131));
 sky130_fd_sc_hd__conb_1 _1184__132 (.HI(net132));
 sky130_fd_sc_hd__conb_1 _1188__133 (.HI(net133));
 sky130_fd_sc_hd__conb_1 _1192__134 (.HI(net134));
 sky130_fd_sc_hd__conb_1 _1196__135 (.HI(net135));
 sky130_fd_sc_hd__conb_1 _1200__136 (.HI(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\mem_right_track_12.DFFR_1_.Q ));
 sky130_fd_sc_hd__clkbuf_1 _0976_ (.A(\mux_right_track_36.out ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(\mux_right_track_34.out ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _0978_ (.A(\mux_right_track_32.out ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _0979_ (.A(\mux_right_track_30.out ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(\mux_right_track_28.out ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _0981_ (.A(\mux_right_track_26.out ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _0982_ (.A(\mux_right_track_24.out ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(\mux_right_track_22.out ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _0984_ (.A(\mux_right_track_20.out ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(\mux_right_track_18.out ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _0986_ (.A(\mux_right_track_16.out ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _0987_ (.A(\mux_right_track_14.out ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _0988_ (.A(\mux_right_track_12.out ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _0989_ (.A(\mux_right_track_10.out ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _0990_ (.A(\mux_right_track_8.out ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(\mux_right_track_6.out ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(\mux_right_track_4.out ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _0993_ (.A(\mux_right_track_2.out ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(\mux_right_track_0.out ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _0995_ (.A(\mux_bottom_track_37.out ),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _0996_ (.A(\mux_bottom_track_35.out ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 _0997_ (.A(\mux_bottom_track_33.out ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(\mux_bottom_track_31.out ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(\mux_bottom_track_29.out ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(\mux_bottom_track_27.out ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(\mux_bottom_track_25.out ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _1002_ (.A(\mux_bottom_track_23.out ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(net28),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _1004_ (.A(\mux_bottom_track_19.out ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _1005_ (.A(\mux_bottom_track_17.out ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(\mux_bottom_track_15.out ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(\mux_bottom_track_13.out ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _1008_ (.A(\mux_bottom_track_11.out ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _1009_ (.A(\mux_bottom_track_9.out ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _1010_ (.A(\mux_bottom_track_7.out ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 _1011_ (.A(\mux_bottom_track_5.out ),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(\mux_bottom_track_3.out ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 _1013_ (.A(\mux_bottom_track_1.out ),
    .X(net81));
 sky130_fd_sc_hd__ebufn_2 _1014_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0177_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1015_ (.A(net100),
    .TE_B(_0178_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1016_ (.A(\mux_right_track_0.INVTX1_1_.out ),
    .TE_B(_0179_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1017_ (.A(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0180_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1018_ (.A(\mux_right_track_0.INVTX1_0_.out ),
    .TE_B(_0181_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1019_ (.A(\mux_right_track_0.INVTX1_2_.out ),
    .TE_B(_0182_),
    .Z(\mux_right_track_0.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1020_ (.A(\mux_right_track_2.INVTX1_1_.out ),
    .TE_B(_0183_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1021_ (.A(net101),
    .TE_B(_0184_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1022_ (.A(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0185_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1023_ (.A(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0186_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1024_ (.A(\mux_right_track_2.INVTX1_2_.out ),
    .TE_B(_0187_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1025_ (.A(\mux_right_track_0.INVTX1_1_.out ),
    .TE_B(_0188_),
    .Z(\mux_right_track_2.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1026_ (.A(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0189_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1027_ (.A(net102),
    .TE_B(_0190_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1028_ (.A(\mux_right_track_24.INVTX1_0_.out ),
    .TE_B(_0191_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1029_ (.A(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0192_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1030_ (.A(\mux_right_track_4.INVTX1_2_.out ),
    .TE_B(_0193_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1031_ (.A(\mux_right_track_2.INVTX1_1_.out ),
    .TE_B(_0194_),
    .Z(\mux_right_track_4.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1032_ (.A(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0195_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1033_ (.A(net103),
    .TE_B(_0196_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1034_ (.A(\mux_right_track_26.INVTX1_0_.out ),
    .TE_B(_0197_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1035_ (.A(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0198_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1036_ (.A(\mux_right_track_6.INVTX1_2_.out ),
    .TE_B(_0199_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1037_ (.A(\mux_right_track_24.INVTX1_0_.out ),
    .TE_B(_0200_),
    .Z(\mux_right_track_6.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1038_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0201_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1039_ (.A(net104),
    .TE_B(_0202_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1040_ (.A(\mux_right_track_10.INVTX1_0_.out ),
    .TE_B(_0203_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1041_ (.A(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0204_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1042_ (.A(\mux_right_track_8.INVTX1_2_.out ),
    .TE_B(_0205_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1043_ (.A(\mux_right_track_26.INVTX1_0_.out ),
    .TE_B(_0206_),
    .Z(\mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1044_ (.A(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0207_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1045_ (.A(net105),
    .TE_B(_0208_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1046_ (.A(\mux_right_track_10.INVTX1_1_.out ),
    .TE_B(_0209_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1047_ (.A(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0210_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1048_ (.A(\mux_right_track_10.INVTX1_2_.out ),
    .TE_B(_0211_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1049_ (.A(\mux_right_track_10.INVTX1_0_.out ),
    .TE_B(_0212_),
    .Z(\mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1050_ (.A(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0213_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1051_ (.A(net106),
    .TE_B(_0214_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1052_ (.A(\mux_right_track_12.INVTX1_1_.out ),
    .TE_B(_0215_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1053_ (.A(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0216_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_2 _1054_ (.A(\mux_right_track_12.INVTX1_2_.out ),
    .TE_B(_0217_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1055_ (.A(\mux_right_track_10.INVTX1_1_.out ),
    .TE_B(_0218_),
    .Z(\mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1056_ (.A(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0219_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1057_ (.A(net107),
    .TE_B(_0220_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1058_ (.A(\mux_right_track_14.INVTX1_1_.out ),
    .TE_B(_0221_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1059_ (.A(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0222_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1060_ (.A(\mux_right_track_14.INVTX1_2_.out ),
    .TE_B(_0223_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1061_ (.A(\mux_right_track_12.INVTX1_1_.out ),
    .TE_B(_0224_),
    .Z(\mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1062_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0225_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1063_ (.A(net108),
    .TE_B(_0226_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1064_ (.A(\mux_right_track_16.INVTX1_1_.out ),
    .TE_B(_0227_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1065_ (.A(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0228_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1066_ (.A(\mux_right_track_16.INVTX1_2_.out ),
    .TE_B(_0229_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1067_ (.A(\mux_right_track_14.INVTX1_1_.out ),
    .TE_B(_0230_),
    .Z(\mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1068_ (.A(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0231_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1069_ (.A(net109),
    .TE_B(_0232_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1070_ (.A(\mux_right_track_16.INVTX1_1_.out ),
    .TE_B(_0233_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1071_ (.A(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0234_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1072_ (.A(\mux_right_track_18.INVTX1_2_.out ),
    .TE_B(_0235_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1073_ (.A(\mux_right_track_0.INVTX1_0_.out ),
    .TE_B(_0236_),
    .Z(\mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1074_ (.A(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0237_),
    .Z(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1075_ (.A(net110),
    .TE_B(_0238_),
    .Z(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1076_ (.A(\mux_right_track_16.INVTX1_1_.out ),
    .TE_B(_0239_),
    .Z(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1077_ (.A(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0240_),
    .Z(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1078_ (.A(\mux_right_track_36.INVTX1_2_.out ),
    .TE_B(_0241_),
    .Z(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1079_ (.A(\mux_right_track_0.INVTX1_0_.out ),
    .TE_B(_0242_),
    .Z(\mux_right_track_36.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1080_ (.A(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0243_),
    .Z(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1081_ (.A(net111),
    .TE_B(_0244_),
    .Z(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1082_ (.A(\mux_bottom_track_3.INVTX1_1_.out ),
    .TE_B(_0245_),
    .Z(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1083_ (.A(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0246_),
    .Z(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1084_ (.A(\mux_bottom_track_23.INVTX1_1_.out ),
    .TE_B(_0247_),
    .Z(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1085_ (.A(\mux_bottom_track_3.INVTX1_0_.out ),
    .TE_B(_0248_),
    .Z(\mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1086_ (.A(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0249_),
    .Z(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1087_ (.A(net112),
    .TE_B(_0250_),
    .Z(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1088_ (.A(\mux_bottom_track_23.INVTX1_1_.out ),
    .TE_B(_0251_),
    .Z(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1089_ (.A(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0252_),
    .Z(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1090_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0253_),
    .Z(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1091_ (.A(\mux_bottom_track_5.INVTX1_0_.out ),
    .TE_B(_0254_),
    .Z(\mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1092_ (.A(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0255_),
    .Z(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1093_ (.A(net113),
    .TE_B(_0256_),
    .Z(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1094_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0257_),
    .Z(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1095_ (.A(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0258_),
    .Z(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1096_ (.A(\mux_bottom_track_27.INVTX1_1_.out ),
    .TE_B(_0259_),
    .Z(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1097_ (.A(\mux_bottom_track_7.INVTX1_0_.out ),
    .TE_B(_0260_),
    .Z(\mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1098_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0261_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1099_ (.A(net114),
    .TE_B(_0262_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1100_ (.A(\mux_bottom_track_27.INVTX1_1_.out ),
    .TE_B(_0263_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1101_ (.A(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0264_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1102_ (.A(\mux_bottom_track_11.INVTX1_1_.out ),
    .TE_B(_0265_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1103_ (.A(\mux_bottom_track_9.INVTX1_0_.out ),
    .TE_B(_0266_),
    .Z(\mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1104_ (.A(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0267_),
    .Z(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1105_ (.A(net115),
    .TE_B(_0268_),
    .Z(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1106_ (.A(\mux_bottom_track_11.INVTX1_1_.out ),
    .TE_B(_0269_),
    .Z(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1107_ (.A(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0270_),
    .Z(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1108_ (.A(\mux_bottom_track_11.INVTX1_2_.out ),
    .TE_B(_0271_),
    .Z(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1109_ (.A(\mux_bottom_track_11.INVTX1_0_.out ),
    .TE_B(_0272_),
    .Z(\mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1110_ (.A(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0273_),
    .Z(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1111_ (.A(net116),
    .TE_B(_0274_),
    .Z(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1112_ (.A(\mux_bottom_track_11.INVTX1_2_.out ),
    .TE_B(_0275_),
    .Z(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1113_ (.A(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0276_),
    .Z(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1114_ (.A(\mux_bottom_track_13.INVTX1_2_.out ),
    .TE_B(_0277_),
    .Z(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1115_ (.A(\mux_bottom_track_13.INVTX1_0_.out ),
    .TE_B(_0278_),
    .Z(\mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1116_ (.A(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0279_),
    .Z(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1117_ (.A(net117),
    .TE_B(_0280_),
    .Z(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1118_ (.A(\mux_bottom_track_13.INVTX1_2_.out ),
    .TE_B(_0281_),
    .Z(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1119_ (.A(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0282_),
    .Z(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1120_ (.A(\mux_bottom_track_15.INVTX1_2_.out ),
    .TE_B(_0283_),
    .Z(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1121_ (.A(\mux_bottom_track_15.INVTX1_0_.out ),
    .TE_B(_0284_),
    .Z(\mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1122_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0285_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1123_ (.A(net118),
    .TE_B(_0286_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1124_ (.A(\mux_bottom_track_15.INVTX1_2_.out ),
    .TE_B(_0287_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1125_ (.A(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0288_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1126_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0289_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1127_ (.A(\mux_bottom_track_17.INVTX1_0_.out ),
    .TE_B(_0290_),
    .Z(\mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1128_ (.A(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0291_),
    .Z(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1129_ (.A(net119),
    .TE_B(_0292_),
    .Z(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1130_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0293_),
    .Z(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1131_ (.A(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0294_),
    .Z(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1132_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0295_),
    .Z(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1133_ (.A(\mux_bottom_track_19.INVTX1_0_.out ),
    .TE_B(_0296_),
    .Z(\mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1134_ (.A(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ),
    .TE_B(_0297_),
    .Z(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1135_ (.A(net120),
    .TE_B(_0298_),
    .Z(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1136_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0299_),
    .Z(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1137_ (.A(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0300_),
    .Z(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out ));
 sky130_fd_sc_hd__ebufn_1 _1138_ (.A(\mux_bottom_track_17.INVTX1_2_.out ),
    .TE_B(_0301_),
    .Z(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1139_ (.A(\mux_bottom_track_37.INVTX1_0_.out ),
    .TE_B(_0302_),
    .Z(\mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1140_ (.A(net121),
    .TE_B(_0303_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1141_ (.A(\mux_right_track_20.INVTX1_1_.out ),
    .TE_B(_0304_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1142_ (.A(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0305_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1143_ (.A(\mux_right_track_0.INVTX1_1_.out ),
    .TE_B(_0306_),
    .Z(\mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1144_ (.A(net122),
    .TE_B(_0307_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1145_ (.A(\mux_right_track_22.INVTX1_1_.out ),
    .TE_B(_0308_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1146_ (.A(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0309_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1147_ (.A(\mux_right_track_2.INVTX1_1_.out ),
    .TE_B(_0310_),
    .Z(\mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1148_ (.A(net123),
    .TE_B(_0311_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1149_ (.A(\mux_right_track_24.INVTX1_1_.out ),
    .TE_B(_0312_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1150_ (.A(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0313_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1151_ (.A(\mux_right_track_24.INVTX1_0_.out ),
    .TE_B(_0314_),
    .Z(\mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1152_ (.A(net124),
    .TE_B(_0315_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1153_ (.A(\mux_right_track_26.INVTX1_1_.out ),
    .TE_B(_0316_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1154_ (.A(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0317_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1155_ (.A(\mux_right_track_26.INVTX1_0_.out ),
    .TE_B(_0318_),
    .Z(\mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1156_ (.A(net125),
    .TE_B(_0319_),
    .Z(\mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1157_ (.A(\mux_right_track_28.INVTX1_1_.out ),
    .TE_B(_0320_),
    .Z(\mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1158_ (.A(\mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0321_),
    .Z(\mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1159_ (.A(\mux_right_track_10.INVTX1_0_.out ),
    .TE_B(_0322_),
    .Z(\mux_right_track_28.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1160_ (.A(net126),
    .TE_B(_0323_),
    .Z(\mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1161_ (.A(\mux_right_track_30.INVTX1_1_.out ),
    .TE_B(_0324_),
    .Z(\mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1162_ (.A(\mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0325_),
    .Z(\mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1163_ (.A(\mux_right_track_10.INVTX1_1_.out ),
    .TE_B(_0326_),
    .Z(\mux_right_track_30.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1164_ (.A(net127),
    .TE_B(_0327_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1165_ (.A(\mux_right_track_32.INVTX1_1_.out ),
    .TE_B(_0328_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1166_ (.A(\mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0329_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1167_ (.A(\mux_right_track_12.INVTX1_1_.out ),
    .TE_B(_0330_),
    .Z(\mux_right_track_32.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1168_ (.A(net128),
    .TE_B(_0331_),
    .Z(\mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1169_ (.A(\mux_right_track_34.INVTX1_1_.out ),
    .TE_B(_0332_),
    .Z(\mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1170_ (.A(\mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0333_),
    .Z(\mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1171_ (.A(\mux_right_track_14.INVTX1_1_.out ),
    .TE_B(_0334_),
    .Z(\mux_right_track_34.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1172_ (.A(net129),
    .TE_B(_0335_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1173_ (.A(\mux_bottom_track_1.INVTX1_1_.out ),
    .TE_B(_0336_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1174_ (.A(\mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0337_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1175_ (.A(\mux_bottom_track_1.INVTX1_0_.out ),
    .TE_B(_0338_),
    .Z(\mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1176_ (.A(net130),
    .TE_B(_0339_),
    .Z(\mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1177_ (.A(\mux_bottom_track_23.INVTX1_1_.out ),
    .TE_B(_0340_),
    .Z(\mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1178_ (.A(\mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0341_),
    .Z(\mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1179_ (.A(\mux_bottom_track_23.INVTX1_0_.out ),
    .TE_B(_0342_),
    .Z(\mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1180_ (.A(net131),
    .TE_B(_0343_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1181_ (.A(\mux_bottom_track_25.INVTX1_1_.out ),
    .TE_B(_0344_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1182_ (.A(\mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0345_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1183_ (.A(\mux_bottom_track_25.INVTX1_0_.out ),
    .TE_B(_0346_),
    .Z(\mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1184_ (.A(net132),
    .TE_B(_0347_),
    .Z(\mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1185_ (.A(\mux_bottom_track_27.INVTX1_1_.out ),
    .TE_B(_0348_),
    .Z(\mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1186_ (.A(\mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0349_),
    .Z(\mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1187_ (.A(\mux_bottom_track_27.INVTX1_0_.out ),
    .TE_B(_0350_),
    .Z(\mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1188_ (.A(net133),
    .TE_B(_0351_),
    .Z(\mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1189_ (.A(\mux_bottom_track_11.INVTX1_1_.out ),
    .TE_B(_0352_),
    .Z(\mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_4 _1190_ (.A(\mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0353_),
    .Z(\mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1191_ (.A(\mux_bottom_track_29.INVTX1_0_.out ),
    .TE_B(_0354_),
    .Z(\mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1192_ (.A(net134),
    .TE_B(_0355_),
    .Z(\mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1193_ (.A(\mux_bottom_track_11.INVTX1_2_.out ),
    .TE_B(_0356_),
    .Z(\mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_1 _1194_ (.A(\mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0357_),
    .Z(\mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1195_ (.A(\mux_bottom_track_31.INVTX1_0_.out ),
    .TE_B(_0358_),
    .Z(\mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1196_ (.A(net135),
    .TE_B(_0359_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1197_ (.A(\mux_bottom_track_13.INVTX1_2_.out ),
    .TE_B(_0360_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1198_ (.A(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0361_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_2 _1199_ (.A(\mux_bottom_track_33.INVTX1_0_.out ),
    .TE_B(_0362_),
    .Z(\mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1200_ (.A(net136),
    .TE_B(_0363_),
    .Z(\mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1201_ (.A(\mux_bottom_track_15.INVTX1_2_.out ),
    .TE_B(_0364_),
    .Z(\mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__ebufn_2 _1202_ (.A(\mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ),
    .TE_B(_0365_),
    .Z(\mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out ));
 sky130_fd_sc_hd__ebufn_1 _1203_ (.A(\mux_bottom_track_35.INVTX1_0_.out ),
    .TE_B(_0366_),
    .Z(\mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(ccff_head),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(chanx_right_in[0]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(chanx_right_in[10]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(chanx_right_in[11]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(chanx_right_in[12]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(chanx_right_in[13]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(chanx_right_in[14]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(chanx_right_in[15]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(chanx_right_in[16]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(chanx_right_in[17]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(chanx_right_in[18]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(chanx_right_in[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(chanx_right_in[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(chanx_right_in[3]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(chanx_right_in[4]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(chanx_right_in[5]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(chanx_right_in[6]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(chanx_right_in[7]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(chanx_right_in[8]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chanx_right_in[9]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(chany_bottom_in[0]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(chany_bottom_in[10]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(chany_bottom_in[11]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(chany_bottom_in[12]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(chany_bottom_in[13]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(chany_bottom_in[14]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chany_bottom_in[15]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(chany_bottom_in[16]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(chany_bottom_in[17]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(chany_bottom_in[18]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(chany_bottom_in[1]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(chany_bottom_in[2]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(chany_bottom_in[3]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(chany_bottom_in[4]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(chany_bottom_in[5]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(chany_bottom_in[6]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(chany_bottom_in[7]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(chany_bottom_in[8]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(chany_bottom_in[9]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(pReset),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(ccff_tail));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(chany_bottom_out[10]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(chany_bottom_out[11]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(chany_bottom_out[12]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(chany_bottom_out[13]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(chany_bottom_out[14]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(chany_bottom_out[15]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(chany_bottom_out[16]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(chany_bottom_out[17]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(chany_bottom_out[18]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(chany_bottom_out[9]));
 sky130_fd_sc_hd__conb_1 _1015__100 (.HI(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\mem_right_track_4.DFFR_1_.Q ));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
endmodule

