magic
tech sky130A
magscale 1 2
timestamp 1674237007
<< obsli1 >>
rect 1090 1959 560818 587337
<< obsm1 >>
rect 0 1712 560818 587448
<< metal2 >>
rect 13528 589000 13584 589600
rect 29628 589000 29684 589600
rect 46372 589000 46428 589600
rect 62472 589000 62528 589600
rect 79216 589000 79272 589600
rect 95316 589000 95372 589600
rect 112060 589000 112116 589600
rect 128160 589000 128216 589600
rect 144260 589000 144316 589600
rect 161004 589000 161060 589600
rect 177104 589000 177160 589600
rect 193848 589000 193904 589600
rect 209948 589000 210004 589600
rect 226048 589000 226104 589600
rect 242792 589000 242848 589600
rect 258892 589000 258948 589600
rect 275636 589000 275692 589600
rect 291736 589000 291792 589600
rect 308480 589000 308536 589600
rect 324580 589000 324636 589600
rect 340680 589000 340736 589600
rect 357424 589000 357480 589600
rect 373524 589000 373580 589600
rect 390268 589000 390324 589600
rect 406368 589000 406424 589600
rect 422468 589000 422524 589600
rect 439212 589000 439268 589600
rect 455312 589000 455368 589600
rect 472056 589000 472112 589600
rect 488156 589000 488212 589600
rect 504900 589000 504956 589600
rect 521000 589000 521056 589600
rect 537100 589000 537156 589600
rect 553844 589000 553900 589600
rect 4 0 60 600
rect 16104 0 16160 600
rect 32204 0 32260 600
rect 48948 0 49004 600
rect 65048 0 65104 600
rect 81792 0 81848 600
rect 97892 0 97948 600
rect 113992 0 114048 600
rect 130736 0 130792 600
rect 146836 0 146892 600
rect 163580 0 163636 600
rect 179680 0 179736 600
rect 195780 0 195836 600
rect 212524 0 212580 600
rect 228624 0 228680 600
rect 245368 0 245424 600
rect 261468 0 261524 600
rect 278212 0 278268 600
rect 294312 0 294368 600
rect 310412 0 310468 600
rect 327156 0 327212 600
rect 343256 0 343312 600
rect 360000 0 360056 600
rect 376100 0 376156 600
rect 392200 0 392256 600
rect 408944 0 409000 600
rect 425044 0 425100 600
rect 441788 0 441844 600
rect 457888 0 457944 600
rect 474632 0 474688 600
rect 490732 0 490788 600
rect 506832 0 506888 600
rect 523576 0 523632 600
rect 539676 0 539732 600
rect 556420 0 556476 600
<< obsm2 >>
rect 6 588944 13472 589000
rect 13640 588944 29572 589000
rect 29740 588944 46316 589000
rect 46484 588944 62416 589000
rect 62584 588944 79160 589000
rect 79328 588944 95260 589000
rect 95428 588944 112004 589000
rect 112172 588944 128104 589000
rect 128272 588944 144204 589000
rect 144372 588944 160948 589000
rect 161116 588944 177048 589000
rect 177216 588944 193792 589000
rect 193960 588944 209892 589000
rect 210060 588944 225992 589000
rect 226160 588944 242736 589000
rect 242904 588944 258836 589000
rect 259004 588944 275580 589000
rect 275748 588944 291680 589000
rect 291848 588944 308424 589000
rect 308592 588944 324524 589000
rect 324692 588944 340624 589000
rect 340792 588944 357368 589000
rect 357536 588944 373468 589000
rect 373636 588944 390212 589000
rect 390380 588944 406312 589000
rect 406480 588944 422412 589000
rect 422580 588944 439156 589000
rect 439324 588944 455256 589000
rect 455424 588944 472000 589000
rect 472168 588944 488100 589000
rect 488268 588944 504844 589000
rect 505012 588944 520944 589000
rect 521112 588944 537044 589000
rect 537212 588944 553788 589000
rect 553956 588944 560522 589000
rect 6 656 560522 588944
rect 116 534 16048 656
rect 16216 534 32148 656
rect 32316 534 48892 656
rect 49060 534 64992 656
rect 65160 534 81736 656
rect 81904 534 97836 656
rect 98004 534 113936 656
rect 114104 534 130680 656
rect 130848 534 146780 656
rect 146948 534 163524 656
rect 163692 534 179624 656
rect 179792 534 195724 656
rect 195892 534 212468 656
rect 212636 534 228568 656
rect 228736 534 245312 656
rect 245480 534 261412 656
rect 261580 534 278156 656
rect 278324 534 294256 656
rect 294424 534 310356 656
rect 310524 534 327100 656
rect 327268 534 343200 656
rect 343368 534 359944 656
rect 360112 534 376044 656
rect 376212 534 392144 656
rect 392312 534 408888 656
rect 409056 534 424988 656
rect 425156 534 441732 656
rect 441900 534 457832 656
rect 458000 534 474576 656
rect 474744 534 490676 656
rect 490844 534 506776 656
rect 506944 534 523520 656
rect 523688 534 539620 656
rect 539788 534 556364 656
rect 556532 534 560522 656
<< metal3 >>
rect 186 587328 786 587448
rect 561186 581208 561786 581328
rect 186 569648 786 569768
rect 561186 563528 561786 563648
rect 186 552648 786 552768
rect 561186 546528 561786 546648
rect 186 534968 786 535088
rect 561186 529528 561786 529648
rect 186 517968 786 518088
rect 561186 511848 561786 511968
rect 186 500968 786 501088
rect 561186 494848 561786 494968
rect 186 483288 786 483408
rect 561186 477168 561786 477288
rect 186 466288 786 466408
rect 561186 460168 561786 460288
rect 186 448608 786 448728
rect 561186 442488 561786 442608
rect 186 431608 786 431728
rect 561186 425488 561786 425608
rect 186 413928 786 414048
rect 561186 408488 561786 408608
rect 186 396928 786 397048
rect 561186 390808 561786 390928
rect 186 379928 786 380048
rect 561186 373808 561786 373928
rect 186 362248 786 362368
rect 561186 356128 561786 356248
rect 186 345248 786 345368
rect 561186 339128 561786 339248
rect 186 327568 786 327688
rect 561186 322128 561786 322248
rect 186 310568 786 310688
rect 561186 304448 561786 304568
rect 186 293568 786 293688
rect 561186 287448 561786 287568
rect 186 275888 786 276008
rect 561186 269768 561786 269888
rect 186 258888 786 259008
rect 561186 252768 561786 252888
rect 186 241208 786 241328
rect 561186 235088 561786 235208
rect 186 224208 786 224328
rect 561186 218088 561786 218208
rect 186 206528 786 206648
rect 561186 201088 561786 201208
rect 186 189528 786 189648
rect 561186 183408 561786 183528
rect 186 172528 786 172648
rect 561186 166408 561786 166528
rect 186 154848 786 154968
rect 561186 148728 561786 148848
rect 186 137848 786 137968
rect 561186 131728 561786 131848
rect 186 120168 786 120288
rect 561186 114728 561786 114848
rect 186 103168 786 103288
rect 561186 97048 561786 97168
rect 186 86168 786 86288
rect 561186 80048 561786 80168
rect 186 68488 786 68608
rect 561186 62368 561786 62488
rect 186 51488 786 51608
rect 561186 45368 561786 45488
rect 186 33808 786 33928
rect 561186 27688 561786 27808
rect 186 16808 786 16928
rect 561186 10688 561786 10808
<< obsm3 >>
rect 866 587248 561186 587421
rect 786 581408 561186 587248
rect 786 581128 561106 581408
rect 786 569848 561186 581128
rect 866 569568 561186 569848
rect 786 563728 561186 569568
rect 786 563448 561106 563728
rect 786 552848 561186 563448
rect 866 552568 561186 552848
rect 786 546728 561186 552568
rect 786 546448 561106 546728
rect 786 535168 561186 546448
rect 866 534888 561186 535168
rect 786 529728 561186 534888
rect 786 529448 561106 529728
rect 786 518168 561186 529448
rect 866 517888 561186 518168
rect 786 512048 561186 517888
rect 786 511768 561106 512048
rect 786 501168 561186 511768
rect 866 500888 561186 501168
rect 786 495048 561186 500888
rect 786 494768 561106 495048
rect 786 483488 561186 494768
rect 866 483208 561186 483488
rect 786 477368 561186 483208
rect 786 477088 561106 477368
rect 786 466488 561186 477088
rect 866 466208 561186 466488
rect 786 460368 561186 466208
rect 786 460088 561106 460368
rect 786 448808 561186 460088
rect 866 448528 561186 448808
rect 786 442688 561186 448528
rect 786 442408 561106 442688
rect 786 431808 561186 442408
rect 866 431528 561186 431808
rect 786 425688 561186 431528
rect 786 425408 561106 425688
rect 786 414128 561186 425408
rect 866 413848 561186 414128
rect 786 408688 561186 413848
rect 786 408408 561106 408688
rect 786 397128 561186 408408
rect 866 396848 561186 397128
rect 786 391008 561186 396848
rect 786 390728 561106 391008
rect 786 380128 561186 390728
rect 866 379848 561186 380128
rect 786 374008 561186 379848
rect 786 373728 561106 374008
rect 786 362448 561186 373728
rect 866 362168 561186 362448
rect 786 356328 561186 362168
rect 786 356048 561106 356328
rect 786 345448 561186 356048
rect 866 345168 561186 345448
rect 786 339328 561186 345168
rect 786 339048 561106 339328
rect 786 327768 561186 339048
rect 866 327488 561186 327768
rect 786 322328 561186 327488
rect 786 322048 561106 322328
rect 786 310768 561186 322048
rect 866 310488 561186 310768
rect 786 304648 561186 310488
rect 786 304368 561106 304648
rect 786 293768 561186 304368
rect 866 293488 561186 293768
rect 786 287648 561186 293488
rect 786 287368 561106 287648
rect 786 276088 561186 287368
rect 866 275808 561186 276088
rect 786 269968 561186 275808
rect 786 269688 561106 269968
rect 786 259088 561186 269688
rect 866 258808 561186 259088
rect 786 252968 561186 258808
rect 786 252688 561106 252968
rect 786 241408 561186 252688
rect 866 241128 561186 241408
rect 786 235288 561186 241128
rect 786 235008 561106 235288
rect 786 224408 561186 235008
rect 866 224128 561186 224408
rect 786 218288 561186 224128
rect 786 218008 561106 218288
rect 786 206728 561186 218008
rect 866 206448 561186 206728
rect 786 201288 561186 206448
rect 786 201008 561106 201288
rect 786 189728 561186 201008
rect 866 189448 561186 189728
rect 786 183608 561186 189448
rect 786 183328 561106 183608
rect 786 172728 561186 183328
rect 866 172448 561186 172728
rect 786 166608 561186 172448
rect 786 166328 561106 166608
rect 786 155048 561186 166328
rect 866 154768 561186 155048
rect 786 148928 561186 154768
rect 786 148648 561106 148928
rect 786 138048 561186 148648
rect 866 137768 561186 138048
rect 786 131928 561186 137768
rect 786 131648 561106 131928
rect 786 120368 561186 131648
rect 866 120088 561186 120368
rect 786 114928 561186 120088
rect 786 114648 561106 114928
rect 786 103368 561186 114648
rect 866 103088 561186 103368
rect 786 97248 561186 103088
rect 786 96968 561106 97248
rect 786 86368 561186 96968
rect 866 86088 561186 86368
rect 786 80248 561186 86088
rect 786 79968 561106 80248
rect 786 68688 561186 79968
rect 866 68408 561186 68688
rect 786 62568 561186 68408
rect 786 62288 561106 62568
rect 786 51688 561186 62288
rect 866 51408 561186 51688
rect 786 45568 561186 51408
rect 786 45288 561106 45568
rect 786 34008 561186 45288
rect 866 33728 561186 34008
rect 786 27888 561186 33728
rect 786 27608 561106 27888
rect 786 17008 561186 27608
rect 866 16728 561186 17008
rect 786 10888 561186 16728
rect 786 10608 561106 10888
rect 786 1943 561186 10608
<< metal4 >>
rect 2494 411016 2814 456808
rect 3230 411016 3550 456808
rect 2494 308744 2814 354536
rect 3230 308744 3550 354536
rect 2494 207016 2814 252808
rect 3230 207016 3550 252808
rect 2494 104744 2814 150536
rect 3230 104744 3550 150536
rect 8330 1928 8650 587368
rect 8990 1928 9310 587368
rect 17330 1928 17650 587368
rect 17990 1928 18310 587368
rect 26330 453444 26650 587368
rect 26330 351444 26650 413868
rect 26330 249444 26650 311868
rect 26330 147444 26650 209868
rect 26330 1928 26650 107868
rect 26990 1928 27310 587368
rect 35330 505089 35650 587368
rect 35990 505089 36310 587368
rect 44330 505089 44650 587368
rect 44990 505089 45310 587368
rect 53330 505089 53650 587368
rect 53990 505089 54310 587368
rect 35330 403089 35650 466359
rect 35990 403089 36310 466359
rect 44330 403089 44650 466359
rect 44990 403089 45310 466359
rect 53330 403089 53650 466359
rect 53990 403089 54310 466359
rect 62330 455444 62650 587368
rect 35330 301089 35650 364359
rect 35990 301089 36310 364359
rect 44330 301089 44650 364359
rect 44990 301089 45310 364359
rect 53330 301089 53650 364359
rect 53990 301089 54310 364359
rect 62330 353444 62650 415868
rect 35330 199089 35650 262359
rect 35990 199089 36310 262359
rect 44330 199089 44650 262359
rect 44990 199089 45310 262359
rect 53330 199089 53650 262359
rect 53990 199089 54310 262359
rect 62330 251444 62650 313868
rect 35330 70444 35650 160359
rect 35990 69953 36310 160359
rect 44330 69953 44650 160359
rect 44990 69953 45310 160359
rect 35330 1928 35650 30868
rect 35990 1928 36310 34079
rect 44330 1928 44650 34079
rect 44990 1928 45310 34079
rect 53330 1928 53650 160359
rect 53990 1928 54310 160359
rect 62330 149444 62650 211868
rect 62330 1928 62650 109868
rect 62990 1928 63310 587368
rect 71330 352681 71650 587368
rect 71990 352681 72310 587368
rect 80330 352681 80650 587368
rect 80990 352681 81310 587368
rect 89330 352681 89650 587368
rect 89990 352681 90310 587368
rect 71330 250681 71650 321567
rect 71990 250681 72310 321567
rect 80330 250681 80650 321567
rect 80990 250681 81310 321567
rect 89330 250681 89650 321567
rect 89990 250681 90310 321567
rect 71330 148681 71650 219567
rect 71990 148681 72310 219567
rect 80330 148681 80650 219567
rect 80990 148681 81310 219567
rect 89330 148681 89650 219567
rect 89990 148681 90310 219567
rect 71330 1928 71650 117567
rect 71990 1928 72310 117567
rect 80330 1928 80650 117567
rect 80990 1928 81310 117567
rect 89330 1928 89650 117567
rect 89990 1928 90310 117567
rect 98330 1928 98650 587368
rect 98990 1928 99310 587368
rect 107330 503865 107650 587368
rect 107990 503865 108310 587368
rect 116330 503865 116650 587368
rect 116990 503865 117310 587368
rect 125330 503865 125650 587368
rect 125990 503865 126310 587368
rect 134330 503865 134650 587368
rect 134990 503865 135310 587368
rect 143330 503865 143650 587368
rect 143990 561444 144310 587368
rect 143990 503865 144310 521868
rect 100934 413192 101254 458440
rect 101670 413192 101990 458440
rect 107330 454137 107650 466767
rect 107990 454137 108310 466767
rect 116330 454137 116650 466767
rect 116990 454137 117310 466767
rect 107330 401865 107650 419351
rect 107990 401865 108310 419351
rect 116330 401865 116650 419351
rect 116990 401865 117310 419351
rect 125330 401865 125650 466767
rect 125990 401865 126310 466767
rect 134330 401865 134650 466767
rect 134990 401865 135310 466767
rect 143330 401865 143650 466767
rect 143990 401865 144310 466767
rect 100934 310920 101254 356712
rect 101670 310920 101990 356712
rect 107330 299865 107650 364767
rect 107990 299865 108310 364767
rect 116330 351865 116650 364767
rect 116990 351865 117310 364767
rect 116330 299865 116650 330543
rect 116990 299865 117310 330543
rect 125330 299865 125650 364767
rect 125990 299865 126310 364767
rect 134330 299865 134650 364767
rect 134990 299865 135310 364767
rect 143330 299865 143650 364767
rect 143990 299865 144310 364767
rect 102406 209192 102726 254440
rect 103142 209192 103462 254440
rect 107330 197865 107650 262767
rect 107990 197865 108310 262767
rect 116330 249865 116650 262767
rect 116990 249865 117310 262767
rect 116330 197865 116650 228543
rect 116990 197865 117310 228543
rect 125330 197865 125650 262767
rect 125990 197865 126310 262767
rect 134330 197865 134650 262767
rect 134990 197865 135310 262767
rect 143330 197865 143650 262767
rect 143990 197865 144310 262767
rect 100934 106920 101254 152712
rect 101670 106920 101990 152712
rect 107330 93865 107650 160767
rect 107990 93865 108310 160767
rect 116330 147865 116650 160767
rect 116990 147865 117310 160767
rect 116330 93865 116650 126543
rect 116990 93865 117310 126543
rect 125330 93865 125650 160767
rect 125990 93865 126310 160767
rect 107330 1928 107650 56359
rect 107990 1928 108310 56359
rect 116330 1928 116650 56359
rect 116990 1928 117310 56359
rect 125330 1928 125650 56359
rect 125990 1928 126310 56359
rect 134330 1928 134650 160767
rect 134990 1928 135310 160767
rect 143330 1928 143650 160767
rect 143990 45444 144310 160767
rect 143990 1928 144310 5868
rect 152330 1928 152650 587368
rect 152990 1928 153310 587368
rect 161330 457089 161650 587368
rect 161990 457089 162310 587368
rect 170330 457089 170650 587368
rect 170990 457089 171310 587368
rect 179330 457089 179650 587368
rect 179990 457089 180310 587368
rect 161330 354409 161650 418903
rect 161990 354409 162310 418903
rect 170330 354409 170650 418903
rect 170990 354409 171310 418903
rect 179330 354409 179650 418903
rect 179990 354409 180310 418903
rect 161330 252409 161650 314999
rect 161990 252409 162310 314999
rect 170330 252409 170650 314999
rect 170990 252409 171310 314999
rect 179330 252409 179650 314999
rect 179990 252409 180310 314999
rect 161330 150409 161650 212999
rect 161990 150409 162310 212999
rect 170330 150409 170650 212999
rect 170990 150409 171310 212999
rect 179330 150409 179650 212999
rect 179990 150409 180310 212999
rect 161330 1928 161650 110999
rect 161990 1928 162310 110999
rect 170330 95225 170650 110999
rect 170990 95225 171310 110999
rect 179330 95225 179650 110999
rect 179990 95225 180310 110999
rect 188330 95225 188650 587368
rect 188990 95225 189310 587368
rect 170330 1928 170650 56359
rect 170990 1928 171310 56359
rect 179330 1928 179650 56359
rect 179990 1928 180310 56359
rect 188330 1928 188650 56359
rect 188990 1928 189310 56359
rect 197330 1928 197650 587368
rect 197990 1928 198310 587368
rect 199742 462696 200062 508488
rect 206330 503865 206650 587368
rect 206990 503865 207310 587368
rect 215330 561444 215650 587368
rect 215330 503865 215650 521868
rect 215990 503865 216310 587368
rect 224330 503865 224650 587368
rect 224990 503865 225310 587368
rect 233330 503865 233650 587368
rect 233990 503865 234310 587368
rect 242330 503865 242650 587368
rect 242990 503865 243310 587368
rect 201398 414824 201718 458440
rect 199742 361512 200062 406216
rect 206330 401865 206650 466767
rect 206990 454137 207310 466767
rect 215330 454137 215650 466767
rect 215990 454137 216310 466767
rect 224330 454137 224650 466767
rect 206990 401865 207310 419351
rect 215330 401865 215650 419351
rect 215990 401865 216310 419351
rect 224330 401865 224650 419351
rect 224990 401865 225310 466767
rect 233330 401865 233650 466767
rect 233990 401865 234310 466767
rect 242330 401865 242650 466767
rect 242990 401865 243310 466767
rect 201398 313640 201718 356168
rect 199742 259240 200062 303944
rect 206330 299865 206650 364767
rect 206990 299865 207310 364767
rect 215330 351865 215650 364767
rect 215990 351865 216310 364767
rect 215330 299865 215650 330543
rect 215990 299865 216310 330543
rect 224330 299865 224650 364767
rect 224990 299865 225310 364767
rect 233330 299865 233650 364767
rect 233990 299865 234310 364767
rect 242330 299865 242650 364767
rect 242990 299865 243310 364767
rect 201398 211368 201718 253896
rect 199742 156968 200062 202760
rect 206330 197865 206650 262767
rect 206990 197865 207310 262767
rect 215330 249865 215650 262767
rect 215990 249865 216310 262767
rect 215330 197865 215650 228543
rect 215990 197865 216310 228543
rect 224330 197865 224650 262767
rect 224990 197865 225310 262767
rect 233330 197865 233650 262767
rect 233990 197865 234310 262767
rect 242330 197865 242650 262767
rect 242990 197865 243310 262767
rect 201398 109096 201718 152712
rect 201398 53608 201718 98312
rect 206330 1928 206650 160767
rect 206990 1928 207310 160767
rect 215330 147865 215650 160767
rect 215990 147865 216310 160767
rect 215330 93865 215650 126543
rect 215990 93865 216310 126543
rect 224330 93865 224650 160767
rect 224990 93865 225310 160767
rect 215330 45444 215650 56359
rect 215330 1928 215650 5868
rect 215990 1928 216310 56359
rect 224330 1928 224650 56359
rect 224990 1928 225310 56359
rect 233330 1928 233650 160767
rect 233990 1928 234310 160767
rect 242330 1928 242650 160767
rect 242990 1928 243310 160767
rect 251330 1928 251650 587368
rect 251990 1928 252310 587368
rect 260330 457089 260650 587368
rect 260990 457089 261310 587368
rect 269330 457089 269650 587368
rect 269990 457089 270310 587368
rect 278330 457089 278650 587368
rect 278990 457089 279310 587368
rect 260330 354409 260650 418903
rect 260990 354409 261310 418903
rect 269330 354409 269650 418903
rect 269990 354409 270310 418903
rect 278330 354409 278650 418903
rect 278990 354409 279310 418903
rect 287330 354409 287650 587368
rect 260330 252409 260650 314999
rect 260990 252409 261310 314999
rect 269330 252409 269650 314999
rect 269990 252409 270310 314999
rect 278330 252409 278650 314999
rect 278990 252409 279310 314999
rect 287330 252409 287650 314999
rect 260330 150409 260650 212999
rect 260990 150409 261310 212999
rect 269330 150409 269650 212999
rect 269990 150409 270310 212999
rect 278330 150409 278650 212999
rect 278990 150409 279310 212999
rect 287330 150409 287650 212999
rect 260330 1928 260650 110999
rect 260990 1928 261310 110999
rect 269330 95225 269650 110999
rect 269990 95225 270310 110999
rect 278330 95225 278650 110999
rect 278990 95225 279310 110999
rect 287330 95225 287650 110999
rect 287990 95225 288310 587368
rect 296330 95225 296650 587368
rect 296990 95225 297310 587368
rect 301494 462696 301814 508488
rect 302230 462696 302550 508488
rect 301494 360968 301814 406760
rect 302230 360968 302550 406760
rect 301494 258696 301814 304488
rect 302230 258696 302550 304488
rect 301494 156968 301814 202760
rect 302230 156968 302550 202760
rect 269330 1928 269650 56359
rect 269990 1928 270310 56359
rect 278330 1928 278650 56359
rect 278990 1928 279310 56359
rect 287330 1928 287650 56359
rect 287990 1928 288310 56359
rect 296330 1928 296650 56359
rect 296990 1928 297310 56359
rect 305330 1928 305650 587368
rect 305990 503865 306310 587368
rect 314330 503865 314650 587368
rect 314990 503865 315310 587368
rect 323330 503865 323650 587368
rect 323990 503865 324310 587368
rect 332330 561444 332650 587368
rect 332330 503865 332650 521868
rect 332990 503865 333310 587368
rect 341330 503865 341650 587368
rect 341990 503865 342310 587368
rect 305990 401865 306310 466767
rect 314330 454137 314650 466767
rect 314990 454137 315310 466767
rect 323330 454137 323650 466767
rect 323990 454137 324310 466767
rect 314330 401865 314650 419351
rect 314990 401865 315310 419351
rect 323330 401865 323650 419351
rect 323990 401865 324310 419351
rect 332330 401865 332650 466767
rect 332990 401865 333310 466767
rect 341330 401865 341650 466767
rect 341990 401865 342310 466767
rect 305990 299865 306310 364767
rect 314330 351865 314650 364767
rect 314990 351865 315310 364767
rect 314330 299865 314650 330543
rect 314990 299865 315310 330543
rect 323330 299865 323650 364767
rect 323990 299865 324310 364767
rect 332330 299865 332650 364767
rect 332990 299865 333310 364767
rect 341330 299865 341650 364767
rect 341990 299865 342310 364767
rect 305990 197865 306310 262767
rect 314330 249865 314650 262767
rect 314990 249865 315310 262767
rect 314330 197865 314650 228543
rect 314990 197865 315310 228543
rect 323330 197865 323650 262767
rect 323990 197865 324310 262767
rect 332330 197865 332650 262767
rect 332990 197865 333310 262767
rect 341330 197865 341650 262767
rect 341990 197865 342310 262767
rect 305990 1928 306310 160767
rect 314330 149865 314650 160767
rect 314990 149865 315310 160767
rect 314330 93865 314650 128543
rect 314990 93865 315310 128543
rect 323330 93865 323650 160767
rect 323990 93865 324310 160767
rect 314330 1928 314650 56359
rect 314990 1928 315310 56359
rect 323330 1928 323650 56359
rect 323990 1928 324310 56359
rect 332330 45444 332650 160767
rect 332330 1928 332650 5868
rect 332990 1928 333310 160767
rect 341330 1928 341650 160767
rect 341990 1928 342310 160767
rect 350330 1928 350650 587368
rect 350990 1928 351310 587368
rect 354486 462696 354806 508488
rect 355222 462696 355542 508488
rect 354486 360968 354806 406760
rect 355222 360968 355542 406760
rect 359330 354409 359650 587368
rect 359990 457089 360310 587368
rect 368330 457089 368650 587368
rect 368990 457089 369310 587368
rect 377330 457089 377650 587368
rect 377990 457089 378310 587368
rect 386330 457089 386650 587368
rect 386990 457089 387310 587368
rect 359990 354409 360310 418903
rect 368330 354409 368650 418903
rect 368990 354409 369310 418903
rect 377330 354409 377650 418903
rect 377990 354409 378310 418903
rect 386330 354409 386650 418903
rect 386990 354409 387310 418903
rect 354486 258696 354806 304488
rect 355222 258696 355542 304488
rect 359330 252409 359650 314999
rect 359990 252409 360310 314999
rect 368330 252409 368650 314999
rect 368990 252409 369310 314999
rect 377330 252409 377650 314999
rect 377990 252409 378310 314999
rect 386330 252409 386650 314999
rect 386990 252409 387310 314999
rect 354486 156968 354806 202760
rect 355222 156968 355542 202760
rect 359330 150409 359650 212999
rect 359990 150409 360310 212999
rect 368330 150409 368650 212999
rect 368990 150409 369310 212999
rect 377330 150409 377650 212999
rect 377990 150409 378310 212999
rect 386330 150409 386650 212999
rect 386990 150409 387310 212999
rect 354302 53608 354622 98312
rect 359330 1928 359650 110999
rect 359990 1928 360310 110999
rect 368330 95225 368650 110999
rect 368990 95225 369310 110999
rect 377330 95225 377650 110999
rect 377990 95225 378310 110999
rect 386330 95225 386650 110999
rect 386990 95225 387310 110999
rect 395330 95225 395650 587368
rect 395990 95225 396310 587368
rect 368330 1928 368650 56359
rect 368990 1928 369310 56359
rect 377330 1928 377650 56359
rect 377990 1928 378310 56359
rect 386330 1928 386650 56359
rect 386990 1928 387310 56359
rect 395330 1928 395650 56359
rect 395990 1928 396310 56359
rect 404330 1928 404650 587368
rect 404990 1928 405310 587368
rect 413330 503865 413650 587368
rect 413990 503865 414310 587368
rect 422330 503865 422650 587368
rect 422990 503865 423310 587368
rect 431330 503865 431650 587368
rect 431990 503865 432310 587368
rect 440330 503865 440650 587368
rect 440990 503865 441310 587368
rect 449330 503865 449650 587368
rect 449990 561444 450310 587368
rect 449990 503865 450310 521868
rect 413330 454137 413650 466767
rect 413990 454137 414310 466767
rect 422330 454137 422650 466767
rect 422990 454137 423310 466767
rect 413330 401865 413650 419351
rect 413990 401865 414310 419351
rect 422330 401865 422650 419351
rect 422990 401865 423310 419351
rect 431330 401865 431650 466767
rect 431990 401865 432310 466767
rect 440330 401865 440650 466767
rect 440990 401865 441310 466767
rect 449330 401865 449650 466767
rect 449990 401865 450310 466767
rect 455502 462696 455822 501416
rect 456238 462696 456558 501416
rect 454398 456168 454718 458440
rect 413330 299865 413650 364767
rect 413990 299865 414310 364767
rect 422330 351865 422650 364767
rect 422990 351865 423310 364767
rect 422330 299865 422650 330543
rect 422990 299865 423310 330543
rect 431330 299865 431650 364767
rect 431990 299865 432310 364767
rect 440330 299865 440650 364767
rect 440990 299865 441310 364767
rect 449330 299865 449650 364767
rect 449990 299865 450310 364767
rect 455502 360968 455822 399688
rect 456238 360968 456558 399688
rect 454030 353896 454350 356712
rect 454766 353896 455086 356712
rect 413330 197865 413650 262767
rect 413990 197865 414310 262767
rect 422330 250465 422650 262767
rect 422990 250465 423310 262767
rect 422330 197865 422650 229143
rect 422990 197865 423310 229143
rect 431330 197865 431650 262767
rect 431990 197865 432310 262767
rect 440330 197865 440650 262767
rect 440990 197865 441310 262767
rect 449330 197865 449650 262767
rect 449990 197865 450310 262767
rect 455502 258696 455822 297416
rect 456238 258696 456558 297416
rect 454030 252168 454350 255528
rect 454766 252168 455086 255528
rect 413330 93865 413650 160767
rect 413990 93865 414310 160767
rect 422330 147865 422650 160767
rect 422990 147865 423310 160767
rect 422330 93865 422650 126543
rect 422990 93865 423310 126543
rect 431330 93865 431650 160767
rect 431990 93865 432310 160767
rect 413330 1928 413650 56359
rect 413990 1928 414310 56359
rect 422330 1928 422650 56359
rect 422990 1928 423310 56359
rect 431330 1928 431650 56359
rect 431990 1928 432310 56359
rect 440330 1928 440650 160767
rect 440990 1928 441310 160767
rect 449330 1928 449650 160767
rect 449990 45444 450310 160767
rect 455502 156968 455822 195688
rect 456238 156968 456558 195688
rect 454030 149896 454350 152712
rect 454766 149896 455086 152712
rect 449990 1928 450310 5868
rect 458330 1928 458650 587368
rect 458990 1928 459310 587368
rect 467330 80537 467650 587368
rect 467990 80537 468310 587368
rect 476330 492649 476650 587368
rect 476990 492649 477310 587368
rect 485330 492649 485650 587368
rect 485990 492649 486310 587368
rect 476330 441649 476650 461399
rect 476990 441649 477310 461399
rect 485330 441649 485650 461399
rect 485990 441649 486310 461399
rect 476330 390649 476650 409719
rect 476990 390649 477310 409719
rect 485330 390649 485650 409719
rect 485990 390649 486310 409719
rect 476330 333665 476650 359399
rect 476990 333665 477310 359399
rect 485330 333665 485650 359399
rect 485990 333665 486310 359399
rect 494330 333665 494650 587368
rect 494990 498444 495310 587368
rect 494990 396444 495310 458868
rect 494990 333665 495310 356868
rect 476330 288649 476650 305951
rect 476990 288649 477310 305951
rect 485330 288649 485650 305951
rect 485990 288649 486310 305951
rect 476330 231665 476650 257399
rect 476990 231665 477310 257399
rect 485330 231665 485650 257399
rect 485990 231665 486310 257399
rect 494330 231665 494650 305951
rect 494990 294444 495310 305951
rect 494990 231665 495310 254868
rect 476330 186649 476650 203951
rect 476990 186649 477310 203951
rect 485330 186649 485650 203951
rect 485990 186649 486310 203951
rect 476330 129665 476650 155399
rect 476990 129665 477310 155399
rect 485330 129665 485650 155399
rect 485990 129665 486310 155399
rect 494330 129665 494650 203951
rect 494990 192444 495310 203951
rect 494990 129665 495310 152868
rect 476330 80537 476650 101951
rect 476990 80537 477310 101951
rect 467330 1928 467650 56087
rect 467990 1928 468310 56087
rect 476330 1928 476650 56087
rect 476990 1928 477310 56087
rect 485330 1928 485650 101951
rect 485990 1928 486310 101951
rect 494330 1928 494650 101951
rect 494990 1928 495310 101951
rect 503330 1928 503650 587368
rect 503990 1928 504310 587368
rect 512330 1928 512650 587368
rect 512990 1928 513310 587368
rect 521330 1928 521650 587368
rect 521990 1928 522310 587368
rect 530330 1928 530650 587368
rect 530990 1928 531310 587368
rect 539330 1928 539650 587368
rect 539990 1928 540310 587368
rect 548330 1928 548650 587368
rect 548990 501444 549310 587368
rect 548990 399444 549310 461868
rect 548990 297444 549310 359868
rect 548990 195444 549310 257868
rect 548990 1928 549310 155868
rect 557330 1928 557650 587368
rect 557990 1928 558310 587368
<< obsm4 >>
rect 5197 2147 8250 587149
rect 8730 2147 8910 587149
rect 9390 2147 17250 587149
rect 17730 2147 17910 587149
rect 18390 453364 26250 587149
rect 26730 453364 26910 587149
rect 18390 413948 26910 453364
rect 18390 351364 26250 413948
rect 26730 351364 26910 413948
rect 18390 311948 26910 351364
rect 18390 249364 26250 311948
rect 26730 249364 26910 311948
rect 18390 209948 26910 249364
rect 18390 147364 26250 209948
rect 26730 147364 26910 209948
rect 18390 107948 26910 147364
rect 18390 2147 26250 107948
rect 26730 2147 26910 107948
rect 27390 505009 35250 587149
rect 35730 505009 35910 587149
rect 36390 505009 44250 587149
rect 44730 505009 44910 587149
rect 45390 505009 53250 587149
rect 53730 505009 53910 587149
rect 54390 505009 62250 587149
rect 27390 466439 62250 505009
rect 27390 403009 35250 466439
rect 35730 403009 35910 466439
rect 36390 403009 44250 466439
rect 44730 403009 44910 466439
rect 45390 403009 53250 466439
rect 53730 403009 53910 466439
rect 54390 455364 62250 466439
rect 62730 455364 62910 587149
rect 54390 415948 62910 455364
rect 54390 403009 62250 415948
rect 27390 364439 62250 403009
rect 27390 301009 35250 364439
rect 35730 301009 35910 364439
rect 36390 301009 44250 364439
rect 44730 301009 44910 364439
rect 45390 301009 53250 364439
rect 53730 301009 53910 364439
rect 54390 353364 62250 364439
rect 62730 353364 62910 415948
rect 54390 313948 62910 353364
rect 54390 301009 62250 313948
rect 27390 262439 62250 301009
rect 27390 199009 35250 262439
rect 35730 199009 35910 262439
rect 36390 199009 44250 262439
rect 44730 199009 44910 262439
rect 45390 199009 53250 262439
rect 53730 199009 53910 262439
rect 54390 251364 62250 262439
rect 62730 251364 62910 313948
rect 54390 211948 62910 251364
rect 54390 199009 62250 211948
rect 27390 160439 62250 199009
rect 27390 70364 35250 160439
rect 35730 70364 35910 160439
rect 27390 69873 35910 70364
rect 36390 69873 44250 160439
rect 44730 69873 44910 160439
rect 45390 69873 53250 160439
rect 27390 34159 53250 69873
rect 27390 30948 35910 34159
rect 27390 2147 35250 30948
rect 35730 2147 35910 30948
rect 36390 2147 44250 34159
rect 44730 2147 44910 34159
rect 45390 2147 53250 34159
rect 53730 2147 53910 160439
rect 54390 149364 62250 160439
rect 62730 149364 62910 211948
rect 54390 109948 62910 149364
rect 54390 2147 62250 109948
rect 62730 2147 62910 109948
rect 63390 352601 71250 587149
rect 71730 352601 71910 587149
rect 72390 352601 80250 587149
rect 80730 352601 80910 587149
rect 81390 352601 89250 587149
rect 89730 352601 89910 587149
rect 90390 352601 98250 587149
rect 63390 321647 98250 352601
rect 63390 250601 71250 321647
rect 71730 250601 71910 321647
rect 72390 250601 80250 321647
rect 80730 250601 80910 321647
rect 81390 250601 89250 321647
rect 89730 250601 89910 321647
rect 90390 250601 98250 321647
rect 63390 219647 98250 250601
rect 63390 148601 71250 219647
rect 71730 148601 71910 219647
rect 72390 148601 80250 219647
rect 80730 148601 80910 219647
rect 81390 148601 89250 219647
rect 89730 148601 89910 219647
rect 90390 148601 98250 219647
rect 63390 117647 98250 148601
rect 63390 2147 71250 117647
rect 71730 2147 71910 117647
rect 72390 2147 80250 117647
rect 80730 2147 80910 117647
rect 81390 2147 89250 117647
rect 89730 2147 89910 117647
rect 90390 2147 98250 117647
rect 98730 2147 98910 587149
rect 99390 503785 107250 587149
rect 107730 503785 107910 587149
rect 108390 503785 116250 587149
rect 116730 503785 116910 587149
rect 117390 503785 125250 587149
rect 125730 503785 125910 587149
rect 126390 503785 134250 587149
rect 134730 503785 134910 587149
rect 135390 503785 143250 587149
rect 143730 561364 143910 587149
rect 144390 561364 152250 587149
rect 143730 521948 152250 561364
rect 143730 503785 143910 521948
rect 144390 503785 152250 521948
rect 99390 466847 152250 503785
rect 99390 458520 107250 466847
rect 99390 413112 100854 458520
rect 101334 413112 101590 458520
rect 102070 454057 107250 458520
rect 107730 454057 107910 466847
rect 108390 454057 116250 466847
rect 116730 454057 116910 466847
rect 117390 454057 125250 466847
rect 102070 419431 125250 454057
rect 102070 413112 107250 419431
rect 99390 401785 107250 413112
rect 107730 401785 107910 419431
rect 108390 401785 116250 419431
rect 116730 401785 116910 419431
rect 117390 401785 125250 419431
rect 125730 401785 125910 466847
rect 126390 401785 134250 466847
rect 134730 401785 134910 466847
rect 135390 401785 143250 466847
rect 143730 401785 143910 466847
rect 144390 401785 152250 466847
rect 99390 364847 152250 401785
rect 99390 356792 107250 364847
rect 99390 310840 100854 356792
rect 101334 310840 101590 356792
rect 102070 310840 107250 356792
rect 99390 299785 107250 310840
rect 107730 299785 107910 364847
rect 108390 351785 116250 364847
rect 116730 351785 116910 364847
rect 117390 351785 125250 364847
rect 108390 330623 125250 351785
rect 108390 299785 116250 330623
rect 116730 299785 116910 330623
rect 117390 299785 125250 330623
rect 125730 299785 125910 364847
rect 126390 299785 134250 364847
rect 134730 299785 134910 364847
rect 135390 299785 143250 364847
rect 143730 299785 143910 364847
rect 144390 299785 152250 364847
rect 99390 262847 152250 299785
rect 99390 254520 107250 262847
rect 99390 209112 102326 254520
rect 102806 209112 103062 254520
rect 103542 209112 107250 254520
rect 99390 197785 107250 209112
rect 107730 197785 107910 262847
rect 108390 249785 116250 262847
rect 116730 249785 116910 262847
rect 117390 249785 125250 262847
rect 108390 228623 125250 249785
rect 108390 197785 116250 228623
rect 116730 197785 116910 228623
rect 117390 197785 125250 228623
rect 125730 197785 125910 262847
rect 126390 197785 134250 262847
rect 134730 197785 134910 262847
rect 135390 197785 143250 262847
rect 143730 197785 143910 262847
rect 144390 197785 152250 262847
rect 99390 160847 152250 197785
rect 99390 152792 107250 160847
rect 99390 106840 100854 152792
rect 101334 106840 101590 152792
rect 102070 106840 107250 152792
rect 99390 93785 107250 106840
rect 107730 93785 107910 160847
rect 108390 147785 116250 160847
rect 116730 147785 116910 160847
rect 117390 147785 125250 160847
rect 108390 126623 125250 147785
rect 108390 93785 116250 126623
rect 116730 93785 116910 126623
rect 117390 93785 125250 126623
rect 125730 93785 125910 160847
rect 126390 93785 134250 160847
rect 99390 56439 134250 93785
rect 99390 2147 107250 56439
rect 107730 2147 107910 56439
rect 108390 2147 116250 56439
rect 116730 2147 116910 56439
rect 117390 2147 125250 56439
rect 125730 2147 125910 56439
rect 126390 2147 134250 56439
rect 134730 2147 134910 160847
rect 135390 2147 143250 160847
rect 143730 45364 143910 160847
rect 144390 45364 152250 160847
rect 143730 5948 152250 45364
rect 143730 2147 143910 5948
rect 144390 2147 152250 5948
rect 152730 2147 152910 587149
rect 153390 457009 161250 587149
rect 161730 457009 161910 587149
rect 162390 457009 170250 587149
rect 170730 457009 170910 587149
rect 171390 457009 179250 587149
rect 179730 457009 179910 587149
rect 180390 457009 188250 587149
rect 153390 418983 188250 457009
rect 153390 354329 161250 418983
rect 161730 354329 161910 418983
rect 162390 354329 170250 418983
rect 170730 354329 170910 418983
rect 171390 354329 179250 418983
rect 179730 354329 179910 418983
rect 180390 354329 188250 418983
rect 153390 315079 188250 354329
rect 153390 252329 161250 315079
rect 161730 252329 161910 315079
rect 162390 252329 170250 315079
rect 170730 252329 170910 315079
rect 171390 252329 179250 315079
rect 179730 252329 179910 315079
rect 180390 252329 188250 315079
rect 153390 213079 188250 252329
rect 153390 150329 161250 213079
rect 161730 150329 161910 213079
rect 162390 150329 170250 213079
rect 170730 150329 170910 213079
rect 171390 150329 179250 213079
rect 179730 150329 179910 213079
rect 180390 150329 188250 213079
rect 153390 111079 188250 150329
rect 153390 2147 161250 111079
rect 161730 2147 161910 111079
rect 162390 95145 170250 111079
rect 170730 95145 170910 111079
rect 171390 95145 179250 111079
rect 179730 95145 179910 111079
rect 180390 95145 188250 111079
rect 188730 95145 188910 587149
rect 189390 95145 197250 587149
rect 162390 56439 197250 95145
rect 162390 2147 170250 56439
rect 170730 2147 170910 56439
rect 171390 2147 179250 56439
rect 179730 2147 179910 56439
rect 180390 2147 188250 56439
rect 188730 2147 188910 56439
rect 189390 2147 197250 56439
rect 197730 2147 197910 587149
rect 198390 508568 206250 587149
rect 198390 462616 199662 508568
rect 200142 503785 206250 508568
rect 206730 503785 206910 587149
rect 207390 561364 215250 587149
rect 215730 561364 215910 587149
rect 207390 521948 215910 561364
rect 207390 503785 215250 521948
rect 215730 503785 215910 521948
rect 216390 503785 224250 587149
rect 224730 503785 224910 587149
rect 225390 503785 233250 587149
rect 233730 503785 233910 587149
rect 234390 503785 242250 587149
rect 242730 503785 242910 587149
rect 243390 503785 251250 587149
rect 200142 466847 251250 503785
rect 200142 462616 206250 466847
rect 198390 458520 206250 462616
rect 198390 414744 201318 458520
rect 201798 414744 206250 458520
rect 198390 406296 206250 414744
rect 198390 361432 199662 406296
rect 200142 401785 206250 406296
rect 206730 454057 206910 466847
rect 207390 454057 215250 466847
rect 215730 454057 215910 466847
rect 216390 454057 224250 466847
rect 224730 454057 224910 466847
rect 206730 419431 224910 454057
rect 206730 401785 206910 419431
rect 207390 401785 215250 419431
rect 215730 401785 215910 419431
rect 216390 401785 224250 419431
rect 224730 401785 224910 419431
rect 225390 401785 233250 466847
rect 233730 401785 233910 466847
rect 234390 401785 242250 466847
rect 242730 401785 242910 466847
rect 243390 401785 251250 466847
rect 200142 364847 251250 401785
rect 200142 361432 206250 364847
rect 198390 356248 206250 361432
rect 198390 313560 201318 356248
rect 201798 313560 206250 356248
rect 198390 304024 206250 313560
rect 198390 259160 199662 304024
rect 200142 299785 206250 304024
rect 206730 299785 206910 364847
rect 207390 351785 215250 364847
rect 215730 351785 215910 364847
rect 216390 351785 224250 364847
rect 207390 330623 224250 351785
rect 207390 299785 215250 330623
rect 215730 299785 215910 330623
rect 216390 299785 224250 330623
rect 224730 299785 224910 364847
rect 225390 299785 233250 364847
rect 233730 299785 233910 364847
rect 234390 299785 242250 364847
rect 242730 299785 242910 364847
rect 243390 299785 251250 364847
rect 200142 262847 251250 299785
rect 200142 259160 206250 262847
rect 198390 253976 206250 259160
rect 198390 211288 201318 253976
rect 201798 211288 206250 253976
rect 198390 202840 206250 211288
rect 198390 156888 199662 202840
rect 200142 197785 206250 202840
rect 206730 197785 206910 262847
rect 207390 249785 215250 262847
rect 215730 249785 215910 262847
rect 216390 249785 224250 262847
rect 207390 228623 224250 249785
rect 207390 197785 215250 228623
rect 215730 197785 215910 228623
rect 216390 197785 224250 228623
rect 224730 197785 224910 262847
rect 225390 197785 233250 262847
rect 233730 197785 233910 262847
rect 234390 197785 242250 262847
rect 242730 197785 242910 262847
rect 243390 197785 251250 262847
rect 200142 160847 251250 197785
rect 200142 156888 206250 160847
rect 198390 152792 206250 156888
rect 198390 109016 201318 152792
rect 201798 109016 206250 152792
rect 198390 98392 206250 109016
rect 198390 53528 201318 98392
rect 201798 53528 206250 98392
rect 198390 2147 206250 53528
rect 206730 2147 206910 160847
rect 207390 147785 215250 160847
rect 215730 147785 215910 160847
rect 216390 147785 224250 160847
rect 207390 126623 224250 147785
rect 207390 93785 215250 126623
rect 215730 93785 215910 126623
rect 216390 93785 224250 126623
rect 224730 93785 224910 160847
rect 225390 93785 233250 160847
rect 207390 56439 233250 93785
rect 207390 45364 215250 56439
rect 215730 45364 215910 56439
rect 207390 5948 215910 45364
rect 207390 2147 215250 5948
rect 215730 2147 215910 5948
rect 216390 2147 224250 56439
rect 224730 2147 224910 56439
rect 225390 2147 233250 56439
rect 233730 2147 233910 160847
rect 234390 2147 242250 160847
rect 242730 2147 242910 160847
rect 243390 2147 251250 160847
rect 251730 2147 251910 587149
rect 252390 457009 260250 587149
rect 260730 457009 260910 587149
rect 261390 457009 269250 587149
rect 269730 457009 269910 587149
rect 270390 457009 278250 587149
rect 278730 457009 278910 587149
rect 279390 457009 287250 587149
rect 252390 418983 287250 457009
rect 252390 354329 260250 418983
rect 260730 354329 260910 418983
rect 261390 354329 269250 418983
rect 269730 354329 269910 418983
rect 270390 354329 278250 418983
rect 278730 354329 278910 418983
rect 279390 354329 287250 418983
rect 287730 354329 287910 587149
rect 252390 315079 287910 354329
rect 252390 252329 260250 315079
rect 260730 252329 260910 315079
rect 261390 252329 269250 315079
rect 269730 252329 269910 315079
rect 270390 252329 278250 315079
rect 278730 252329 278910 315079
rect 279390 252329 287250 315079
rect 287730 252329 287910 315079
rect 252390 213079 287910 252329
rect 252390 150329 260250 213079
rect 260730 150329 260910 213079
rect 261390 150329 269250 213079
rect 269730 150329 269910 213079
rect 270390 150329 278250 213079
rect 278730 150329 278910 213079
rect 279390 150329 287250 213079
rect 287730 150329 287910 213079
rect 252390 111079 287910 150329
rect 252390 2147 260250 111079
rect 260730 2147 260910 111079
rect 261390 95145 269250 111079
rect 269730 95145 269910 111079
rect 270390 95145 278250 111079
rect 278730 95145 278910 111079
rect 279390 95145 287250 111079
rect 287730 95145 287910 111079
rect 288390 95145 296250 587149
rect 296730 95145 296910 587149
rect 297390 508568 305250 587149
rect 297390 462616 301414 508568
rect 301894 462616 302150 508568
rect 302630 462616 305250 508568
rect 297390 406840 305250 462616
rect 297390 360888 301414 406840
rect 301894 360888 302150 406840
rect 302630 360888 305250 406840
rect 297390 304568 305250 360888
rect 297390 258616 301414 304568
rect 301894 258616 302150 304568
rect 302630 258616 305250 304568
rect 297390 202840 305250 258616
rect 297390 156888 301414 202840
rect 301894 156888 302150 202840
rect 302630 156888 305250 202840
rect 297390 95145 305250 156888
rect 261390 56439 305250 95145
rect 261390 2147 269250 56439
rect 269730 2147 269910 56439
rect 270390 2147 278250 56439
rect 278730 2147 278910 56439
rect 279390 2147 287250 56439
rect 287730 2147 287910 56439
rect 288390 2147 296250 56439
rect 296730 2147 296910 56439
rect 297390 2147 305250 56439
rect 305730 503785 305910 587149
rect 306390 503785 314250 587149
rect 314730 503785 314910 587149
rect 315390 503785 323250 587149
rect 323730 503785 323910 587149
rect 324390 561364 332250 587149
rect 332730 561364 332910 587149
rect 324390 521948 332910 561364
rect 324390 503785 332250 521948
rect 332730 503785 332910 521948
rect 333390 503785 341250 587149
rect 341730 503785 341910 587149
rect 342390 503785 350250 587149
rect 305730 466847 350250 503785
rect 305730 401785 305910 466847
rect 306390 454057 314250 466847
rect 314730 454057 314910 466847
rect 315390 454057 323250 466847
rect 323730 454057 323910 466847
rect 324390 454057 332250 466847
rect 306390 419431 332250 454057
rect 306390 401785 314250 419431
rect 314730 401785 314910 419431
rect 315390 401785 323250 419431
rect 323730 401785 323910 419431
rect 324390 401785 332250 419431
rect 332730 401785 332910 466847
rect 333390 401785 341250 466847
rect 341730 401785 341910 466847
rect 342390 401785 350250 466847
rect 305730 364847 350250 401785
rect 305730 299785 305910 364847
rect 306390 351785 314250 364847
rect 314730 351785 314910 364847
rect 315390 351785 323250 364847
rect 306390 330623 323250 351785
rect 306390 299785 314250 330623
rect 314730 299785 314910 330623
rect 315390 299785 323250 330623
rect 323730 299785 323910 364847
rect 324390 299785 332250 364847
rect 332730 299785 332910 364847
rect 333390 299785 341250 364847
rect 341730 299785 341910 364847
rect 342390 299785 350250 364847
rect 305730 262847 350250 299785
rect 305730 197785 305910 262847
rect 306390 249785 314250 262847
rect 314730 249785 314910 262847
rect 315390 249785 323250 262847
rect 306390 228623 323250 249785
rect 306390 197785 314250 228623
rect 314730 197785 314910 228623
rect 315390 197785 323250 228623
rect 323730 197785 323910 262847
rect 324390 197785 332250 262847
rect 332730 197785 332910 262847
rect 333390 197785 341250 262847
rect 341730 197785 341910 262847
rect 342390 197785 350250 262847
rect 305730 160847 350250 197785
rect 305730 2147 305910 160847
rect 306390 149785 314250 160847
rect 314730 149785 314910 160847
rect 315390 149785 323250 160847
rect 306390 128623 323250 149785
rect 306390 93785 314250 128623
rect 314730 93785 314910 128623
rect 315390 93785 323250 128623
rect 323730 93785 323910 160847
rect 324390 93785 332250 160847
rect 306390 56439 332250 93785
rect 306390 2147 314250 56439
rect 314730 2147 314910 56439
rect 315390 2147 323250 56439
rect 323730 2147 323910 56439
rect 324390 45364 332250 56439
rect 332730 45364 332910 160847
rect 324390 5948 332910 45364
rect 324390 2147 332250 5948
rect 332730 2147 332910 5948
rect 333390 2147 341250 160847
rect 341730 2147 341910 160847
rect 342390 2147 350250 160847
rect 350730 2147 350910 587149
rect 351390 508568 359250 587149
rect 351390 462616 354406 508568
rect 354886 462616 355142 508568
rect 355622 462616 359250 508568
rect 351390 406840 359250 462616
rect 351390 360888 354406 406840
rect 354886 360888 355142 406840
rect 355622 360888 359250 406840
rect 351390 354329 359250 360888
rect 359730 457009 359910 587149
rect 360390 457009 368250 587149
rect 368730 457009 368910 587149
rect 369390 457009 377250 587149
rect 377730 457009 377910 587149
rect 378390 457009 386250 587149
rect 386730 457009 386910 587149
rect 387390 457009 395250 587149
rect 359730 418983 395250 457009
rect 359730 354329 359910 418983
rect 360390 354329 368250 418983
rect 368730 354329 368910 418983
rect 369390 354329 377250 418983
rect 377730 354329 377910 418983
rect 378390 354329 386250 418983
rect 386730 354329 386910 418983
rect 387390 354329 395250 418983
rect 351390 315079 395250 354329
rect 351390 304568 359250 315079
rect 351390 258616 354406 304568
rect 354886 258616 355142 304568
rect 355622 258616 359250 304568
rect 351390 252329 359250 258616
rect 359730 252329 359910 315079
rect 360390 252329 368250 315079
rect 368730 252329 368910 315079
rect 369390 252329 377250 315079
rect 377730 252329 377910 315079
rect 378390 252329 386250 315079
rect 386730 252329 386910 315079
rect 387390 252329 395250 315079
rect 351390 213079 395250 252329
rect 351390 202840 359250 213079
rect 351390 156888 354406 202840
rect 354886 156888 355142 202840
rect 355622 156888 359250 202840
rect 351390 150329 359250 156888
rect 359730 150329 359910 213079
rect 360390 150329 368250 213079
rect 368730 150329 368910 213079
rect 369390 150329 377250 213079
rect 377730 150329 377910 213079
rect 378390 150329 386250 213079
rect 386730 150329 386910 213079
rect 387390 150329 395250 213079
rect 351390 111079 395250 150329
rect 351390 98392 359250 111079
rect 351390 53528 354222 98392
rect 354702 53528 359250 98392
rect 351390 2147 359250 53528
rect 359730 2147 359910 111079
rect 360390 95145 368250 111079
rect 368730 95145 368910 111079
rect 369390 95145 377250 111079
rect 377730 95145 377910 111079
rect 378390 95145 386250 111079
rect 386730 95145 386910 111079
rect 387390 95145 395250 111079
rect 395730 95145 395910 587149
rect 396390 95145 404250 587149
rect 360390 56439 404250 95145
rect 360390 2147 368250 56439
rect 368730 2147 368910 56439
rect 369390 2147 377250 56439
rect 377730 2147 377910 56439
rect 378390 2147 386250 56439
rect 386730 2147 386910 56439
rect 387390 2147 395250 56439
rect 395730 2147 395910 56439
rect 396390 2147 404250 56439
rect 404730 2147 404910 587149
rect 405390 503785 413250 587149
rect 413730 503785 413910 587149
rect 414390 503785 422250 587149
rect 422730 503785 422910 587149
rect 423390 503785 431250 587149
rect 431730 503785 431910 587149
rect 432390 503785 440250 587149
rect 440730 503785 440910 587149
rect 441390 503785 449250 587149
rect 449730 561364 449910 587149
rect 450390 561364 458250 587149
rect 449730 521948 458250 561364
rect 449730 503785 449910 521948
rect 450390 503785 458250 521948
rect 405390 501496 458250 503785
rect 405390 466847 455422 501496
rect 405390 454057 413250 466847
rect 413730 454057 413910 466847
rect 414390 454057 422250 466847
rect 422730 454057 422910 466847
rect 423390 454057 431250 466847
rect 405390 419431 431250 454057
rect 405390 401785 413250 419431
rect 413730 401785 413910 419431
rect 414390 401785 422250 419431
rect 422730 401785 422910 419431
rect 423390 401785 431250 419431
rect 431730 401785 431910 466847
rect 432390 401785 440250 466847
rect 440730 401785 440910 466847
rect 441390 401785 449250 466847
rect 449730 401785 449910 466847
rect 450390 462616 455422 466847
rect 455902 462616 456158 501496
rect 456638 462616 458250 501496
rect 450390 458520 458250 462616
rect 450390 456088 454318 458520
rect 454798 456088 458250 458520
rect 450390 401785 458250 456088
rect 405390 399768 458250 401785
rect 405390 364847 455422 399768
rect 405390 299785 413250 364847
rect 413730 299785 413910 364847
rect 414390 351785 422250 364847
rect 422730 351785 422910 364847
rect 423390 351785 431250 364847
rect 414390 330623 431250 351785
rect 414390 299785 422250 330623
rect 422730 299785 422910 330623
rect 423390 299785 431250 330623
rect 431730 299785 431910 364847
rect 432390 299785 440250 364847
rect 440730 299785 440910 364847
rect 441390 299785 449250 364847
rect 449730 299785 449910 364847
rect 450390 360888 455422 364847
rect 455902 360888 456158 399768
rect 456638 360888 458250 399768
rect 450390 356792 458250 360888
rect 450390 353816 453950 356792
rect 454430 353816 454686 356792
rect 455166 353816 458250 356792
rect 450390 299785 458250 353816
rect 405390 297496 458250 299785
rect 405390 262847 455422 297496
rect 405390 197785 413250 262847
rect 413730 197785 413910 262847
rect 414390 250385 422250 262847
rect 422730 250385 422910 262847
rect 423390 250385 431250 262847
rect 414390 229223 431250 250385
rect 414390 197785 422250 229223
rect 422730 197785 422910 229223
rect 423390 197785 431250 229223
rect 431730 197785 431910 262847
rect 432390 197785 440250 262847
rect 440730 197785 440910 262847
rect 441390 197785 449250 262847
rect 449730 197785 449910 262847
rect 450390 258616 455422 262847
rect 455902 258616 456158 297496
rect 456638 258616 458250 297496
rect 450390 255608 458250 258616
rect 450390 252088 453950 255608
rect 454430 252088 454686 255608
rect 455166 252088 458250 255608
rect 450390 197785 458250 252088
rect 405390 195768 458250 197785
rect 405390 160847 455422 195768
rect 405390 93785 413250 160847
rect 413730 93785 413910 160847
rect 414390 147785 422250 160847
rect 422730 147785 422910 160847
rect 423390 147785 431250 160847
rect 414390 126623 431250 147785
rect 414390 93785 422250 126623
rect 422730 93785 422910 126623
rect 423390 93785 431250 126623
rect 431730 93785 431910 160847
rect 432390 93785 440250 160847
rect 405390 56439 440250 93785
rect 405390 2147 413250 56439
rect 413730 2147 413910 56439
rect 414390 2147 422250 56439
rect 422730 2147 422910 56439
rect 423390 2147 431250 56439
rect 431730 2147 431910 56439
rect 432390 2147 440250 56439
rect 440730 2147 440910 160847
rect 441390 2147 449250 160847
rect 449730 45364 449910 160847
rect 450390 156888 455422 160847
rect 455902 156888 456158 195768
rect 456638 156888 458250 195768
rect 450390 152792 458250 156888
rect 450390 149816 453950 152792
rect 454430 149816 454686 152792
rect 455166 149816 458250 152792
rect 450390 45364 458250 149816
rect 449730 5948 458250 45364
rect 449730 2147 449910 5948
rect 450390 2147 458250 5948
rect 458730 2147 458910 587149
rect 459390 80457 467250 587149
rect 467730 80457 467910 587149
rect 468390 492569 476250 587149
rect 476730 492569 476910 587149
rect 477390 492569 485250 587149
rect 485730 492569 485910 587149
rect 486390 492569 494250 587149
rect 468390 461479 494250 492569
rect 468390 441569 476250 461479
rect 476730 441569 476910 461479
rect 477390 441569 485250 461479
rect 485730 441569 485910 461479
rect 486390 441569 494250 461479
rect 468390 409799 494250 441569
rect 468390 390569 476250 409799
rect 476730 390569 476910 409799
rect 477390 390569 485250 409799
rect 485730 390569 485910 409799
rect 486390 390569 494250 409799
rect 468390 359479 494250 390569
rect 468390 333585 476250 359479
rect 476730 333585 476910 359479
rect 477390 333585 485250 359479
rect 485730 333585 485910 359479
rect 486390 333585 494250 359479
rect 494730 498364 494910 587149
rect 495390 498364 503250 587149
rect 494730 458948 503250 498364
rect 494730 396364 494910 458948
rect 495390 396364 503250 458948
rect 494730 356948 503250 396364
rect 494730 333585 494910 356948
rect 495390 333585 503250 356948
rect 468390 306031 503250 333585
rect 468390 288569 476250 306031
rect 476730 288569 476910 306031
rect 477390 288569 485250 306031
rect 485730 288569 485910 306031
rect 486390 288569 494250 306031
rect 468390 257479 494250 288569
rect 468390 231585 476250 257479
rect 476730 231585 476910 257479
rect 477390 231585 485250 257479
rect 485730 231585 485910 257479
rect 486390 231585 494250 257479
rect 494730 294364 494910 306031
rect 495390 294364 503250 306031
rect 494730 254948 503250 294364
rect 494730 231585 494910 254948
rect 495390 231585 503250 254948
rect 468390 204031 503250 231585
rect 468390 186569 476250 204031
rect 476730 186569 476910 204031
rect 477390 186569 485250 204031
rect 485730 186569 485910 204031
rect 486390 186569 494250 204031
rect 468390 155479 494250 186569
rect 468390 129585 476250 155479
rect 476730 129585 476910 155479
rect 477390 129585 485250 155479
rect 485730 129585 485910 155479
rect 486390 129585 494250 155479
rect 494730 192364 494910 204031
rect 495390 192364 503250 204031
rect 494730 152948 503250 192364
rect 494730 129585 494910 152948
rect 495390 129585 503250 152948
rect 468390 102031 503250 129585
rect 468390 80457 476250 102031
rect 476730 80457 476910 102031
rect 477390 80457 485250 102031
rect 459390 56167 485250 80457
rect 459390 2147 467250 56167
rect 467730 2147 467910 56167
rect 468390 2147 476250 56167
rect 476730 2147 476910 56167
rect 477390 2147 485250 56167
rect 485730 2147 485910 102031
rect 486390 2147 494250 102031
rect 494730 2147 494910 102031
rect 495390 2147 503250 102031
rect 503730 2147 503910 587149
rect 504390 2147 512250 587149
rect 512730 2147 512910 587149
rect 513390 2147 521250 587149
rect 521730 2147 521910 587149
rect 522390 2147 530250 587149
rect 530730 2147 530910 587149
rect 531390 2147 539250 587149
rect 539730 2147 539910 587149
rect 540390 2147 548250 587149
rect 548730 501364 548910 587149
rect 548730 461948 549234 501364
rect 548730 399364 548910 461948
rect 548730 359948 549234 399364
rect 548730 297364 548910 359948
rect 548730 257948 549234 297364
rect 548730 195364 548910 257948
rect 548730 155948 549234 195364
rect 548730 2147 548910 155948
<< metal5 >>
rect 1042 581876 560866 582196
rect 1042 581216 560866 581536
rect 1042 570876 560866 571196
rect 1042 570216 560866 570536
rect 1042 559876 560866 560196
rect 1042 559216 560866 559536
rect 1042 548876 560866 549196
rect 1042 548216 560866 548536
rect 1042 537876 560866 538196
rect 1042 537216 560866 537536
rect 1042 526876 560866 527196
rect 1042 526216 560866 526536
rect 1042 515876 560866 516196
rect 1042 515216 560866 515536
rect 1042 504876 560866 505196
rect 1042 504216 560866 504536
rect 1042 493876 560866 494196
rect 1042 493216 560866 493536
rect 1042 482876 560866 483196
rect 1042 482216 560866 482536
rect 1042 471876 560866 472196
rect 1042 471216 560866 471536
rect 1042 460876 560866 461196
rect 1042 460216 560866 460536
rect 1042 449876 560866 450196
rect 1042 449216 560866 449536
rect 1042 438876 560866 439196
rect 1042 438216 560866 438536
rect 1042 427876 560866 428196
rect 1042 427216 560866 427536
rect 1042 416876 560866 417196
rect 1042 416216 560866 416536
rect 1042 405876 560866 406196
rect 1042 405216 560866 405536
rect 1042 394876 560866 395196
rect 1042 394216 560866 394536
rect 1042 383876 560866 384196
rect 1042 383216 560866 383536
rect 1042 372876 560866 373196
rect 1042 372216 560866 372536
rect 1042 361876 560866 362196
rect 1042 361216 560866 361536
rect 1042 350876 560866 351196
rect 1042 350216 560866 350536
rect 1042 339876 560866 340196
rect 1042 339216 560866 339536
rect 1042 328876 560866 329196
rect 1042 328216 560866 328536
rect 1042 317876 560866 318196
rect 1042 317216 560866 317536
rect 1042 306876 560866 307196
rect 1042 306216 560866 306536
rect 1042 295876 560866 296196
rect 1042 295216 560866 295536
rect 1042 284876 560866 285196
rect 1042 284216 560866 284536
rect 1042 273876 560866 274196
rect 1042 273216 560866 273536
rect 1042 262876 560866 263196
rect 1042 262216 560866 262536
rect 1042 251876 560866 252196
rect 1042 251216 560866 251536
rect 1042 240876 560866 241196
rect 1042 240216 560866 240536
rect 1042 229876 560866 230196
rect 1042 229216 560866 229536
rect 1042 218876 560866 219196
rect 1042 218216 560866 218536
rect 1042 207876 560866 208196
rect 1042 207216 560866 207536
rect 1042 196876 560866 197196
rect 1042 196216 560866 196536
rect 1042 185876 560866 186196
rect 1042 185216 560866 185536
rect 1042 174876 560866 175196
rect 1042 174216 560866 174536
rect 1042 163876 560866 164196
rect 1042 163216 560866 163536
rect 1042 152876 560866 153196
rect 1042 152216 560866 152536
rect 1042 141876 560866 142196
rect 1042 141216 560866 141536
rect 1042 130876 560866 131196
rect 1042 130216 560866 130536
rect 1042 119876 560866 120196
rect 1042 119216 560866 119536
rect 1042 108876 560866 109196
rect 1042 108216 560866 108536
rect 1042 97876 560866 98196
rect 1042 97216 560866 97536
rect 1042 86876 560866 87196
rect 1042 86216 560866 86536
rect 1042 75876 560866 76196
rect 1042 75216 560866 75536
rect 1042 64876 560866 65196
rect 1042 64216 560866 64536
rect 1042 53876 560866 54196
rect 1042 53216 560866 53536
rect 1042 42876 560866 43196
rect 1042 42216 560866 42536
rect 1042 31876 560866 32196
rect 1042 31216 560866 31536
rect 1042 20876 560866 21196
rect 1042 20216 560866 20536
rect 1042 9876 560866 10196
rect 1042 9216 560866 9536
<< labels >>
rlabel metal3 s 186 327568 786 327688 6 ccff_head
port 1 nsew signal input
rlabel metal2 s 79216 589000 79272 589600 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 561186 408488 561786 408608 6 clk
port 3 nsew signal input
rlabel metal2 s 81792 0 81848 600 6 gfpga_pad_GPIO_PAD_in[0]
port 4 nsew signal input
rlabel metal2 s 474632 0 474688 600 6 gfpga_pad_GPIO_PAD_in[10]
port 5 nsew signal input
rlabel metal2 s 390268 589000 390324 589600 6 gfpga_pad_GPIO_PAD_in[11]
port 6 nsew signal input
rlabel metal2 s 324580 589000 324636 589600 6 gfpga_pad_GPIO_PAD_in[12]
port 7 nsew signal input
rlabel metal2 s 291736 589000 291792 589600 6 gfpga_pad_GPIO_PAD_in[13]
port 8 nsew signal input
rlabel metal2 s 425044 0 425100 600 6 gfpga_pad_GPIO_PAD_in[14]
port 9 nsew signal input
rlabel metal2 s 455312 589000 455368 589600 6 gfpga_pad_GPIO_PAD_in[15]
port 10 nsew signal input
rlabel metal3 s 186 120168 786 120288 6 gfpga_pad_GPIO_PAD_in[16]
port 11 nsew signal input
rlabel metal3 s 186 466288 786 466408 6 gfpga_pad_GPIO_PAD_in[17]
port 12 nsew signal input
rlabel metal2 s 163580 0 163636 600 6 gfpga_pad_GPIO_PAD_in[18]
port 13 nsew signal input
rlabel metal2 s 537100 589000 537156 589600 6 gfpga_pad_GPIO_PAD_in[19]
port 14 nsew signal input
rlabel metal3 s 186 172528 786 172648 6 gfpga_pad_GPIO_PAD_in[1]
port 15 nsew signal input
rlabel metal2 s 343256 0 343312 600 6 gfpga_pad_GPIO_PAD_in[20]
port 16 nsew signal input
rlabel metal2 s 46372 589000 46428 589600 6 gfpga_pad_GPIO_PAD_in[21]
port 17 nsew signal input
rlabel metal2 s 488156 589000 488212 589600 6 gfpga_pad_GPIO_PAD_in[22]
port 18 nsew signal input
rlabel metal3 s 186 241208 786 241328 6 gfpga_pad_GPIO_PAD_in[23]
port 19 nsew signal input
rlabel metal3 s 561186 252768 561786 252888 6 gfpga_pad_GPIO_PAD_in[24]
port 20 nsew signal input
rlabel metal2 s 521000 589000 521056 589600 6 gfpga_pad_GPIO_PAD_in[25]
port 21 nsew signal input
rlabel metal2 s 179680 0 179736 600 6 gfpga_pad_GPIO_PAD_in[26]
port 22 nsew signal input
rlabel metal3 s 186 293568 786 293688 6 gfpga_pad_GPIO_PAD_in[27]
port 23 nsew signal input
rlabel metal3 s 186 431608 786 431728 6 gfpga_pad_GPIO_PAD_in[28]
port 24 nsew signal input
rlabel metal2 s 62472 589000 62528 589600 6 gfpga_pad_GPIO_PAD_in[29]
port 25 nsew signal input
rlabel metal3 s 561186 442488 561786 442608 6 gfpga_pad_GPIO_PAD_in[2]
port 26 nsew signal input
rlabel metal3 s 186 68488 786 68608 6 gfpga_pad_GPIO_PAD_in[30]
port 27 nsew signal input
rlabel metal2 s 193848 589000 193904 589600 6 gfpga_pad_GPIO_PAD_in[31]
port 28 nsew signal input
rlabel metal3 s 186 310568 786 310688 6 gfpga_pad_GPIO_PAD_in[32]
port 29 nsew signal input
rlabel metal3 s 561186 27688 561786 27808 6 gfpga_pad_GPIO_PAD_in[33]
port 30 nsew signal input
rlabel metal3 s 561186 183408 561786 183528 6 gfpga_pad_GPIO_PAD_in[34]
port 31 nsew signal input
rlabel metal3 s 561186 235088 561786 235208 6 gfpga_pad_GPIO_PAD_in[35]
port 32 nsew signal input
rlabel metal3 s 561186 269768 561786 269888 6 gfpga_pad_GPIO_PAD_in[36]
port 33 nsew signal input
rlabel metal2 s 245368 0 245424 600 6 gfpga_pad_GPIO_PAD_in[37]
port 34 nsew signal input
rlabel metal2 s 275636 589000 275692 589600 6 gfpga_pad_GPIO_PAD_in[38]
port 35 nsew signal input
rlabel metal2 s 490732 0 490788 600 6 gfpga_pad_GPIO_PAD_in[39]
port 36 nsew signal input
rlabel metal3 s 561186 10688 561786 10808 6 gfpga_pad_GPIO_PAD_in[3]
port 37 nsew signal input
rlabel metal3 s 561186 304448 561786 304568 6 gfpga_pad_GPIO_PAD_in[40]
port 38 nsew signal input
rlabel metal2 s 258892 589000 258948 589600 6 gfpga_pad_GPIO_PAD_in[41]
port 39 nsew signal input
rlabel metal2 s 242792 589000 242848 589600 6 gfpga_pad_GPIO_PAD_in[42]
port 40 nsew signal input
rlabel metal3 s 186 413928 786 414048 6 gfpga_pad_GPIO_PAD_in[43]
port 41 nsew signal input
rlabel metal2 s 357424 589000 357480 589600 6 gfpga_pad_GPIO_PAD_in[44]
port 42 nsew signal input
rlabel metal2 s 360000 0 360056 600 6 gfpga_pad_GPIO_PAD_in[45]
port 43 nsew signal input
rlabel metal2 s 294312 0 294368 600 6 gfpga_pad_GPIO_PAD_in[46]
port 44 nsew signal input
rlabel metal2 s 112060 589000 112116 589600 6 gfpga_pad_GPIO_PAD_in[47]
port 45 nsew signal input
rlabel metal3 s 561186 356128 561786 356248 6 gfpga_pad_GPIO_PAD_in[48]
port 46 nsew signal input
rlabel metal3 s 186 569648 786 569768 6 gfpga_pad_GPIO_PAD_in[49]
port 47 nsew signal input
rlabel metal2 s 130736 0 130792 600 6 gfpga_pad_GPIO_PAD_in[4]
port 48 nsew signal input
rlabel metal2 s 472056 589000 472112 589600 6 gfpga_pad_GPIO_PAD_in[50]
port 49 nsew signal input
rlabel metal3 s 561186 511848 561786 511968 6 gfpga_pad_GPIO_PAD_in[51]
port 50 nsew signal input
rlabel metal3 s 186 345248 786 345368 6 gfpga_pad_GPIO_PAD_in[52]
port 51 nsew signal input
rlabel metal2 s 146836 0 146892 600 6 gfpga_pad_GPIO_PAD_in[53]
port 52 nsew signal input
rlabel metal3 s 186 587328 786 587448 6 gfpga_pad_GPIO_PAD_in[54]
port 53 nsew signal input
rlabel metal3 s 561186 166408 561786 166528 6 gfpga_pad_GPIO_PAD_in[55]
port 54 nsew signal input
rlabel metal2 s 177104 589000 177160 589600 6 gfpga_pad_GPIO_PAD_in[56]
port 55 nsew signal input
rlabel metal2 s 556420 0 556476 600 6 gfpga_pad_GPIO_PAD_in[57]
port 56 nsew signal input
rlabel metal3 s 561186 477168 561786 477288 6 gfpga_pad_GPIO_PAD_in[58]
port 57 nsew signal input
rlabel metal3 s 561186 80048 561786 80168 6 gfpga_pad_GPIO_PAD_in[59]
port 58 nsew signal input
rlabel metal2 s 553844 589000 553900 589600 6 gfpga_pad_GPIO_PAD_in[5]
port 59 nsew signal input
rlabel metal3 s 561186 460168 561786 460288 6 gfpga_pad_GPIO_PAD_in[60]
port 60 nsew signal input
rlabel metal3 s 561186 114728 561786 114848 6 gfpga_pad_GPIO_PAD_in[61]
port 61 nsew signal input
rlabel metal2 s 228624 0 228680 600 6 gfpga_pad_GPIO_PAD_in[62]
port 62 nsew signal input
rlabel metal3 s 186 379928 786 380048 6 gfpga_pad_GPIO_PAD_in[63]
port 63 nsew signal input
rlabel metal2 s 16104 0 16160 600 6 gfpga_pad_GPIO_PAD_in[6]
port 64 nsew signal input
rlabel metal3 s 186 258888 786 259008 6 gfpga_pad_GPIO_PAD_in[7]
port 65 nsew signal input
rlabel metal2 s 408944 0 409000 600 6 gfpga_pad_GPIO_PAD_in[8]
port 66 nsew signal input
rlabel metal3 s 186 103168 786 103288 6 gfpga_pad_GPIO_PAD_in[9]
port 67 nsew signal input
rlabel metal2 s 128160 589000 128216 589600 6 gfpga_pad_GPIO_PAD_out[0]
port 68 nsew signal output
rlabel metal3 s 561186 546528 561786 546648 6 gfpga_pad_GPIO_PAD_out[10]
port 69 nsew signal output
rlabel metal3 s 186 396928 786 397048 6 gfpga_pad_GPIO_PAD_out[11]
port 70 nsew signal output
rlabel metal3 s 186 137848 786 137968 6 gfpga_pad_GPIO_PAD_out[12]
port 71 nsew signal output
rlabel metal2 s 29628 589000 29684 589600 6 gfpga_pad_GPIO_PAD_out[13]
port 72 nsew signal output
rlabel metal2 s 161004 589000 161060 589600 6 gfpga_pad_GPIO_PAD_out[14]
port 73 nsew signal output
rlabel metal2 s 209948 589000 210004 589600 6 gfpga_pad_GPIO_PAD_out[15]
port 74 nsew signal output
rlabel metal3 s 186 206528 786 206648 6 gfpga_pad_GPIO_PAD_out[16]
port 75 nsew signal output
rlabel metal3 s 186 86168 786 86288 6 gfpga_pad_GPIO_PAD_out[17]
port 76 nsew signal output
rlabel metal3 s 561186 201088 561786 201208 6 gfpga_pad_GPIO_PAD_out[18]
port 77 nsew signal output
rlabel metal3 s 561186 563528 561786 563648 6 gfpga_pad_GPIO_PAD_out[19]
port 78 nsew signal output
rlabel metal2 s 48948 0 49004 600 6 gfpga_pad_GPIO_PAD_out[1]
port 79 nsew signal output
rlabel metal3 s 561186 45368 561786 45488 6 gfpga_pad_GPIO_PAD_out[20]
port 80 nsew signal output
rlabel metal3 s 561186 218088 561786 218208 6 gfpga_pad_GPIO_PAD_out[21]
port 81 nsew signal output
rlabel metal2 s 373524 589000 373580 589600 6 gfpga_pad_GPIO_PAD_out[22]
port 82 nsew signal output
rlabel metal3 s 561186 131728 561786 131848 6 gfpga_pad_GPIO_PAD_out[23]
port 83 nsew signal output
rlabel metal2 s 523576 0 523632 600 6 gfpga_pad_GPIO_PAD_out[24]
port 84 nsew signal output
rlabel metal2 s 261468 0 261524 600 6 gfpga_pad_GPIO_PAD_out[25]
port 85 nsew signal output
rlabel metal3 s 561186 322128 561786 322248 6 gfpga_pad_GPIO_PAD_out[26]
port 86 nsew signal output
rlabel metal3 s 561186 581208 561786 581328 6 gfpga_pad_GPIO_PAD_out[27]
port 87 nsew signal output
rlabel metal3 s 186 224208 786 224328 6 gfpga_pad_GPIO_PAD_out[28]
port 88 nsew signal output
rlabel metal3 s 186 275888 786 276008 6 gfpga_pad_GPIO_PAD_out[29]
port 89 nsew signal output
rlabel metal3 s 186 51488 786 51608 6 gfpga_pad_GPIO_PAD_out[2]
port 90 nsew signal output
rlabel metal2 s 539676 0 539732 600 6 gfpga_pad_GPIO_PAD_out[30]
port 91 nsew signal output
rlabel metal2 s 226048 589000 226104 589600 6 gfpga_pad_GPIO_PAD_out[31]
port 92 nsew signal output
rlabel metal2 s 441788 0 441844 600 6 gfpga_pad_GPIO_PAD_out[32]
port 93 nsew signal output
rlabel metal2 s 65048 0 65104 600 6 gfpga_pad_GPIO_PAD_out[33]
port 94 nsew signal output
rlabel metal2 s 212524 0 212580 600 6 gfpga_pad_GPIO_PAD_out[34]
port 95 nsew signal output
rlabel metal3 s 561186 62368 561786 62488 6 gfpga_pad_GPIO_PAD_out[35]
port 96 nsew signal output
rlabel metal3 s 561186 425488 561786 425608 6 gfpga_pad_GPIO_PAD_out[36]
port 97 nsew signal output
rlabel metal3 s 186 16808 786 16928 6 gfpga_pad_GPIO_PAD_out[37]
port 98 nsew signal output
rlabel metal2 s 457888 0 457944 600 6 gfpga_pad_GPIO_PAD_out[38]
port 99 nsew signal output
rlabel metal3 s 186 362248 786 362368 6 gfpga_pad_GPIO_PAD_out[39]
port 100 nsew signal output
rlabel metal3 s 561186 148728 561786 148848 6 gfpga_pad_GPIO_PAD_out[3]
port 101 nsew signal output
rlabel metal3 s 186 483288 786 483408 6 gfpga_pad_GPIO_PAD_out[40]
port 102 nsew signal output
rlabel metal3 s 561186 339128 561786 339248 6 gfpga_pad_GPIO_PAD_out[41]
port 103 nsew signal output
rlabel metal3 s 561186 494848 561786 494968 6 gfpga_pad_GPIO_PAD_out[42]
port 104 nsew signal output
rlabel metal2 s 506832 0 506888 600 6 gfpga_pad_GPIO_PAD_out[43]
port 105 nsew signal output
rlabel metal3 s 561186 529528 561786 529648 6 gfpga_pad_GPIO_PAD_out[44]
port 106 nsew signal output
rlabel metal3 s 186 33808 786 33928 6 gfpga_pad_GPIO_PAD_out[45]
port 107 nsew signal output
rlabel metal3 s 186 517968 786 518088 6 gfpga_pad_GPIO_PAD_out[46]
port 108 nsew signal output
rlabel metal3 s 186 189528 786 189648 6 gfpga_pad_GPIO_PAD_out[47]
port 109 nsew signal output
rlabel metal2 s 4 0 60 600 6 gfpga_pad_GPIO_PAD_out[48]
port 110 nsew signal output
rlabel metal2 s 376100 0 376156 600 6 gfpga_pad_GPIO_PAD_out[49]
port 111 nsew signal output
rlabel metal3 s 186 552648 786 552768 6 gfpga_pad_GPIO_PAD_out[4]
port 112 nsew signal output
rlabel metal2 s 144260 589000 144316 589600 6 gfpga_pad_GPIO_PAD_out[50]
port 113 nsew signal output
rlabel metal2 s 340680 589000 340736 589600 6 gfpga_pad_GPIO_PAD_out[51]
port 114 nsew signal output
rlabel metal3 s 186 448608 786 448728 6 gfpga_pad_GPIO_PAD_out[52]
port 115 nsew signal output
rlabel metal2 s 97892 0 97948 600 6 gfpga_pad_GPIO_PAD_out[53]
port 116 nsew signal output
rlabel metal2 s 32204 0 32260 600 6 gfpga_pad_GPIO_PAD_out[54]
port 117 nsew signal output
rlabel metal2 s 439212 589000 439268 589600 6 gfpga_pad_GPIO_PAD_out[55]
port 118 nsew signal output
rlabel metal2 s 308480 589000 308536 589600 6 gfpga_pad_GPIO_PAD_out[56]
port 119 nsew signal output
rlabel metal2 s 278212 0 278268 600 6 gfpga_pad_GPIO_PAD_out[57]
port 120 nsew signal output
rlabel metal2 s 504900 589000 504956 589600 6 gfpga_pad_GPIO_PAD_out[58]
port 121 nsew signal output
rlabel metal3 s 561186 97048 561786 97168 6 gfpga_pad_GPIO_PAD_out[59]
port 122 nsew signal output
rlabel metal3 s 186 534968 786 535088 6 gfpga_pad_GPIO_PAD_out[5]
port 123 nsew signal output
rlabel metal3 s 561186 373808 561786 373928 6 gfpga_pad_GPIO_PAD_out[60]
port 124 nsew signal output
rlabel metal2 s 113992 0 114048 600 6 gfpga_pad_GPIO_PAD_out[61]
port 125 nsew signal output
rlabel metal2 s 195780 0 195836 600 6 gfpga_pad_GPIO_PAD_out[62]
port 126 nsew signal output
rlabel metal2 s 310412 0 310468 600 6 gfpga_pad_GPIO_PAD_out[63]
port 127 nsew signal output
rlabel metal3 s 561186 390808 561786 390928 6 gfpga_pad_GPIO_PAD_out[6]
port 128 nsew signal output
rlabel metal2 s 327156 0 327212 600 6 gfpga_pad_GPIO_PAD_out[7]
port 129 nsew signal output
rlabel metal2 s 422468 589000 422524 589600 6 gfpga_pad_GPIO_PAD_out[8]
port 130 nsew signal output
rlabel metal2 s 406368 589000 406424 589600 6 gfpga_pad_GPIO_PAD_out[9]
port 131 nsew signal output
rlabel metal2 s 13528 589000 13584 589600 6 pReset
port 132 nsew signal input
rlabel metal2 s 95316 589000 95372 589600 6 prog_clk
port 133 nsew signal input
rlabel metal2 s 392200 0 392256 600 6 reset
port 134 nsew signal input
rlabel metal3 s 186 154848 786 154968 6 set
port 135 nsew signal input
rlabel metal3 s 186 500968 786 501088 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 8330 1928 8650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 17330 1928 17650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 26330 1928 26650 107868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 26330 147444 26650 209868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 26330 249444 26650 311868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 26330 351444 26650 413868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 26330 453444 26650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 35330 1928 35650 30868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 35330 70444 35650 160359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 35330 199089 35650 262359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 35330 301089 35650 364359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 35330 403089 35650 466359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 35330 505089 35650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 44330 1928 44650 34079 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 44330 69953 44650 160359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 44330 199089 44650 262359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 44330 301089 44650 364359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 44330 403089 44650 466359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 44330 505089 44650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 53330 1928 53650 160359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 53330 199089 53650 262359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 53330 301089 53650 364359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 53330 403089 53650 466359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 53330 505089 53650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 62330 1928 62650 109868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 62330 149444 62650 211868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 62330 251444 62650 313868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 62330 353444 62650 415868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 62330 455444 62650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 71330 1928 71650 117567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 71330 148681 71650 219567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 71330 250681 71650 321567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 71330 352681 71650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 80330 1928 80650 117567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 80330 148681 80650 219567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 80330 250681 80650 321567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 80330 352681 80650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 89330 1928 89650 117567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 89330 148681 89650 219567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 89330 250681 89650 321567 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 89330 352681 89650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 98330 1928 98650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 1928 107650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 93865 107650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 197865 107650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 299865 107650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 401865 107650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 454137 107650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 107330 503865 107650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 1928 116650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 93865 116650 126543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 147865 116650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 197865 116650 228543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 249865 116650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 299865 116650 330543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 351865 116650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 401865 116650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 454137 116650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 116330 503865 116650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 125330 1928 125650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 125330 93865 125650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 125330 197865 125650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 125330 299865 125650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 125330 401865 125650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 125330 503865 125650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 134330 1928 134650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 134330 197865 134650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 134330 299865 134650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 134330 401865 134650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 134330 503865 134650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 143330 1928 143650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 143330 197865 143650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 143330 299865 143650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 143330 401865 143650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 143330 503865 143650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 152330 1928 152650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 161330 1928 161650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 161330 150409 161650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 161330 252409 161650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 161330 354409 161650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 161330 457089 161650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 170330 1928 170650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 170330 95225 170650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 170330 150409 170650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 170330 252409 170650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 170330 354409 170650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 170330 457089 170650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 179330 1928 179650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 179330 95225 179650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 179330 150409 179650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 179330 252409 179650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 179330 354409 179650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 179330 457089 179650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 188330 1928 188650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 188330 95225 188650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 197330 1928 197650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 206330 1928 206650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 206330 197865 206650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 206330 299865 206650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 206330 401865 206650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 206330 503865 206650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 1928 215650 5868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 45444 215650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 93865 215650 126543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 147865 215650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 197865 215650 228543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 249865 215650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 299865 215650 330543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 351865 215650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 401865 215650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 454137 215650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 503865 215650 521868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 215330 561444 215650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 1928 224650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 93865 224650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 197865 224650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 299865 224650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 401865 224650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 454137 224650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 224330 503865 224650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 233330 1928 233650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 233330 197865 233650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 233330 299865 233650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 233330 401865 233650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 233330 503865 233650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 242330 1928 242650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 242330 197865 242650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 242330 299865 242650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 242330 401865 242650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 242330 503865 242650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 251330 1928 251650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 260330 1928 260650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 260330 150409 260650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 260330 252409 260650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 260330 354409 260650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 260330 457089 260650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 269330 1928 269650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 269330 95225 269650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 269330 150409 269650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 269330 252409 269650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 269330 354409 269650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 269330 457089 269650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 278330 1928 278650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 278330 95225 278650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 278330 150409 278650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 278330 252409 278650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 278330 354409 278650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 278330 457089 278650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 287330 1928 287650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 287330 95225 287650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 287330 150409 287650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 287330 252409 287650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 287330 354409 287650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 296330 1928 296650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 296330 95225 296650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 305330 1928 305650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 1928 314650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 93865 314650 128543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 149865 314650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 197865 314650 228543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 249865 314650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 299865 314650 330543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 351865 314650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 401865 314650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 454137 314650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 314330 503865 314650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 1928 323650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 93865 323650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 197865 323650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 299865 323650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 401865 323650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 454137 323650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 323330 503865 323650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 1928 332650 5868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 45444 332650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 197865 332650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 299865 332650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 401865 332650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 503865 332650 521868 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 332330 561444 332650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 341330 1928 341650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 341330 197865 341650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 341330 299865 341650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 341330 401865 341650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 341330 503865 341650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 350330 1928 350650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 359330 1928 359650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 359330 150409 359650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 359330 252409 359650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 359330 354409 359650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 368330 1928 368650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 368330 95225 368650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 368330 150409 368650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 368330 252409 368650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 368330 354409 368650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 368330 457089 368650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 377330 1928 377650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 377330 95225 377650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 377330 150409 377650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 377330 252409 377650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 377330 354409 377650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 377330 457089 377650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 386330 1928 386650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 386330 95225 386650 110999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 386330 150409 386650 212999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 386330 252409 386650 314999 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 386330 354409 386650 418903 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 386330 457089 386650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 395330 1928 395650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 395330 95225 395650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 404330 1928 404650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 1928 413650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 93865 413650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 197865 413650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 299865 413650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 401865 413650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 454137 413650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 413330 503865 413650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 1928 422650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 93865 422650 126543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 147865 422650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 197865 422650 229143 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 250465 422650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 299865 422650 330543 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 351865 422650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 401865 422650 419351 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 454137 422650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 422330 503865 422650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 431330 1928 431650 56359 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 431330 93865 431650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 431330 197865 431650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 431330 299865 431650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 431330 401865 431650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 431330 503865 431650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 440330 1928 440650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 440330 197865 440650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 440330 299865 440650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 440330 401865 440650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 440330 503865 440650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 449330 1928 449650 160767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 449330 197865 449650 262767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 449330 299865 449650 364767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 449330 401865 449650 466767 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 449330 503865 449650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 458330 1928 458650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 467330 1928 467650 56087 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 467330 80537 467650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 1928 476650 56087 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 80537 476650 101951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 129665 476650 155399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 186649 476650 203951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 231665 476650 257399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 288649 476650 305951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 333665 476650 359399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 390649 476650 409719 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 441649 476650 461399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 476330 492649 476650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 1928 485650 101951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 129665 485650 155399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 186649 485650 203951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 231665 485650 257399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 288649 485650 305951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 333665 485650 359399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 390649 485650 409719 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 441649 485650 461399 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 485330 492649 485650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 494330 1928 494650 101951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 494330 129665 494650 203951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 494330 231665 494650 305951 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 494330 333665 494650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 503330 1928 503650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 512330 1928 512650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 521330 1928 521650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 530330 1928 530650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 539330 1928 539650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 548330 1928 548650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 557330 1928 557650 587368 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 9216 560866 9536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 20216 560866 20536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 31216 560866 31536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 42216 560866 42536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 53216 560866 53536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 64216 560866 64536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 75216 560866 75536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 86216 560866 86536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 97216 560866 97536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 108216 560866 108536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 119216 560866 119536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 130216 560866 130536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 141216 560866 141536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 152216 560866 152536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 163216 560866 163536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 174216 560866 174536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 185216 560866 185536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 196216 560866 196536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 207216 560866 207536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 218216 560866 218536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 229216 560866 229536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 240216 560866 240536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 251216 560866 251536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 262216 560866 262536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 273216 560866 273536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 284216 560866 284536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 295216 560866 295536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 306216 560866 306536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 317216 560866 317536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 328216 560866 328536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 339216 560866 339536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 350216 560866 350536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 361216 560866 361536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 372216 560866 372536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 383216 560866 383536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 394216 560866 394536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 405216 560866 405536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 416216 560866 416536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 427216 560866 427536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 438216 560866 438536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 449216 560866 449536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 460216 560866 460536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 471216 560866 471536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 482216 560866 482536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 493216 560866 493536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 504216 560866 504536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 515216 560866 515536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 526216 560866 526536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 537216 560866 537536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 548216 560866 548536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 559216 560866 559536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 570216 560866 570536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal5 s 1042 581216 560866 581536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 2494 104744 2814 150536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 102406 209192 102726 254440 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 201398 53608 201718 98312 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 301494 156968 301814 202760 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 354486 258696 354806 304488 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 454030 353896 454350 356712 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 2494 207016 2814 252808 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 100934 106920 101254 152712 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 199742 156968 200062 202760 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 301494 258696 301814 304488 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 354302 53608 354622 98312 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 454398 456168 454718 458440 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 2494 308744 2814 354536 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 100934 413192 101254 458440 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 201398 109096 201718 152712 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 301494 360968 301814 406760 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 354486 156968 354806 202760 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 454030 252168 454350 255528 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 2494 411016 2814 456808 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 100934 310920 101254 356712 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 201398 211368 201718 253896 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 301494 462696 301814 508488 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 354486 360968 354806 406760 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 454030 149896 454350 152712 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 199742 259240 200062 303944 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 354486 462696 354806 508488 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 455502 156968 455822 195688 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 201398 313640 201718 356168 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 455502 258696 455822 297416 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 199742 361512 200062 406216 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 455502 462696 455822 501416 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 201398 414824 201718 458440 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 455502 360968 455822 399688 6 vccd1
port 136 nsew signal bidirectional
rlabel metal4 s 199742 462696 200062 508488 6 vccd1
port 136 nsew signal bidirectional
rlabel metal3 s 561186 287448 561786 287568 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 8990 1928 9310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 17990 1928 18310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 26990 1928 27310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 35990 1928 36310 34079 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 35990 69953 36310 160359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 35990 199089 36310 262359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 35990 301089 36310 364359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 35990 403089 36310 466359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 35990 505089 36310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 44990 1928 45310 34079 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 44990 69953 45310 160359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 44990 199089 45310 262359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 44990 301089 45310 364359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 44990 403089 45310 466359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 44990 505089 45310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 53990 1928 54310 160359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 53990 199089 54310 262359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 53990 301089 54310 364359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 53990 403089 54310 466359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 53990 505089 54310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 62990 1928 63310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 71990 1928 72310 117567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 71990 148681 72310 219567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 71990 250681 72310 321567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 71990 352681 72310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 80990 1928 81310 117567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 80990 148681 81310 219567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 80990 250681 81310 321567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 80990 352681 81310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 89990 1928 90310 117567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 89990 148681 90310 219567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 89990 250681 90310 321567 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 89990 352681 90310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 98990 1928 99310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 1928 108310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 93865 108310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 197865 108310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 299865 108310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 401865 108310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 454137 108310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 107990 503865 108310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 1928 117310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 93865 117310 126543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 147865 117310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 197865 117310 228543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 249865 117310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 299865 117310 330543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 351865 117310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 401865 117310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 454137 117310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 116990 503865 117310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 125990 1928 126310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 125990 93865 126310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 125990 197865 126310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 125990 299865 126310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 125990 401865 126310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 125990 503865 126310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 134990 1928 135310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 134990 197865 135310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 134990 299865 135310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 134990 401865 135310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 134990 503865 135310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 1928 144310 5868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 45444 144310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 197865 144310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 299865 144310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 401865 144310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 503865 144310 521868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 143990 561444 144310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 152990 1928 153310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 161990 1928 162310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 161990 150409 162310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 161990 252409 162310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 161990 354409 162310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 161990 457089 162310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 170990 1928 171310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 170990 95225 171310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 170990 150409 171310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 170990 252409 171310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 170990 354409 171310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 170990 457089 171310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 179990 1928 180310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 179990 95225 180310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 179990 150409 180310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 179990 252409 180310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 179990 354409 180310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 179990 457089 180310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 188990 1928 189310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 188990 95225 189310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 197990 1928 198310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 206990 1928 207310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 206990 197865 207310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 206990 299865 207310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 206990 401865 207310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 206990 454137 207310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 206990 503865 207310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 1928 216310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 93865 216310 126543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 147865 216310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 197865 216310 228543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 249865 216310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 299865 216310 330543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 351865 216310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 401865 216310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 454137 216310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 215990 503865 216310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 224990 1928 225310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 224990 93865 225310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 224990 197865 225310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 224990 299865 225310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 224990 401865 225310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 224990 503865 225310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 233990 1928 234310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 233990 197865 234310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 233990 299865 234310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 233990 401865 234310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 233990 503865 234310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 242990 1928 243310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 242990 197865 243310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 242990 299865 243310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 242990 401865 243310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 242990 503865 243310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 251990 1928 252310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 260990 1928 261310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 260990 150409 261310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 260990 252409 261310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 260990 354409 261310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 260990 457089 261310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 269990 1928 270310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 269990 95225 270310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 269990 150409 270310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 269990 252409 270310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 269990 354409 270310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 269990 457089 270310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 278990 1928 279310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 278990 95225 279310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 278990 150409 279310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 278990 252409 279310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 278990 354409 279310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 278990 457089 279310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 287990 1928 288310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 287990 95225 288310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 296990 1928 297310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 296990 95225 297310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 305990 1928 306310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 305990 197865 306310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 305990 299865 306310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 305990 401865 306310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 305990 503865 306310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 1928 315310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 93865 315310 128543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 149865 315310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 197865 315310 228543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 249865 315310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 299865 315310 330543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 351865 315310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 401865 315310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 454137 315310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 314990 503865 315310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 1928 324310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 93865 324310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 197865 324310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 299865 324310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 401865 324310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 454137 324310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 323990 503865 324310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 332990 1928 333310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 332990 197865 333310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 332990 299865 333310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 332990 401865 333310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 332990 503865 333310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 341990 1928 342310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 341990 197865 342310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 341990 299865 342310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 341990 401865 342310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 341990 503865 342310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 350990 1928 351310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 359990 1928 360310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 359990 150409 360310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 359990 252409 360310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 359990 354409 360310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 359990 457089 360310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 368990 1928 369310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 368990 95225 369310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 368990 150409 369310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 368990 252409 369310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 368990 354409 369310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 368990 457089 369310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 377990 1928 378310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 377990 95225 378310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 377990 150409 378310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 377990 252409 378310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 377990 354409 378310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 377990 457089 378310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 386990 1928 387310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 386990 95225 387310 110999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 386990 150409 387310 212999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 386990 252409 387310 314999 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 386990 354409 387310 418903 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 386990 457089 387310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 395990 1928 396310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 395990 95225 396310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 404990 1928 405310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 1928 414310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 93865 414310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 197865 414310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 299865 414310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 401865 414310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 454137 414310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 413990 503865 414310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 1928 423310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 93865 423310 126543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 147865 423310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 197865 423310 229143 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 250465 423310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 299865 423310 330543 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 351865 423310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 401865 423310 419351 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 454137 423310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 422990 503865 423310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 431990 1928 432310 56359 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 431990 93865 432310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 431990 197865 432310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 431990 299865 432310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 431990 401865 432310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 431990 503865 432310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 440990 1928 441310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 440990 197865 441310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 440990 299865 441310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 440990 401865 441310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 440990 503865 441310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 1928 450310 5868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 45444 450310 160767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 197865 450310 262767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 299865 450310 364767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 401865 450310 466767 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 503865 450310 521868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 449990 561444 450310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 458990 1928 459310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 467990 1928 468310 56087 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 467990 80537 468310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 1928 477310 56087 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 80537 477310 101951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 129665 477310 155399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 186649 477310 203951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 231665 477310 257399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 288649 477310 305951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 333665 477310 359399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 390649 477310 409719 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 441649 477310 461399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 476990 492649 477310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 1928 486310 101951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 129665 486310 155399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 186649 486310 203951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 231665 486310 257399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 288649 486310 305951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 333665 486310 359399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 390649 486310 409719 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 441649 486310 461399 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 485990 492649 486310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 1928 495310 101951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 129665 495310 152868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 192444 495310 203951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 231665 495310 254868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 294444 495310 305951 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 333665 495310 356868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 396444 495310 458868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 494990 498444 495310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 503990 1928 504310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 512990 1928 513310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 521990 1928 522310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 530990 1928 531310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 539990 1928 540310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 548990 1928 549310 155868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 548990 195444 549310 257868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 548990 297444 549310 359868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 548990 399444 549310 461868 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 548990 501444 549310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 557990 1928 558310 587368 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 9876 560866 10196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 20876 560866 21196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 31876 560866 32196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 42876 560866 43196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 53876 560866 54196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 64876 560866 65196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 75876 560866 76196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 86876 560866 87196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 97876 560866 98196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 108876 560866 109196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 119876 560866 120196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 130876 560866 131196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 141876 560866 142196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 152876 560866 153196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 163876 560866 164196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 174876 560866 175196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 185876 560866 186196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 196876 560866 197196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 207876 560866 208196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 218876 560866 219196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 229876 560866 230196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 240876 560866 241196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 251876 560866 252196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 262876 560866 263196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 273876 560866 274196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 284876 560866 285196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 295876 560866 296196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 306876 560866 307196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 317876 560866 318196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 328876 560866 329196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 339876 560866 340196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 350876 560866 351196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 361876 560866 362196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 372876 560866 373196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 383876 560866 384196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 394876 560866 395196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 405876 560866 406196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 416876 560866 417196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 427876 560866 428196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 438876 560866 439196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 449876 560866 450196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 460876 560866 461196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 471876 560866 472196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 482876 560866 483196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 493876 560866 494196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 504876 560866 505196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 515876 560866 516196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 526876 560866 527196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 537876 560866 538196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 548876 560866 549196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 559876 560866 560196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 570876 560866 571196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal5 s 1042 581876 560866 582196 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 3230 104744 3550 150536 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 103142 209192 103462 254440 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 302230 156968 302550 202760 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 355222 258696 355542 304488 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 454766 353896 455086 356712 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 3230 207016 3550 252808 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 101670 106920 101990 152712 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 302230 258696 302550 304488 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 3230 308744 3550 354536 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 101670 413192 101990 458440 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 302230 360968 302550 406760 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 355222 156968 355542 202760 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 454766 252168 455086 255528 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 3230 411016 3550 456808 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 101670 310920 101990 356712 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 302230 462696 302550 508488 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 355222 360968 355542 406760 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 454766 149896 455086 152712 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 355222 462696 355542 508488 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 456238 156968 456558 195688 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 456238 258696 456558 297416 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 456238 462696 456558 501416 6 vssd1
port 137 nsew signal bidirectional
rlabel metal4 s 456238 360968 456558 399688 6 vssd1
port 137 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 561786 589600
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 104779648
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/fpga_top/runs/23_01_20_11_39/results/signoff/fpga_top.magic.gds
string GDS_START 37707536
<< end >>

