VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_right
  CLASS BLOCK ;
  FOREIGN grid_io_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 115.640 199.000 116.240 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 1.000 51.890 4.000 ;
    END
  END ccff_tail
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 163.240 4.000 163.840 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 27.240 4.000 27.840 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 1.000 154.930 4.000 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 81.640 4.000 82.240 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 54.440 4.000 55.040 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 199.000 61.840 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 196.000 67.990 199.000 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN left_width_0_height_0_subtile_0__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 196.000 171.030 199.000 ;
    END
  END left_width_0_height_0_subtile_0__pin_inpad_0_
  PIN left_width_0_height_0_subtile_0__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 196.000 196.790 199.000 ;
    END
  END left_width_0_height_0_subtile_0__pin_outpad_0_
  PIN left_width_0_height_0_subtile_1__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 196.000 145.270 199.000 ;
    END
  END left_width_0_height_0_subtile_1__pin_inpad_0_
  PIN left_width_0_height_0_subtile_1__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 199.000 7.440 ;
    END
  END left_width_0_height_0_subtile_1__pin_outpad_0_
  PIN left_width_0_height_0_subtile_2__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1.000 129.170 4.000 ;
    END
  END left_width_0_height_0_subtile_2__pin_inpad_0_
  PIN left_width_0_height_0_subtile_2__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 196.000 16.470 199.000 ;
    END
  END left_width_0_height_0_subtile_2__pin_outpad_0_
  PIN left_width_0_height_0_subtile_3__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1.000 180.690 4.000 ;
    END
  END left_width_0_height_0_subtile_3__pin_inpad_0_
  PIN left_width_0_height_0_subtile_3__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 196.000 119.510 199.000 ;
    END
  END left_width_0_height_0_subtile_3__pin_outpad_0_
  PIN left_width_0_height_0_subtile_4__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1.000 26.130 4.000 ;
    END
  END left_width_0_height_0_subtile_4__pin_inpad_0_
  PIN left_width_0_height_0_subtile_4__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 196.000 42.230 199.000 ;
    END
  END left_width_0_height_0_subtile_4__pin_outpad_0_
  PIN left_width_0_height_0_subtile_5__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.040 199.000 34.640 ;
    END
  END left_width_0_height_0_subtile_5__pin_inpad_0_
  PIN left_width_0_height_0_subtile_5__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1.000 77.650 4.000 ;
    END
  END left_width_0_height_0_subtile_5__pin_outpad_0_
  PIN left_width_0_height_0_subtile_6__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 142.840 199.000 143.440 ;
    END
  END left_width_0_height_0_subtile_6__pin_inpad_0_
  PIN left_width_0_height_0_subtile_6__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.040 199.000 170.640 ;
    END
  END left_width_0_height_0_subtile_6__pin_outpad_0_
  PIN left_width_0_height_0_subtile_7__pin_inpad_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 136.040 4.000 136.640 ;
    END
  END left_width_0_height_0_subtile_7__pin_inpad_0_
  PIN left_width_0_height_0_subtile_7__pin_outpad_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 196.000 93.750 199.000 ;
    END
  END left_width_0_height_0_subtile_7__pin_outpad_0_
  PIN pReset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1.000 103.410 4.000 ;
    END
  END pReset
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 108.840 4.000 109.440 ;
    END
  END prog_clk
  PIN vccd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.440 4.000 191.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 199.000 89.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 0.070 6.500 196.810 187.920 ;
      LAYER met2 ;
        RECT 0.100 195.720 15.910 196.000 ;
        RECT 16.750 195.720 41.670 196.000 ;
        RECT 42.510 195.720 67.430 196.000 ;
        RECT 68.270 195.720 93.190 196.000 ;
        RECT 94.030 195.720 118.950 196.000 ;
        RECT 119.790 195.720 144.710 196.000 ;
        RECT 145.550 195.720 170.470 196.000 ;
        RECT 171.310 195.720 196.230 196.000 ;
        RECT 0.100 4.280 196.780 195.720 ;
        RECT 0.650 3.670 25.570 4.280 ;
        RECT 26.410 3.670 51.330 4.280 ;
        RECT 52.170 3.670 77.090 4.280 ;
        RECT 77.930 3.670 102.850 4.280 ;
        RECT 103.690 3.670 128.610 4.280 ;
        RECT 129.450 3.670 154.370 4.280 ;
        RECT 155.210 3.670 180.130 4.280 ;
        RECT 180.970 3.670 196.780 4.280 ;
      LAYER met3 ;
        RECT 4.000 171.040 196.000 187.845 ;
        RECT 4.000 169.640 195.600 171.040 ;
        RECT 4.000 164.240 196.000 169.640 ;
        RECT 4.400 162.840 196.000 164.240 ;
        RECT 4.000 143.840 196.000 162.840 ;
        RECT 4.000 142.440 195.600 143.840 ;
        RECT 4.000 137.040 196.000 142.440 ;
        RECT 4.400 135.640 196.000 137.040 ;
        RECT 4.000 116.640 196.000 135.640 ;
        RECT 4.000 115.240 195.600 116.640 ;
        RECT 4.000 109.840 196.000 115.240 ;
        RECT 4.400 108.440 196.000 109.840 ;
        RECT 4.000 89.440 196.000 108.440 ;
        RECT 4.000 88.040 195.600 89.440 ;
        RECT 4.000 82.640 196.000 88.040 ;
        RECT 4.400 81.240 196.000 82.640 ;
        RECT 4.000 62.240 196.000 81.240 ;
        RECT 4.000 60.840 195.600 62.240 ;
        RECT 4.000 55.440 196.000 60.840 ;
        RECT 4.400 54.040 196.000 55.440 ;
        RECT 4.000 35.040 196.000 54.040 ;
        RECT 4.000 33.640 195.600 35.040 ;
        RECT 4.000 28.240 196.000 33.640 ;
        RECT 4.400 26.840 196.000 28.240 ;
        RECT 4.000 7.840 196.000 26.840 ;
        RECT 4.000 6.975 195.600 7.840 ;
  END
END grid_io_right
END LIBRARY

