magic
tech sky130A
magscale 1 2
timestamp 1674175171
<< viali >>
rect 3157 37349 3191 37383
rect 17141 37349 17175 37383
rect 1593 37281 1627 37315
rect 3985 37281 4019 37315
rect 6561 37281 6595 37315
rect 9137 37281 9171 37315
rect 22661 37281 22695 37315
rect 24869 37281 24903 37315
rect 27813 37281 27847 37315
rect 1869 37213 1903 37247
rect 2973 37213 3007 37247
rect 4261 37213 4295 37247
rect 5457 37213 5491 37247
rect 6837 37213 6871 37247
rect 8033 37213 8067 37247
rect 9413 37213 9447 37247
rect 10425 37213 10459 37247
rect 11897 37213 11931 37247
rect 12541 37213 12575 37247
rect 14289 37213 14323 37247
rect 14657 37213 14691 37247
rect 14933 37213 14967 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 22201 37213 22235 37247
rect 22937 37213 22971 37247
rect 24685 37213 24719 37247
rect 25881 37213 25915 37247
rect 26341 37213 26375 37247
rect 28089 37213 28123 37247
rect 29929 37213 29963 37247
rect 30573 37213 30607 37247
rect 31033 37213 31067 37247
rect 32321 37213 32355 37247
rect 33057 37213 33091 37247
rect 34897 37213 34931 37247
rect 36185 37213 36219 37247
rect 37473 37213 37507 37247
rect 16957 37145 16991 37179
rect 5273 37077 5307 37111
rect 7849 37077 7883 37111
rect 10609 37077 10643 37111
rect 11713 37077 11747 37111
rect 12357 37077 12391 37111
rect 14105 37077 14139 37111
rect 15117 37077 15151 37111
rect 18153 37077 18187 37111
rect 20269 37077 20303 37111
rect 22017 37077 22051 37111
rect 25697 37077 25731 37111
rect 26525 37077 26559 37111
rect 29745 37077 29779 37111
rect 30389 37077 30423 37111
rect 31217 37077 31251 37111
rect 32505 37077 32539 37111
rect 33241 37077 33275 37111
rect 35081 37077 35115 37111
rect 36369 37077 36403 37111
rect 37657 37077 37691 37111
rect 1777 36873 1811 36907
rect 17693 36873 17727 36907
rect 19625 36873 19659 36907
rect 29193 36873 29227 36907
rect 31401 36873 31435 36907
rect 38117 36805 38151 36839
rect 1593 36737 1627 36771
rect 2513 36737 2547 36771
rect 3157 36737 3191 36771
rect 9321 36737 9355 36771
rect 13185 36737 13219 36771
rect 17049 36737 17083 36771
rect 17877 36737 17911 36771
rect 19441 36737 19475 36771
rect 23489 36737 23523 36771
rect 28457 36737 28491 36771
rect 28733 36737 28767 36771
rect 29377 36737 29411 36771
rect 31585 36737 31619 36771
rect 35725 36737 35759 36771
rect 36369 36737 36403 36771
rect 2329 36601 2363 36635
rect 13001 36601 13035 36635
rect 2973 36533 3007 36567
rect 9137 36533 9171 36567
rect 16865 36533 16899 36567
rect 23305 36533 23339 36567
rect 35541 36533 35575 36567
rect 36461 36533 36495 36567
rect 38209 36533 38243 36567
rect 37473 36329 37507 36363
rect 36645 36261 36679 36295
rect 1777 36125 1811 36159
rect 36829 36125 36863 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 1593 35989 1627 36023
rect 38209 35989 38243 36023
rect 12541 35785 12575 35819
rect 1777 35649 1811 35683
rect 12725 35649 12759 35683
rect 36921 35649 36955 35683
rect 38025 35649 38059 35683
rect 1593 35445 1627 35479
rect 36737 35445 36771 35479
rect 38209 35445 38243 35479
rect 38301 35037 38335 35071
rect 38117 34901 38151 34935
rect 1593 34561 1627 34595
rect 38025 34561 38059 34595
rect 1777 34357 1811 34391
rect 38209 34357 38243 34391
rect 4537 33609 4571 33643
rect 4721 33473 4755 33507
rect 28181 33065 28215 33099
rect 37381 33065 37415 33099
rect 1593 32861 1627 32895
rect 4169 32861 4203 32895
rect 28365 32861 28399 32895
rect 37565 32861 37599 32895
rect 38117 32793 38151 32827
rect 1777 32725 1811 32759
rect 3985 32725 4019 32759
rect 38209 32725 38243 32759
rect 13921 32521 13955 32555
rect 36829 32521 36863 32555
rect 1593 32385 1627 32419
rect 13829 32385 13863 32419
rect 15301 32385 15335 32419
rect 36737 32385 36771 32419
rect 38117 32385 38151 32419
rect 1777 32181 1811 32215
rect 15393 32181 15427 32215
rect 38209 32181 38243 32215
rect 23029 31977 23063 32011
rect 5917 31841 5951 31875
rect 19625 31841 19659 31875
rect 21741 31841 21775 31875
rect 5825 31773 5859 31807
rect 19533 31773 19567 31807
rect 20637 31773 20671 31807
rect 20821 31773 20855 31807
rect 21649 31773 21683 31807
rect 22937 31773 22971 31807
rect 26709 31773 26743 31807
rect 26525 31637 26559 31671
rect 33333 31433 33367 31467
rect 5733 31297 5767 31331
rect 25697 31297 25731 31331
rect 33517 31297 33551 31331
rect 5825 31093 5859 31127
rect 25789 31093 25823 31127
rect 1593 30685 1627 30719
rect 6837 30685 6871 30719
rect 8033 30685 8067 30719
rect 11069 30685 11103 30719
rect 29745 30685 29779 30719
rect 30481 30685 30515 30719
rect 38025 30685 38059 30719
rect 6929 30617 6963 30651
rect 30573 30617 30607 30651
rect 1777 30549 1811 30583
rect 8125 30549 8159 30583
rect 11161 30549 11195 30583
rect 29837 30549 29871 30583
rect 38209 30549 38243 30583
rect 6653 30277 6687 30311
rect 3893 30209 3927 30243
rect 6561 30209 6595 30243
rect 13277 30209 13311 30243
rect 25421 30209 25455 30243
rect 27169 30209 27203 30243
rect 3709 30073 3743 30107
rect 13093 30073 13127 30107
rect 25237 30073 25271 30107
rect 27261 30005 27295 30039
rect 33793 29801 33827 29835
rect 1777 29597 1811 29631
rect 7849 29597 7883 29631
rect 10609 29597 10643 29631
rect 33977 29597 34011 29631
rect 38025 29597 38059 29631
rect 1593 29461 1627 29495
rect 7941 29461 7975 29495
rect 10701 29461 10735 29495
rect 38209 29461 38243 29495
rect 1593 29121 1627 29155
rect 14565 29121 14599 29155
rect 15485 29121 15519 29155
rect 38025 29121 38059 29155
rect 14657 29053 14691 29087
rect 1777 28985 1811 29019
rect 15577 28985 15611 29019
rect 38209 28985 38243 29019
rect 11897 28509 11931 28543
rect 18061 28509 18095 28543
rect 11989 28373 12023 28407
rect 18153 28373 18187 28407
rect 35081 28169 35115 28203
rect 15209 28033 15243 28067
rect 23673 28033 23707 28067
rect 35265 28033 35299 28067
rect 15301 27829 15335 27863
rect 23765 27829 23799 27863
rect 1777 27421 1811 27455
rect 38301 27421 38335 27455
rect 1593 27285 1627 27319
rect 38117 27285 38151 27319
rect 6837 27081 6871 27115
rect 35357 27081 35391 27115
rect 6745 26945 6779 26979
rect 13001 26945 13035 26979
rect 13645 26945 13679 26979
rect 22109 26945 22143 26979
rect 35265 26945 35299 26979
rect 22293 26809 22327 26843
rect 12817 26741 12851 26775
rect 13461 26741 13495 26775
rect 34897 26537 34931 26571
rect 1593 26469 1627 26503
rect 13553 26469 13587 26503
rect 15025 26469 15059 26503
rect 15669 26469 15703 26503
rect 1777 26333 1811 26367
rect 12173 26333 12207 26367
rect 13737 26333 13771 26367
rect 14289 26333 14323 26367
rect 15209 26333 15243 26367
rect 15853 26333 15887 26367
rect 18061 26333 18095 26367
rect 35081 26333 35115 26367
rect 38301 26333 38335 26367
rect 12265 26265 12299 26299
rect 14381 26265 14415 26299
rect 17877 26197 17911 26231
rect 38117 26197 38151 26231
rect 28089 25993 28123 26027
rect 13737 25857 13771 25891
rect 17877 25857 17911 25891
rect 18889 25857 18923 25891
rect 27997 25857 28031 25891
rect 13553 25653 13587 25687
rect 17969 25653 18003 25687
rect 18981 25653 19015 25687
rect 28089 25449 28123 25483
rect 14289 25245 14323 25279
rect 15485 25245 15519 25279
rect 16129 25245 16163 25279
rect 17233 25245 17267 25279
rect 27997 25245 28031 25279
rect 38025 25245 38059 25279
rect 18245 25177 18279 25211
rect 18337 25177 18371 25211
rect 18889 25177 18923 25211
rect 14381 25109 14415 25143
rect 15577 25109 15611 25143
rect 16221 25109 16255 25143
rect 17049 25109 17083 25143
rect 38209 25109 38243 25143
rect 14381 24837 14415 24871
rect 17049 24837 17083 24871
rect 1593 24769 1627 24803
rect 7389 24769 7423 24803
rect 9229 24769 9263 24803
rect 14933 24769 14967 24803
rect 15485 24769 15519 24803
rect 16129 24769 16163 24803
rect 22753 24769 22787 24803
rect 23397 24769 23431 24803
rect 13553 24701 13587 24735
rect 14289 24701 14323 24735
rect 16957 24701 16991 24735
rect 7481 24633 7515 24667
rect 17509 24633 17543 24667
rect 22569 24633 22603 24667
rect 1777 24565 1811 24599
rect 9045 24565 9079 24599
rect 15577 24565 15611 24599
rect 16221 24565 16255 24599
rect 23213 24565 23247 24599
rect 10701 24293 10735 24327
rect 15853 24293 15887 24327
rect 12265 24225 12299 24259
rect 15025 24225 15059 24259
rect 15485 24225 15519 24259
rect 15669 24225 15703 24259
rect 16773 24225 16807 24259
rect 16957 24225 16991 24259
rect 20545 24225 20579 24259
rect 1593 24157 1627 24191
rect 9321 24157 9355 24191
rect 10149 24157 10183 24191
rect 10609 24157 10643 24191
rect 11253 24157 11287 24191
rect 17417 24157 17451 24191
rect 18429 24157 18463 24191
rect 37473 24157 37507 24191
rect 37749 24157 37783 24191
rect 12357 24089 12391 24123
rect 13277 24089 13311 24123
rect 14381 24089 14415 24123
rect 14473 24089 14507 24123
rect 19533 24089 19567 24123
rect 19625 24089 19659 24123
rect 1777 24021 1811 24055
rect 9413 24021 9447 24055
rect 9965 24021 9999 24055
rect 11345 24021 11379 24055
rect 18521 24021 18555 24055
rect 22661 24021 22695 24055
rect 22109 23817 22143 23851
rect 30757 23817 30791 23851
rect 10425 23749 10459 23783
rect 10977 23749 11011 23783
rect 15117 23749 15151 23783
rect 17141 23749 17175 23783
rect 17877 23749 17911 23783
rect 7573 23681 7607 23715
rect 8401 23681 8435 23715
rect 13829 23681 13863 23715
rect 14013 23681 14047 23715
rect 16129 23681 16163 23715
rect 17049 23681 17083 23715
rect 18889 23681 18923 23715
rect 22017 23681 22051 23715
rect 22661 23681 22695 23715
rect 22845 23681 22879 23715
rect 25789 23681 25823 23715
rect 30665 23681 30699 23715
rect 10333 23613 10367 23647
rect 12725 23613 12759 23647
rect 12909 23613 12943 23647
rect 15025 23613 15059 23647
rect 17785 23613 17819 23647
rect 18061 23613 18095 23647
rect 7665 23545 7699 23579
rect 13369 23545 13403 23579
rect 14197 23545 14231 23579
rect 15577 23545 15611 23579
rect 8217 23477 8251 23511
rect 16221 23477 16255 23511
rect 18981 23477 19015 23511
rect 23029 23477 23063 23511
rect 25605 23477 25639 23511
rect 8401 23205 8435 23239
rect 16037 23205 16071 23239
rect 10793 23137 10827 23171
rect 12265 23137 12299 23171
rect 18245 23137 18279 23171
rect 18521 23137 18555 23171
rect 7757 23069 7791 23103
rect 8585 23069 8619 23103
rect 9137 23069 9171 23103
rect 10701 23069 10735 23103
rect 12081 23069 12115 23103
rect 20177 23069 20211 23103
rect 21097 23069 21131 23103
rect 21649 23069 21683 23103
rect 7849 23001 7883 23035
rect 15853 23001 15887 23035
rect 18337 23001 18371 23035
rect 9229 22933 9263 22967
rect 12725 22933 12759 22967
rect 13185 22933 13219 22967
rect 14749 22933 14783 22967
rect 20269 22933 20303 22967
rect 20913 22933 20947 22967
rect 21741 22933 21775 22967
rect 2329 22729 2363 22763
rect 8401 22729 8435 22763
rect 14381 22729 14415 22763
rect 20269 22729 20303 22763
rect 29193 22729 29227 22763
rect 10609 22661 10643 22695
rect 15761 22661 15795 22695
rect 17141 22661 17175 22695
rect 17693 22661 17727 22695
rect 23489 22661 23523 22695
rect 25053 22661 25087 22695
rect 1685 22593 1719 22627
rect 2513 22593 2547 22627
rect 7205 22593 7239 22627
rect 8309 22593 8343 22627
rect 9137 22593 9171 22627
rect 9781 22593 9815 22627
rect 12081 22593 12115 22627
rect 13645 22593 13679 22627
rect 14289 22593 14323 22627
rect 14933 22593 14967 22627
rect 19809 22593 19843 22627
rect 20913 22593 20947 22627
rect 22201 22593 22235 22627
rect 29101 22593 29135 22627
rect 38025 22593 38059 22627
rect 10517 22525 10551 22559
rect 12265 22525 12299 22559
rect 15669 22525 15703 22559
rect 15945 22525 15979 22559
rect 17049 22525 17083 22559
rect 19625 22525 19659 22559
rect 23397 22525 23431 22559
rect 24317 22525 24351 22559
rect 24961 22525 24995 22559
rect 25237 22525 25271 22559
rect 9229 22457 9263 22491
rect 11069 22457 11103 22491
rect 12449 22457 12483 22491
rect 38209 22457 38243 22491
rect 1777 22389 1811 22423
rect 7021 22389 7055 22423
rect 9873 22389 9907 22423
rect 13737 22389 13771 22423
rect 15025 22389 15059 22423
rect 21005 22389 21039 22423
rect 22017 22389 22051 22423
rect 13185 22185 13219 22219
rect 12817 22049 12851 22083
rect 14749 22049 14783 22083
rect 15761 22049 15795 22083
rect 18245 22049 18279 22083
rect 18521 22049 18555 22083
rect 19533 22049 19567 22083
rect 20177 22049 20211 22083
rect 21373 22049 21407 22083
rect 23305 22049 23339 22083
rect 1961 21981 1995 22015
rect 7297 21981 7331 22015
rect 12173 21981 12207 22015
rect 13001 21981 13035 22015
rect 23949 21981 23983 22015
rect 31493 21981 31527 22015
rect 38301 21981 38335 22015
rect 10701 21913 10735 21947
rect 10793 21913 10827 21947
rect 11713 21913 11747 21947
rect 14841 21913 14875 21947
rect 16313 21913 16347 21947
rect 16405 21913 16439 21947
rect 16957 21913 16991 21947
rect 18337 21913 18371 21947
rect 19618 21913 19652 21947
rect 21097 21913 21131 21947
rect 21189 21913 21223 21947
rect 22661 21913 22695 21947
rect 22753 21913 22787 21947
rect 1777 21845 1811 21879
rect 7113 21845 7147 21879
rect 12265 21845 12299 21879
rect 23765 21845 23799 21879
rect 31585 21845 31619 21879
rect 38117 21845 38151 21879
rect 11161 21641 11195 21675
rect 17509 21641 17543 21675
rect 22017 21641 22051 21675
rect 22661 21641 22695 21675
rect 12357 21573 12391 21607
rect 13737 21573 13771 21607
rect 13829 21573 13863 21607
rect 15301 21573 15335 21607
rect 16221 21573 16255 21607
rect 20085 21573 20119 21607
rect 21189 21573 21223 21607
rect 27537 21573 27571 21607
rect 27629 21573 27663 21607
rect 1593 21505 1627 21539
rect 7205 21505 7239 21539
rect 8493 21505 8527 21539
rect 9137 21505 9171 21539
rect 10701 21505 10735 21539
rect 16857 21503 16891 21537
rect 17693 21505 17727 21539
rect 18613 21505 18647 21539
rect 21097 21505 21131 21539
rect 23397 21505 23431 21539
rect 23581 21505 23615 21539
rect 24593 21505 24627 21539
rect 25513 21505 25547 21539
rect 31217 21505 31251 21539
rect 9229 21437 9263 21471
rect 10517 21437 10551 21471
rect 12265 21437 12299 21471
rect 12541 21437 12575 21471
rect 15209 21437 15243 21471
rect 19257 21437 19291 21471
rect 19993 21437 20027 21471
rect 20269 21437 20303 21471
rect 28549 21437 28583 21471
rect 14289 21369 14323 21403
rect 25605 21369 25639 21403
rect 1777 21301 1811 21335
rect 7297 21301 7331 21335
rect 8585 21301 8619 21335
rect 16957 21301 16991 21335
rect 18705 21301 18739 21335
rect 24041 21301 24075 21335
rect 24685 21301 24719 21335
rect 31309 21301 31343 21335
rect 1593 21097 1627 21131
rect 8493 21097 8527 21131
rect 24593 21097 24627 21131
rect 6653 21029 6687 21063
rect 13645 21029 13679 21063
rect 20085 21029 20119 21063
rect 27721 21029 27755 21063
rect 12357 20961 12391 20995
rect 13093 20961 13127 20995
rect 13277 20961 13311 20995
rect 14565 20961 14599 20995
rect 14749 20961 14783 20995
rect 15853 20961 15887 20995
rect 16865 20961 16899 20995
rect 17417 20961 17451 20995
rect 19533 20961 19567 20995
rect 20729 20961 20763 20995
rect 20913 20961 20947 20995
rect 1777 20893 1811 20927
rect 7389 20893 7423 20927
rect 8401 20893 8435 20927
rect 9689 20893 9723 20927
rect 15209 20893 15243 20927
rect 22937 20893 22971 20927
rect 23121 20893 23155 20927
rect 24777 20893 24811 20927
rect 26801 20893 26835 20927
rect 26893 20893 26927 20927
rect 33977 20893 34011 20927
rect 38025 20893 38059 20927
rect 6101 20825 6135 20859
rect 6193 20825 6227 20859
rect 10425 20825 10459 20859
rect 10517 20825 10551 20859
rect 11437 20825 11471 20859
rect 15945 20825 15979 20859
rect 17509 20825 17543 20859
rect 18429 20825 18463 20859
rect 19625 20825 19659 20859
rect 23581 20825 23615 20859
rect 27537 20825 27571 20859
rect 7205 20757 7239 20791
rect 9781 20757 9815 20791
rect 21373 20757 21407 20791
rect 33793 20757 33827 20791
rect 38209 20757 38243 20791
rect 12173 20553 12207 20587
rect 12817 20553 12851 20587
rect 17049 20553 17083 20587
rect 24133 20553 24167 20587
rect 7021 20485 7055 20519
rect 7113 20485 7147 20519
rect 8677 20485 8711 20519
rect 10333 20485 10367 20519
rect 10885 20485 10919 20519
rect 14749 20485 14783 20519
rect 15301 20485 15335 20519
rect 17693 20485 17727 20519
rect 20085 20485 20119 20519
rect 23397 20485 23431 20519
rect 12081 20417 12115 20451
rect 12725 20417 12759 20451
rect 13461 20417 13495 20451
rect 15761 20417 15795 20451
rect 16957 20417 16991 20451
rect 17601 20417 17635 20451
rect 19165 20417 19199 20451
rect 21281 20417 21315 20451
rect 24041 20417 24075 20451
rect 29193 20417 29227 20451
rect 33977 20417 34011 20451
rect 8033 20349 8067 20383
rect 8585 20349 8619 20383
rect 8861 20349 8895 20383
rect 10241 20349 10275 20383
rect 14657 20349 14691 20383
rect 19993 20349 20027 20383
rect 20545 20281 20579 20315
rect 23581 20281 23615 20315
rect 13553 20213 13587 20247
rect 15853 20213 15887 20247
rect 19257 20213 19291 20247
rect 21097 20213 21131 20247
rect 29009 20213 29043 20247
rect 33793 20213 33827 20247
rect 8033 20009 8067 20043
rect 16589 20009 16623 20043
rect 19533 20009 19567 20043
rect 20821 20009 20855 20043
rect 9229 19941 9263 19975
rect 12081 19941 12115 19975
rect 21281 19941 21315 19975
rect 27077 19941 27111 19975
rect 10241 19873 10275 19907
rect 12725 19873 12759 19907
rect 13737 19873 13771 19907
rect 15025 19873 15059 19907
rect 16129 19873 16163 19907
rect 16313 19873 16347 19907
rect 20177 19873 20211 19907
rect 20361 19873 20395 19907
rect 26893 19873 26927 19907
rect 28549 19873 28583 19907
rect 7941 19805 7975 19839
rect 9137 19805 9171 19839
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 14289 19805 14323 19839
rect 15669 19805 15703 19839
rect 19441 19805 19475 19839
rect 21465 19805 21499 19839
rect 22661 19805 22695 19839
rect 26709 19805 26743 19839
rect 27813 19805 27847 19839
rect 28457 19805 28491 19839
rect 30849 19805 30883 19839
rect 6837 19737 6871 19771
rect 6929 19737 6963 19771
rect 7481 19737 7515 19771
rect 11529 19737 11563 19771
rect 11621 19737 11655 19771
rect 12817 19737 12851 19771
rect 15117 19737 15151 19771
rect 17325 19737 17359 19771
rect 17509 19737 17543 19771
rect 27905 19737 27939 19771
rect 10885 19669 10919 19703
rect 14381 19669 14415 19703
rect 22477 19669 22511 19703
rect 30941 19669 30975 19703
rect 1593 19465 1627 19499
rect 5825 19465 5859 19499
rect 7757 19465 7791 19499
rect 9137 19465 9171 19499
rect 9781 19465 9815 19499
rect 12173 19397 12207 19431
rect 13737 19397 13771 19431
rect 14657 19397 14691 19431
rect 15209 19397 15243 19431
rect 15301 19397 15335 19431
rect 16221 19397 16255 19431
rect 17969 19397 18003 19431
rect 1777 19329 1811 19363
rect 4813 19329 4847 19363
rect 6009 19329 6043 19363
rect 7113 19329 7147 19363
rect 7205 19329 7239 19363
rect 7941 19329 7975 19363
rect 9045 19329 9079 19363
rect 9689 19329 9723 19363
rect 10425 19329 10459 19363
rect 10517 19329 10551 19363
rect 16957 19329 16991 19363
rect 22017 19329 22051 19363
rect 28733 19329 28767 19363
rect 30113 19329 30147 19363
rect 30205 19329 30239 19363
rect 38117 19329 38151 19363
rect 8401 19261 8435 19295
rect 12081 19261 12115 19295
rect 13093 19261 13127 19295
rect 13645 19261 13679 19295
rect 17877 19261 17911 19295
rect 18245 19261 18279 19295
rect 19441 19261 19475 19295
rect 4629 19125 4663 19159
rect 17049 19125 17083 19159
rect 22109 19125 22143 19159
rect 28549 19125 28583 19159
rect 38209 19125 38243 19159
rect 6469 18921 6503 18955
rect 7849 18921 7883 18955
rect 9229 18785 9263 18819
rect 9505 18785 9539 18819
rect 10701 18785 10735 18819
rect 11069 18785 11103 18819
rect 12725 18785 12759 18819
rect 13645 18785 13679 18819
rect 15025 18785 15059 18819
rect 19533 18785 19567 18819
rect 19809 18785 19843 18819
rect 22477 18785 22511 18819
rect 4721 18717 4755 18751
rect 6009 18717 6043 18751
rect 6653 18717 6687 18751
rect 7113 18717 7147 18751
rect 7757 18717 7791 18751
rect 8401 18717 8435 18751
rect 11989 18717 12023 18751
rect 14829 18717 14863 18751
rect 16037 18717 16071 18751
rect 16681 18717 16715 18751
rect 17509 18717 17543 18751
rect 18705 18717 18739 18751
rect 21189 18717 21223 18751
rect 23765 18717 23799 18751
rect 24777 18717 24811 18751
rect 25421 18717 25455 18751
rect 26157 18717 26191 18751
rect 27261 18717 27295 18751
rect 9321 18649 9355 18683
rect 10793 18649 10827 18683
rect 12081 18649 12115 18683
rect 12817 18649 12851 18683
rect 18797 18649 18831 18683
rect 19625 18649 19659 18683
rect 22569 18649 22603 18683
rect 23121 18649 23155 18683
rect 4537 18581 4571 18615
rect 5825 18581 5859 18615
rect 7205 18581 7239 18615
rect 8493 18581 8527 18615
rect 15485 18581 15519 18615
rect 16129 18581 16163 18615
rect 16773 18581 16807 18615
rect 17601 18581 17635 18615
rect 21281 18581 21315 18615
rect 23581 18581 23615 18615
rect 24869 18581 24903 18615
rect 25513 18581 25547 18615
rect 26249 18581 26283 18615
rect 27077 18581 27111 18615
rect 28089 18581 28123 18615
rect 5825 18377 5859 18411
rect 8493 18377 8527 18411
rect 11805 18377 11839 18411
rect 13001 18377 13035 18411
rect 18521 18377 18555 18411
rect 21281 18377 21315 18411
rect 4353 18309 4387 18343
rect 9137 18309 9171 18343
rect 13645 18309 13679 18343
rect 14565 18309 14599 18343
rect 15754 18309 15788 18343
rect 17049 18309 17083 18343
rect 22201 18309 22235 18343
rect 24869 18309 24903 18343
rect 26065 18309 26099 18343
rect 27261 18309 27295 18343
rect 27353 18309 27387 18343
rect 1777 18241 1811 18275
rect 6009 18241 6043 18275
rect 7113 18241 7147 18275
rect 7757 18241 7791 18275
rect 8401 18241 8435 18275
rect 9045 18241 9079 18275
rect 9689 18241 9723 18275
rect 10517 18241 10551 18275
rect 10977 18241 11011 18275
rect 11713 18241 11747 18275
rect 12541 18241 12575 18275
rect 18429 18241 18463 18275
rect 19625 18241 19659 18275
rect 20453 18241 20487 18275
rect 21189 18241 21223 18275
rect 23765 18241 23799 18275
rect 28365 18241 28399 18275
rect 28549 18241 28583 18275
rect 4261 18173 4295 18207
rect 4905 18173 4939 18207
rect 12357 18173 12391 18207
rect 13553 18173 13587 18207
rect 15669 18173 15703 18207
rect 16957 18173 16991 18207
rect 17233 18173 17267 18207
rect 22109 18173 22143 18207
rect 23121 18173 23155 18207
rect 23581 18173 23615 18207
rect 24777 18173 24811 18207
rect 25053 18173 25087 18207
rect 25973 18173 26007 18207
rect 26617 18173 26651 18207
rect 7849 18105 7883 18139
rect 11069 18105 11103 18139
rect 16221 18105 16255 18139
rect 27813 18105 27847 18139
rect 1593 18037 1627 18071
rect 7205 18037 7239 18071
rect 9781 18037 9815 18071
rect 10333 18037 10367 18071
rect 19717 18037 19751 18071
rect 20545 18037 20579 18071
rect 24225 18037 24259 18071
rect 29009 18037 29043 18071
rect 7573 17833 7607 17867
rect 11713 17833 11747 17867
rect 14473 17833 14507 17867
rect 22845 17833 22879 17867
rect 25605 17833 25639 17867
rect 32137 17833 32171 17867
rect 13645 17765 13679 17799
rect 15669 17765 15703 17799
rect 4353 17697 4387 17731
rect 7389 17697 7423 17731
rect 10333 17697 10367 17731
rect 13093 17697 13127 17731
rect 17417 17697 17451 17731
rect 24869 17697 24903 17731
rect 26249 17697 26283 17731
rect 26893 17697 26927 17731
rect 5917 17629 5951 17663
rect 6561 17629 6595 17663
rect 7205 17629 7239 17663
rect 8401 17629 8435 17663
rect 10793 17629 10827 17663
rect 11897 17629 11931 17663
rect 12357 17629 12391 17663
rect 14381 17629 14415 17663
rect 16221 17629 16255 17663
rect 18521 17629 18555 17663
rect 19533 17629 19567 17663
rect 20545 17629 20579 17663
rect 22753 17629 22787 17663
rect 25513 17629 25547 17663
rect 27721 17629 27755 17663
rect 29745 17629 29779 17663
rect 32321 17629 32355 17663
rect 9689 17561 9723 17595
rect 9781 17561 9815 17595
rect 11069 17561 11103 17595
rect 13185 17561 13219 17595
rect 15117 17561 15151 17595
rect 15209 17561 15243 17595
rect 17509 17561 17543 17595
rect 18061 17561 18095 17595
rect 26341 17561 26375 17595
rect 6009 17493 6043 17527
rect 6653 17493 6687 17527
rect 8493 17493 8527 17527
rect 12449 17493 12483 17527
rect 16313 17493 16347 17527
rect 18613 17493 18647 17527
rect 19625 17493 19659 17527
rect 20637 17493 20671 17527
rect 27537 17493 27571 17527
rect 29837 17493 29871 17527
rect 25237 17289 25271 17323
rect 7481 17221 7515 17255
rect 9505 17221 9539 17255
rect 10609 17221 10643 17255
rect 11161 17221 11195 17255
rect 14381 17221 14415 17255
rect 15761 17221 15795 17255
rect 18061 17221 18095 17255
rect 19257 17221 19291 17255
rect 20453 17221 20487 17255
rect 23397 17221 23431 17255
rect 23489 17221 23523 17255
rect 25973 17221 26007 17255
rect 26065 17221 26099 17255
rect 27905 17221 27939 17255
rect 28457 17221 28491 17255
rect 1869 17153 1903 17187
rect 3525 17153 3559 17187
rect 4169 17153 4203 17187
rect 4997 17153 5031 17187
rect 5825 17153 5859 17187
rect 6653 17153 6687 17187
rect 8861 17153 8895 17187
rect 9045 17153 9079 17187
rect 11989 17153 12023 17187
rect 12633 17153 12667 17187
rect 13277 17153 13311 17187
rect 17233 17153 17267 17187
rect 24501 17153 24535 17187
rect 25145 17153 25179 17187
rect 29285 17153 29319 17187
rect 38301 17153 38335 17187
rect 1593 17085 1627 17119
rect 7389 17085 7423 17119
rect 10517 17085 10551 17119
rect 13461 17085 13495 17119
rect 14289 17085 14323 17119
rect 14565 17085 14599 17119
rect 15669 17085 15703 17119
rect 16313 17085 16347 17119
rect 17969 17085 18003 17119
rect 19165 17085 19199 17119
rect 20361 17085 20395 17119
rect 21005 17085 21039 17119
rect 24041 17085 24075 17119
rect 26617 17085 26651 17119
rect 27813 17085 27847 17119
rect 29101 17085 29135 17119
rect 5917 17017 5951 17051
rect 7941 17017 7975 17051
rect 12081 17017 12115 17051
rect 18521 17017 18555 17051
rect 19717 17017 19751 17051
rect 29469 17017 29503 17051
rect 3617 16949 3651 16983
rect 4261 16949 4295 16983
rect 4813 16949 4847 16983
rect 6745 16949 6779 16983
rect 12725 16949 12759 16983
rect 17325 16949 17359 16983
rect 24593 16949 24627 16983
rect 38117 16949 38151 16983
rect 18797 16745 18831 16779
rect 19809 16745 19843 16779
rect 26157 16745 26191 16779
rect 10241 16677 10275 16711
rect 13461 16677 13495 16711
rect 29837 16677 29871 16711
rect 9689 16609 9723 16643
rect 11529 16609 11563 16643
rect 11805 16609 11839 16643
rect 12909 16609 12943 16643
rect 15117 16609 15151 16643
rect 20545 16609 20579 16643
rect 20821 16609 20855 16643
rect 3249 16541 3283 16575
rect 4537 16541 4571 16575
rect 5181 16541 5215 16575
rect 5825 16541 5859 16575
rect 6469 16541 6503 16575
rect 7113 16541 7147 16575
rect 7757 16541 7791 16575
rect 7849 16541 7883 16575
rect 8401 16541 8435 16575
rect 10793 16541 10827 16575
rect 14381 16541 14415 16575
rect 16773 16541 16807 16575
rect 17417 16541 17451 16575
rect 18245 16541 18279 16575
rect 18705 16541 18739 16575
rect 19717 16541 19751 16575
rect 23489 16541 23523 16575
rect 24593 16541 24627 16575
rect 26065 16541 26099 16575
rect 27169 16541 27203 16575
rect 29745 16541 29779 16575
rect 7205 16473 7239 16507
rect 9781 16473 9815 16507
rect 11621 16473 11655 16507
rect 13001 16473 13035 16507
rect 15209 16473 15243 16507
rect 16129 16473 16163 16507
rect 16865 16473 16899 16507
rect 20637 16473 20671 16507
rect 21741 16473 21775 16507
rect 21833 16473 21867 16507
rect 22385 16473 22419 16507
rect 24685 16473 24719 16507
rect 2421 16405 2455 16439
rect 3065 16405 3099 16439
rect 4629 16405 4663 16439
rect 5273 16405 5307 16439
rect 5917 16405 5951 16439
rect 6561 16405 6595 16439
rect 8493 16405 8527 16439
rect 10885 16405 10919 16439
rect 14473 16405 14507 16439
rect 17509 16405 17543 16439
rect 18061 16405 18095 16439
rect 22845 16405 22879 16439
rect 23581 16405 23615 16439
rect 27261 16405 27295 16439
rect 2697 16201 2731 16235
rect 8309 16201 8343 16235
rect 16221 16201 16255 16235
rect 4721 16133 4755 16167
rect 5457 16133 5491 16167
rect 9597 16133 9631 16167
rect 9689 16133 9723 16167
rect 13185 16133 13219 16167
rect 13277 16133 13311 16167
rect 17141 16133 17175 16167
rect 20361 16133 20395 16167
rect 22845 16133 22879 16167
rect 22937 16133 22971 16167
rect 24501 16133 24535 16167
rect 26065 16133 26099 16167
rect 26617 16133 26651 16167
rect 1593 16065 1627 16099
rect 2881 16065 2915 16099
rect 3525 16065 3559 16099
rect 3985 16065 4019 16099
rect 4629 16065 4663 16099
rect 6929 16065 6963 16099
rect 7573 16065 7607 16099
rect 8217 16065 8251 16099
rect 8861 16065 8895 16099
rect 12173 16065 12207 16099
rect 15209 16065 15243 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 17969 16065 18003 16099
rect 19073 16065 19107 16099
rect 22017 16065 22051 16099
rect 38301 16065 38335 16099
rect 5365 15997 5399 16031
rect 6009 15997 6043 16031
rect 10609 15997 10643 16031
rect 12357 15997 12391 16031
rect 14197 15997 14231 16031
rect 15025 15997 15059 16031
rect 20269 15997 20303 16031
rect 20913 15997 20947 16031
rect 23121 15997 23155 16031
rect 24409 15997 24443 16031
rect 25421 15997 25455 16031
rect 25973 15997 26007 16031
rect 4077 15929 4111 15963
rect 7665 15929 7699 15963
rect 15393 15929 15427 15963
rect 22109 15929 22143 15963
rect 1777 15861 1811 15895
rect 3341 15861 3375 15895
rect 7021 15861 7055 15895
rect 8953 15861 8987 15895
rect 18061 15861 18095 15895
rect 19165 15861 19199 15895
rect 38117 15861 38151 15895
rect 1961 15657 1995 15691
rect 16773 15657 16807 15691
rect 20821 15657 20855 15691
rect 21649 15657 21683 15691
rect 29101 15657 29135 15691
rect 18337 15589 18371 15623
rect 6469 15521 6503 15555
rect 12081 15521 12115 15555
rect 13093 15521 13127 15555
rect 14933 15521 14967 15555
rect 15393 15521 15427 15555
rect 16405 15521 16439 15555
rect 16589 15521 16623 15555
rect 17785 15521 17819 15555
rect 19625 15521 19659 15555
rect 22753 15521 22787 15555
rect 29837 15521 29871 15555
rect 30113 15521 30147 15555
rect 37749 15521 37783 15555
rect 2145 15453 2179 15487
rect 3249 15453 3283 15487
rect 4261 15453 4295 15487
rect 6285 15453 6319 15487
rect 7757 15453 7791 15487
rect 8401 15453 8435 15487
rect 11069 15453 11103 15487
rect 13553 15453 13587 15487
rect 20269 15453 20303 15487
rect 20729 15453 20763 15487
rect 21557 15453 21591 15487
rect 23397 15453 23431 15487
rect 23857 15453 23891 15487
rect 24593 15453 24627 15487
rect 25237 15453 25271 15487
rect 29009 15453 29043 15487
rect 37473 15453 37507 15487
rect 2605 15385 2639 15419
rect 4997 15385 5031 15419
rect 5089 15385 5123 15419
rect 5641 15385 5675 15419
rect 7849 15385 7883 15419
rect 9781 15385 9815 15419
rect 9873 15385 9907 15419
rect 10425 15385 10459 15419
rect 11345 15385 11379 15419
rect 12173 15385 12207 15419
rect 15025 15385 15059 15419
rect 17877 15385 17911 15419
rect 19717 15385 19751 15419
rect 22845 15385 22879 15419
rect 24685 15385 24719 15419
rect 29929 15385 29963 15419
rect 3341 15317 3375 15351
rect 4353 15317 4387 15351
rect 6929 15317 6963 15351
rect 8493 15317 8527 15351
rect 13645 15317 13679 15351
rect 23949 15317 23983 15351
rect 25329 15317 25363 15351
rect 2053 15113 2087 15147
rect 9597 15113 9631 15147
rect 27537 15113 27571 15147
rect 28089 15113 28123 15147
rect 10333 15045 10367 15079
rect 12541 15045 12575 15079
rect 13369 15045 13403 15079
rect 13921 15045 13955 15079
rect 15301 15045 15335 15079
rect 17417 15045 17451 15079
rect 18613 15045 18647 15079
rect 21005 15045 21039 15079
rect 22201 15045 22235 15079
rect 23673 15045 23707 15079
rect 23765 15045 23799 15079
rect 1961 14977 1995 15011
rect 2605 14977 2639 15011
rect 3249 14977 3283 15011
rect 3893 14977 3927 15011
rect 4537 14977 4571 15011
rect 5181 14977 5215 15011
rect 5825 14977 5859 15011
rect 6929 14977 6963 15011
rect 7573 14977 7607 15011
rect 8217 14977 8251 15011
rect 8861 14977 8895 15011
rect 9505 14977 9539 15011
rect 12265 14977 12299 15011
rect 14381 14977 14415 15011
rect 19625 14977 19659 15011
rect 20269 14977 20303 15011
rect 20913 14977 20947 15011
rect 26249 14977 26283 15011
rect 27445 14977 27479 15011
rect 28273 14977 28307 15011
rect 28917 14977 28951 15011
rect 38025 14977 38059 15011
rect 10241 14909 10275 14943
rect 13277 14909 13311 14943
rect 15209 14909 15243 14943
rect 16221 14909 16255 14943
rect 17325 14909 17359 14943
rect 17601 14909 17635 14943
rect 18521 14909 18555 14943
rect 19165 14909 19199 14943
rect 22109 14909 22143 14943
rect 23121 14909 23155 14943
rect 23949 14909 23983 14943
rect 30113 14909 30147 14943
rect 3985 14841 4019 14875
rect 8953 14841 8987 14875
rect 10793 14841 10827 14875
rect 20361 14841 20395 14875
rect 2697 14773 2731 14807
rect 3341 14773 3375 14807
rect 4629 14773 4663 14807
rect 5273 14773 5307 14807
rect 5917 14773 5951 14807
rect 7021 14773 7055 14807
rect 7665 14773 7699 14807
rect 8309 14773 8343 14807
rect 14565 14773 14599 14807
rect 19717 14773 19751 14807
rect 26065 14773 26099 14807
rect 28733 14773 28767 14807
rect 37841 14773 37875 14807
rect 9505 14569 9539 14603
rect 21649 14569 21683 14603
rect 26249 14569 26283 14603
rect 30389 14501 30423 14535
rect 2789 14433 2823 14467
rect 4445 14433 4479 14467
rect 7205 14433 7239 14467
rect 10793 14433 10827 14467
rect 12725 14433 12759 14467
rect 17785 14433 17819 14467
rect 18705 14433 18739 14467
rect 20545 14433 20579 14467
rect 23489 14433 23523 14467
rect 30021 14433 30055 14467
rect 30205 14433 30239 14467
rect 1593 14365 1627 14399
rect 6469 14365 6503 14399
rect 7113 14365 7147 14399
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 9413 14365 9447 14399
rect 10057 14365 10091 14399
rect 14289 14365 14323 14399
rect 17509 14365 17543 14399
rect 18429 14365 18463 14399
rect 21557 14365 21591 14399
rect 24593 14365 24627 14399
rect 25237 14365 25271 14399
rect 26157 14365 26191 14399
rect 27261 14365 27295 14399
rect 27721 14365 27755 14399
rect 28365 14365 28399 14399
rect 2881 14297 2915 14331
rect 3433 14297 3467 14331
rect 4537 14297 4571 14331
rect 5457 14297 5491 14331
rect 6561 14297 6595 14331
rect 10885 14297 10919 14331
rect 11805 14297 11839 14331
rect 12817 14297 12851 14331
rect 13737 14297 13771 14331
rect 15025 14297 15059 14331
rect 15669 14297 15703 14331
rect 16405 14297 16439 14331
rect 19533 14297 19567 14331
rect 19625 14297 19659 14331
rect 22845 14297 22879 14331
rect 22937 14297 22971 14331
rect 27813 14297 27847 14331
rect 1777 14229 1811 14263
rect 7849 14229 7883 14263
rect 8493 14229 8527 14263
rect 10149 14229 10183 14263
rect 24685 14229 24719 14263
rect 25329 14229 25363 14263
rect 27077 14229 27111 14263
rect 28457 14229 28491 14263
rect 5917 14025 5951 14059
rect 6653 14025 6687 14059
rect 24869 14025 24903 14059
rect 25513 14025 25547 14059
rect 3341 13957 3375 13991
rect 4629 13957 4663 13991
rect 7297 13957 7331 13991
rect 10241 13957 10275 13991
rect 12541 13957 12575 13991
rect 12633 13957 12667 13991
rect 14197 13957 14231 13991
rect 15761 13957 15795 13991
rect 16313 13957 16347 13991
rect 17049 13957 17083 13991
rect 17601 13957 17635 13991
rect 18981 13957 19015 13991
rect 19901 13957 19935 13991
rect 20545 13957 20579 13991
rect 23397 13957 23431 13991
rect 27353 13957 27387 13991
rect 29469 13957 29503 13991
rect 1593 13889 1627 13923
rect 2513 13889 2547 13923
rect 4537 13889 4571 13923
rect 5181 13889 5215 13923
rect 5825 13889 5859 13923
rect 6561 13889 6595 13923
rect 7205 13889 7239 13923
rect 7849 13889 7883 13923
rect 8493 13889 8527 13923
rect 9781 13889 9815 13923
rect 11805 13889 11839 13923
rect 11897 13889 11931 13923
rect 18153 13889 18187 13923
rect 22017 13889 22051 13923
rect 24777 13889 24811 13923
rect 25421 13889 25455 13923
rect 27905 13889 27939 13923
rect 37749 13889 37783 13923
rect 3249 13821 3283 13855
rect 3525 13821 3559 13855
rect 5273 13821 5307 13855
rect 8585 13821 8619 13855
rect 9137 13821 9171 13855
rect 9321 13821 9355 13855
rect 11069 13821 11103 13855
rect 13553 13821 13587 13855
rect 14105 13821 14139 13855
rect 15117 13821 15151 13855
rect 15669 13821 15703 13855
rect 16957 13821 16991 13855
rect 18245 13821 18279 13855
rect 18889 13821 18923 13855
rect 20453 13821 20487 13855
rect 21373 13821 21407 13855
rect 23305 13821 23339 13855
rect 24317 13821 24351 13855
rect 27261 13821 27295 13855
rect 29377 13821 29411 13855
rect 29653 13821 29687 13855
rect 37473 13821 37507 13855
rect 1777 13685 1811 13719
rect 2605 13685 2639 13719
rect 7941 13685 7975 13719
rect 22109 13685 22143 13719
rect 13001 13481 13035 13515
rect 2881 13345 2915 13379
rect 4629 13345 4663 13379
rect 7297 13345 7331 13379
rect 9781 13345 9815 13379
rect 10057 13345 10091 13379
rect 13645 13345 13679 13379
rect 18797 13345 18831 13379
rect 28365 13345 28399 13379
rect 4537 13277 4571 13311
rect 5365 13277 5399 13311
rect 6009 13277 6043 13311
rect 6101 13277 6135 13311
rect 8401 13277 8435 13311
rect 11253 13277 11287 13311
rect 13553 13277 13587 13311
rect 21189 13277 21223 13311
rect 21833 13277 21867 13311
rect 22477 13277 22511 13311
rect 23121 13277 23155 13311
rect 23765 13277 23799 13311
rect 1869 13209 1903 13243
rect 1961 13209 1995 13243
rect 6745 13209 6779 13243
rect 6837 13209 6871 13243
rect 9873 13209 9907 13243
rect 11529 13209 11563 13243
rect 14381 13209 14415 13243
rect 14473 13209 14507 13243
rect 15393 13209 15427 13243
rect 16221 13209 16255 13243
rect 16313 13209 16347 13243
rect 17233 13209 17267 13243
rect 17785 13209 17819 13243
rect 17877 13209 17911 13243
rect 19717 13209 19751 13243
rect 19809 13209 19843 13243
rect 20729 13209 20763 13243
rect 23213 13209 23247 13243
rect 24685 13209 24719 13243
rect 24777 13209 24811 13243
rect 25697 13209 25731 13243
rect 26249 13209 26283 13243
rect 26341 13209 26375 13243
rect 27261 13209 27295 13243
rect 28089 13209 28123 13243
rect 28181 13209 28215 13243
rect 5457 13141 5491 13175
rect 8493 13141 8527 13175
rect 21281 13141 21315 13175
rect 21925 13141 21959 13175
rect 22569 13141 22603 13175
rect 23857 13141 23891 13175
rect 23581 12937 23615 12971
rect 29469 12937 29503 12971
rect 6837 12869 6871 12903
rect 7389 12869 7423 12903
rect 8033 12869 8067 12903
rect 14841 12869 14875 12903
rect 21189 12869 21223 12903
rect 22385 12869 22419 12903
rect 22477 12869 22511 12903
rect 24869 12869 24903 12903
rect 27445 12869 27479 12903
rect 28365 12869 28399 12903
rect 1593 12801 1627 12835
rect 2789 12801 2823 12835
rect 3433 12801 3467 12835
rect 4077 12801 4111 12835
rect 4721 12801 4755 12835
rect 5365 12801 5399 12835
rect 11713 12801 11747 12835
rect 12357 12801 12391 12835
rect 14565 12801 14599 12835
rect 16865 12801 16899 12835
rect 20453 12801 20487 12835
rect 21097 12801 21131 12835
rect 23489 12801 23523 12835
rect 24133 12801 24167 12835
rect 24777 12801 24811 12835
rect 38025 12801 38059 12835
rect 6745 12733 6779 12767
rect 7941 12733 7975 12767
rect 8953 12733 8987 12767
rect 9413 12733 9447 12767
rect 9689 12733 9723 12767
rect 12633 12733 12667 12767
rect 16313 12733 16347 12767
rect 17049 12733 17083 12767
rect 17969 12733 18003 12767
rect 18245 12733 18279 12767
rect 19717 12733 19751 12767
rect 27353 12733 27387 12767
rect 28825 12733 28859 12767
rect 29009 12733 29043 12767
rect 4169 12665 4203 12699
rect 5457 12665 5491 12699
rect 11161 12665 11195 12699
rect 22937 12665 22971 12699
rect 1777 12597 1811 12631
rect 2881 12597 2915 12631
rect 3525 12597 3559 12631
rect 4813 12597 4847 12631
rect 11805 12597 11839 12631
rect 14105 12597 14139 12631
rect 20545 12597 20579 12631
rect 24225 12597 24259 12631
rect 38209 12597 38243 12631
rect 2421 12393 2455 12427
rect 15926 12393 15960 12427
rect 27077 12393 27111 12427
rect 28365 12393 28399 12427
rect 17417 12325 17451 12359
rect 4629 12257 4663 12291
rect 5457 12257 5491 12291
rect 9505 12257 9539 12291
rect 13737 12257 13771 12291
rect 15669 12257 15703 12291
rect 22293 12257 22327 12291
rect 27629 12257 27663 12291
rect 30849 12257 30883 12291
rect 2329 12189 2363 12223
rect 6101 12189 6135 12223
rect 8401 12189 8435 12223
rect 11989 12189 12023 12223
rect 14749 12189 14783 12223
rect 18429 12189 18463 12223
rect 19533 12189 19567 12223
rect 22937 12189 22971 12223
rect 23397 12189 23431 12223
rect 24593 12189 24627 12223
rect 26157 12189 26191 12223
rect 26985 12189 27019 12223
rect 28273 12189 28307 12223
rect 4721 12121 4755 12155
rect 6377 12121 6411 12155
rect 9781 12121 9815 12155
rect 12265 12121 12299 12155
rect 15025 12121 15059 12155
rect 18521 12121 18555 12155
rect 19809 12121 19843 12155
rect 22385 12121 22419 12155
rect 24685 12121 24719 12155
rect 29837 12121 29871 12155
rect 29929 12121 29963 12155
rect 7849 12053 7883 12087
rect 8493 12053 8527 12087
rect 11253 12053 11287 12087
rect 21281 12053 21315 12087
rect 23489 12053 23523 12087
rect 26249 12053 26283 12087
rect 1593 11849 1627 11883
rect 3249 11849 3283 11883
rect 4629 11849 4663 11883
rect 16313 11849 16347 11883
rect 25789 11849 25823 11883
rect 35725 11849 35759 11883
rect 5273 11781 5307 11815
rect 10241 11781 10275 11815
rect 18521 11781 18555 11815
rect 20913 11781 20947 11815
rect 22293 11781 22327 11815
rect 23029 11781 23063 11815
rect 27261 11781 27295 11815
rect 27353 11781 27387 11815
rect 1777 11713 1811 11747
rect 3433 11713 3467 11747
rect 4077 11713 4111 11747
rect 4537 11713 4571 11747
rect 5181 11713 5215 11747
rect 5825 11713 5859 11747
rect 6745 11713 6779 11747
rect 7389 11713 7423 11747
rect 12081 11713 12115 11747
rect 14565 11713 14599 11747
rect 16865 11713 16899 11747
rect 18245 11713 18279 11747
rect 22201 11713 22235 11747
rect 24409 11713 24443 11747
rect 25053 11713 25087 11747
rect 25697 11713 25731 11747
rect 35909 11713 35943 11747
rect 7665 11645 7699 11679
rect 10149 11645 10183 11679
rect 11161 11645 11195 11679
rect 12357 11645 12391 11679
rect 14105 11645 14139 11679
rect 14841 11645 14875 11679
rect 17049 11645 17083 11679
rect 20269 11645 20303 11679
rect 20821 11645 20855 11679
rect 21097 11645 21131 11679
rect 22937 11645 22971 11679
rect 23949 11645 23983 11679
rect 27537 11645 27571 11679
rect 3893 11577 3927 11611
rect 5917 11577 5951 11611
rect 25145 11577 25179 11611
rect 6837 11509 6871 11543
rect 9137 11509 9171 11543
rect 24501 11509 24535 11543
rect 4261 11305 4295 11339
rect 8585 11305 8619 11339
rect 9413 11305 9447 11339
rect 13461 11305 13495 11339
rect 16852 11305 16886 11339
rect 18337 11305 18371 11339
rect 19980 11305 20014 11339
rect 21465 11305 21499 11339
rect 26893 11305 26927 11339
rect 33241 11305 33275 11339
rect 10057 11237 10091 11271
rect 1869 11169 1903 11203
rect 10609 11169 10643 11203
rect 12633 11169 12667 11203
rect 14289 11169 14323 11203
rect 14565 11169 14599 11203
rect 16037 11169 16071 11203
rect 16589 11169 16623 11203
rect 19717 11169 19751 11203
rect 1593 11101 1627 11135
rect 4169 11101 4203 11135
rect 4813 11101 4847 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 9321 11101 9355 11135
rect 9965 11101 9999 11135
rect 13369 11101 13403 11135
rect 22017 11101 22051 11135
rect 24593 11101 24627 11135
rect 25237 11101 25271 11135
rect 26801 11101 26835 11135
rect 33149 11101 33183 11135
rect 38301 11101 38335 11135
rect 4905 11033 4939 11067
rect 5457 11033 5491 11067
rect 7113 11033 7147 11067
rect 10885 11033 10919 11067
rect 22293 11033 22327 11067
rect 25329 11033 25363 11067
rect 2881 10965 2915 10999
rect 23765 10965 23799 10999
rect 24685 10965 24719 10999
rect 38117 10965 38151 10999
rect 4261 10761 4295 10795
rect 5273 10761 5307 10795
rect 6653 10761 6687 10795
rect 12725 10761 12759 10795
rect 15025 10761 15059 10795
rect 16221 10761 16255 10795
rect 18613 10761 18647 10795
rect 17141 10693 17175 10727
rect 27261 10693 27295 10727
rect 27997 10693 28031 10727
rect 1593 10625 1627 10659
rect 2697 10625 2731 10659
rect 4169 10625 4203 10659
rect 5181 10625 5215 10659
rect 5825 10625 5859 10659
rect 6561 10625 6595 10659
rect 7197 10625 7231 10659
rect 7856 10625 7890 10659
rect 10149 10625 10183 10659
rect 10793 10625 10827 10659
rect 11805 10625 11839 10659
rect 12633 10625 12667 10659
rect 16129 10625 16163 10659
rect 22017 10625 22051 10659
rect 27169 10625 27203 10659
rect 38025 10625 38059 10659
rect 1777 10557 1811 10591
rect 2881 10557 2915 10591
rect 8125 10557 8159 10591
rect 13277 10557 13311 10591
rect 13553 10557 13587 10591
rect 16865 10557 16899 10591
rect 19257 10557 19291 10591
rect 19533 10557 19567 10591
rect 21281 10557 21315 10591
rect 22293 10557 22327 10591
rect 23765 10557 23799 10591
rect 27905 10557 27939 10591
rect 10241 10489 10275 10523
rect 28457 10489 28491 10523
rect 2237 10421 2271 10455
rect 3065 10421 3099 10455
rect 5917 10421 5951 10455
rect 7297 10421 7331 10455
rect 9597 10421 9631 10455
rect 10885 10421 10919 10455
rect 11897 10421 11931 10455
rect 38209 10421 38243 10455
rect 1961 10217 1995 10251
rect 2513 10217 2547 10251
rect 3157 10217 3191 10251
rect 6285 10217 6319 10251
rect 8585 10217 8619 10251
rect 37841 10217 37875 10251
rect 11437 10149 11471 10183
rect 17693 10149 17727 10183
rect 18245 10149 18279 10183
rect 21373 10149 21407 10183
rect 30389 10149 30423 10183
rect 5641 10081 5675 10115
rect 9965 10081 9999 10115
rect 11897 10081 11931 10115
rect 15025 10081 15059 10115
rect 15945 10081 15979 10115
rect 19901 10081 19935 10115
rect 23305 10081 23339 10115
rect 1869 10013 1903 10047
rect 2697 10013 2731 10047
rect 3341 10013 3375 10047
rect 4169 10013 4203 10047
rect 5549 10013 5583 10047
rect 6193 10013 6227 10047
rect 6837 10013 6871 10047
rect 9689 10013 9723 10047
rect 18153 10013 18187 10047
rect 19625 10013 19659 10047
rect 22569 10013 22603 10047
rect 24593 10013 24627 10047
rect 25237 10013 25271 10047
rect 38025 10013 38059 10047
rect 7113 9945 7147 9979
rect 12173 9945 12207 9979
rect 14289 9945 14323 9979
rect 16221 9945 16255 9979
rect 21833 9945 21867 9979
rect 23397 9945 23431 9979
rect 23949 9945 23983 9979
rect 29837 9945 29871 9979
rect 29929 9945 29963 9979
rect 3985 9877 4019 9911
rect 13645 9877 13679 9911
rect 24685 9877 24719 9911
rect 25329 9877 25363 9911
rect 27445 9877 27479 9911
rect 1869 9673 1903 9707
rect 29929 9673 29963 9707
rect 13461 9605 13495 9639
rect 16221 9605 16255 9639
rect 19901 9605 19935 9639
rect 24133 9605 24167 9639
rect 24777 9605 24811 9639
rect 24869 9605 24903 9639
rect 27445 9605 27479 9639
rect 27537 9605 27571 9639
rect 2053 9537 2087 9571
rect 2513 9537 2547 9571
rect 3157 9537 3191 9571
rect 7205 9537 7239 9571
rect 11713 9537 11747 9571
rect 12541 9537 12575 9571
rect 13185 9537 13219 9571
rect 15485 9537 15519 9571
rect 16129 9537 16163 9571
rect 22477 9537 22511 9571
rect 23121 9537 23155 9571
rect 24041 9537 24075 9571
rect 25881 9537 25915 9571
rect 28917 9537 28951 9571
rect 29837 9537 29871 9571
rect 2605 9469 2639 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 7481 9469 7515 9503
rect 9413 9469 9447 9503
rect 9689 9469 9723 9503
rect 15577 9469 15611 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 19625 9469 19659 9503
rect 21373 9469 21407 9503
rect 27997 9469 28031 9503
rect 6009 9401 6043 9435
rect 8953 9401 8987 9435
rect 23213 9401 23247 9435
rect 25329 9401 25363 9435
rect 3249 9333 3283 9367
rect 11161 9333 11195 9367
rect 12633 9333 12667 9367
rect 14933 9333 14967 9367
rect 18613 9333 18647 9367
rect 22569 9333 22603 9367
rect 25973 9333 26007 9367
rect 29009 9333 29043 9367
rect 2697 9129 2731 9163
rect 4997 9129 5031 9163
rect 11437 9129 11471 9163
rect 14381 9129 14415 9163
rect 16865 9129 16899 9163
rect 18521 9129 18555 9163
rect 13645 9061 13679 9095
rect 24041 9061 24075 9095
rect 11897 8993 11931 9027
rect 15117 8993 15151 9027
rect 19809 8993 19843 9027
rect 20085 8993 20119 9027
rect 22293 8993 22327 9027
rect 22569 8993 22603 9027
rect 26525 8993 26559 9027
rect 2053 8925 2087 8959
rect 2881 8925 2915 8959
rect 3985 8925 4019 8959
rect 4905 8925 4939 8959
rect 5733 8925 5767 8959
rect 6745 8925 6779 8959
rect 9696 8925 9730 8959
rect 14289 8925 14323 8959
rect 18429 8925 18463 8959
rect 24593 8925 24627 8959
rect 25237 8925 25271 8959
rect 34897 8925 34931 8959
rect 38025 8925 38059 8959
rect 7021 8857 7055 8891
rect 9965 8857 9999 8891
rect 12173 8857 12207 8891
rect 15393 8857 15427 8891
rect 21833 8857 21867 8891
rect 25329 8857 25363 8891
rect 26157 8857 26191 8891
rect 26249 8857 26283 8891
rect 2145 8789 2179 8823
rect 4077 8789 4111 8823
rect 5549 8789 5583 8823
rect 8493 8789 8527 8823
rect 24685 8789 24719 8823
rect 34989 8789 35023 8823
rect 38209 8789 38243 8823
rect 6009 8585 6043 8619
rect 28365 8585 28399 8619
rect 29653 8585 29687 8619
rect 36093 8585 36127 8619
rect 2145 8517 2179 8551
rect 12449 8517 12483 8551
rect 13461 8517 13495 8551
rect 23673 8517 23707 8551
rect 25237 8517 25271 8551
rect 26157 8517 26191 8551
rect 2329 8449 2363 8483
rect 2973 8449 3007 8483
rect 3433 8449 3467 8483
rect 7205 8449 7239 8483
rect 9413 8449 9447 8483
rect 11161 8449 11195 8483
rect 11713 8449 11747 8483
rect 13185 8449 13219 8483
rect 17233 8449 17267 8483
rect 19533 8449 19567 8483
rect 28273 8449 28307 8483
rect 28917 8449 28951 8483
rect 29561 8449 29595 8483
rect 36277 8449 36311 8483
rect 3525 8381 3559 8415
rect 4261 8381 4295 8415
rect 4537 8381 4571 8415
rect 7481 8381 7515 8415
rect 17509 8381 17543 8415
rect 21281 8381 21315 8415
rect 23581 8381 23615 8415
rect 24041 8381 24075 8415
rect 25145 8381 25179 8415
rect 27169 8381 27203 8415
rect 27353 8381 27387 8415
rect 29009 8381 29043 8415
rect 2789 8313 2823 8347
rect 27813 8313 27847 8347
rect 8953 8245 8987 8279
rect 14933 8245 14967 8279
rect 18981 8245 19015 8279
rect 19790 8245 19824 8279
rect 2513 8041 2547 8075
rect 4077 8041 4111 8075
rect 4892 8041 4926 8075
rect 6377 8041 6411 8075
rect 12725 7973 12759 8007
rect 17969 7973 18003 8007
rect 4629 7905 4663 7939
rect 6837 7905 6871 7939
rect 7113 7905 7147 7939
rect 10977 7905 11011 7939
rect 16221 7905 16255 7939
rect 16497 7905 16531 7939
rect 19533 7905 19567 7939
rect 19809 7905 19843 7939
rect 21557 7905 21591 7939
rect 27537 7905 27571 7939
rect 28549 7905 28583 7939
rect 29193 7905 29227 7939
rect 2053 7837 2087 7871
rect 2697 7837 2731 7871
rect 3341 7837 3375 7871
rect 3985 7837 4019 7871
rect 13277 7837 13311 7871
rect 18521 7837 18555 7871
rect 23397 7837 23431 7871
rect 38025 7837 38059 7871
rect 11253 7769 11287 7803
rect 13369 7769 13403 7803
rect 14749 7769 14783 7803
rect 15485 7769 15519 7803
rect 24685 7769 24719 7803
rect 24777 7769 24811 7803
rect 25697 7769 25731 7803
rect 26433 7769 26467 7803
rect 26525 7769 26559 7803
rect 27077 7769 27111 7803
rect 28641 7769 28675 7803
rect 1869 7701 1903 7735
rect 3157 7701 3191 7735
rect 8585 7701 8619 7735
rect 18613 7701 18647 7735
rect 23489 7701 23523 7735
rect 38209 7701 38243 7735
rect 2881 7497 2915 7531
rect 4537 7497 4571 7531
rect 21189 7497 21223 7531
rect 24961 7497 24995 7531
rect 27261 7497 27295 7531
rect 5825 7429 5859 7463
rect 6653 7429 6687 7463
rect 8033 7429 8067 7463
rect 10241 7429 10275 7463
rect 13277 7429 13311 7463
rect 23213 7429 23247 7463
rect 24225 7429 24259 7463
rect 1869 7361 1903 7395
rect 3065 7361 3099 7395
rect 3801 7361 3835 7395
rect 4445 7361 4479 7395
rect 5089 7361 5123 7395
rect 6561 7361 6595 7395
rect 11989 7361 12023 7395
rect 15025 7361 15059 7395
rect 24869 7361 24903 7395
rect 25513 7361 25547 7395
rect 26157 7361 26191 7395
rect 27169 7361 27203 7395
rect 38301 7361 38335 7395
rect 1593 7293 1627 7327
rect 7757 7293 7791 7327
rect 9781 7293 9815 7327
rect 10977 7293 11011 7327
rect 11713 7293 11747 7327
rect 13001 7293 13035 7327
rect 16865 7293 16899 7327
rect 17141 7293 17175 7327
rect 19441 7293 19475 7327
rect 23121 7293 23155 7327
rect 25605 7293 25639 7327
rect 23673 7225 23707 7259
rect 3893 7157 3927 7191
rect 18613 7157 18647 7191
rect 19704 7157 19738 7191
rect 26249 7157 26283 7191
rect 38117 7157 38151 7191
rect 4892 6953 4926 6987
rect 15380 6953 15414 6987
rect 19980 6953 20014 6987
rect 29009 6953 29043 6987
rect 2237 6885 2271 6919
rect 16865 6885 16899 6919
rect 29745 6885 29779 6919
rect 4629 6817 4663 6851
rect 6837 6817 6871 6851
rect 7113 6817 7147 6851
rect 9321 6817 9355 6851
rect 10241 6817 10275 6851
rect 10517 6817 10551 6851
rect 11989 6817 12023 6851
rect 18797 6817 18831 6851
rect 19717 6817 19751 6851
rect 21925 6817 21959 6851
rect 27813 6817 27847 6851
rect 27997 6817 28031 6851
rect 1777 6749 1811 6783
rect 2421 6749 2455 6783
rect 3065 6749 3099 6783
rect 4169 6749 4203 6783
rect 9229 6749 9263 6783
rect 13277 6749 13311 6783
rect 15117 6749 15151 6783
rect 17971 6749 18005 6783
rect 26525 6749 26559 6783
rect 27169 6749 27203 6783
rect 28457 6749 28491 6783
rect 29193 6749 29227 6783
rect 29929 6749 29963 6783
rect 33241 6749 33275 6783
rect 12541 6681 12575 6715
rect 22201 6681 22235 6715
rect 25053 6681 25087 6715
rect 25145 6681 25179 6715
rect 26065 6681 26099 6715
rect 27261 6681 27295 6715
rect 1593 6613 1627 6647
rect 2881 6613 2915 6647
rect 3985 6613 4019 6647
rect 6377 6613 6411 6647
rect 8585 6613 8619 6647
rect 21465 6613 21499 6647
rect 23673 6613 23707 6647
rect 26617 6613 26651 6647
rect 33333 6613 33367 6647
rect 6009 6409 6043 6443
rect 16129 6409 16163 6443
rect 27261 6409 27295 6443
rect 27905 6409 27939 6443
rect 29193 6409 29227 6443
rect 29837 6409 29871 6443
rect 4537 6341 4571 6375
rect 14289 6341 14323 6375
rect 23029 6341 23063 6375
rect 23121 6341 23155 6375
rect 28549 6341 28583 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 3249 6273 3283 6307
rect 3525 6273 3559 6307
rect 4261 6273 4295 6307
rect 6837 6273 6871 6307
rect 9413 6273 9447 6307
rect 12265 6273 12299 6307
rect 16313 6273 16347 6307
rect 16865 6273 16899 6307
rect 21465 6273 21499 6307
rect 22293 6273 22327 6307
rect 24501 6273 24535 6307
rect 25145 6273 25179 6307
rect 25789 6273 25823 6307
rect 25881 6273 25915 6307
rect 26433 6273 26467 6307
rect 27169 6273 27203 6307
rect 27813 6273 27847 6307
rect 28457 6273 28491 6307
rect 29101 6273 29135 6307
rect 29745 6273 29779 6307
rect 30573 6273 30607 6307
rect 7113 6205 7147 6239
rect 9689 6205 9723 6239
rect 12541 6205 12575 6239
rect 17141 6205 17175 6239
rect 19441 6205 19475 6239
rect 19717 6205 19751 6239
rect 24041 6205 24075 6239
rect 1777 6137 1811 6171
rect 8585 6137 8619 6171
rect 18613 6137 18647 6171
rect 2513 6069 2547 6103
rect 3709 6069 3743 6103
rect 11161 6069 11195 6103
rect 22385 6069 22419 6103
rect 24593 6069 24627 6103
rect 25237 6069 25271 6103
rect 26525 6069 26559 6103
rect 30389 6069 30423 6103
rect 27169 5865 27203 5899
rect 29101 5865 29135 5899
rect 17693 5797 17727 5831
rect 18429 5797 18463 5831
rect 26525 5797 26559 5831
rect 29745 5797 29779 5831
rect 2881 5729 2915 5763
rect 4261 5729 4295 5763
rect 6653 5729 6687 5763
rect 9137 5729 9171 5763
rect 10885 5729 10919 5763
rect 11437 5729 11471 5763
rect 16865 5729 16899 5763
rect 19809 5729 19843 5763
rect 24685 5729 24719 5763
rect 25881 5729 25915 5763
rect 1593 5661 1627 5695
rect 2605 5661 2639 5695
rect 3985 5661 4019 5695
rect 14657 5661 14691 5695
rect 15117 5661 15151 5695
rect 17509 5661 17543 5695
rect 18245 5661 18279 5695
rect 22017 5661 22051 5695
rect 23765 5661 23799 5695
rect 25329 5661 25363 5695
rect 25789 5661 25823 5695
rect 26433 5661 26467 5695
rect 27077 5661 27111 5695
rect 27721 5661 27755 5695
rect 27813 5661 27847 5695
rect 28365 5661 28399 5695
rect 29009 5661 29043 5695
rect 29929 5661 29963 5695
rect 30389 5661 30423 5695
rect 31033 5661 31067 5695
rect 31861 5661 31895 5695
rect 35541 5661 35575 5695
rect 38025 5661 38059 5695
rect 6929 5593 6963 5627
rect 9413 5593 9447 5627
rect 11713 5593 11747 5627
rect 13461 5593 13495 5627
rect 15393 5593 15427 5627
rect 20085 5593 20119 5627
rect 22753 5593 22787 5627
rect 24777 5593 24811 5627
rect 28457 5593 28491 5627
rect 30481 5593 30515 5627
rect 31125 5593 31159 5627
rect 1777 5525 1811 5559
rect 5733 5525 5767 5559
rect 8401 5525 8435 5559
rect 14473 5525 14507 5559
rect 21557 5525 21591 5559
rect 23857 5525 23891 5559
rect 31677 5525 31711 5559
rect 35357 5525 35391 5559
rect 38209 5525 38243 5559
rect 25973 5321 26007 5355
rect 29653 5321 29687 5355
rect 31585 5321 31619 5355
rect 7297 5253 7331 5287
rect 10425 5253 10459 5287
rect 12541 5253 12575 5287
rect 14749 5253 14783 5287
rect 19441 5253 19475 5287
rect 27261 5253 27295 5287
rect 27353 5253 27387 5287
rect 27905 5253 27939 5287
rect 28549 5253 28583 5287
rect 30297 5253 30331 5287
rect 1593 5185 1627 5219
rect 2881 5185 2915 5219
rect 4261 5185 4295 5219
rect 6561 5185 6595 5219
rect 8401 5185 8435 5219
rect 11161 5185 11195 5219
rect 12265 5185 12299 5219
rect 19165 5185 19199 5219
rect 22017 5185 22051 5219
rect 24593 5185 24627 5219
rect 25237 5185 25271 5219
rect 25881 5185 25915 5219
rect 29561 5185 29595 5219
rect 30205 5185 30239 5219
rect 30849 5185 30883 5219
rect 31493 5185 31527 5219
rect 32321 5185 32355 5219
rect 3709 5117 3743 5151
rect 4537 5117 4571 5151
rect 6009 5117 6043 5151
rect 8677 5117 8711 5151
rect 14473 5117 14507 5151
rect 16957 5117 16991 5151
rect 17233 5117 17267 5151
rect 20913 5117 20947 5151
rect 22293 5117 22327 5151
rect 28457 5117 28491 5151
rect 14013 5049 14047 5083
rect 18705 5049 18739 5083
rect 24685 5049 24719 5083
rect 29009 5049 29043 5083
rect 1777 4981 1811 5015
rect 10977 4981 11011 5015
rect 16221 4981 16255 5015
rect 23765 4981 23799 5015
rect 25329 4981 25363 5015
rect 30941 4981 30975 5015
rect 32413 4981 32447 5015
rect 7941 4777 7975 4811
rect 8401 4777 8435 4811
rect 11529 4777 11563 4811
rect 21189 4777 21223 4811
rect 28733 4777 28767 4811
rect 31769 4777 31803 4811
rect 3433 4709 3467 4743
rect 13737 4709 13771 4743
rect 27445 4709 27479 4743
rect 32321 4709 32355 4743
rect 33609 4709 33643 4743
rect 1961 4641 1995 4675
rect 3985 4641 4019 4675
rect 6193 4641 6227 4675
rect 9781 4641 9815 4675
rect 11989 4641 12023 4675
rect 15301 4641 15335 4675
rect 17049 4641 17083 4675
rect 18797 4641 18831 4675
rect 21649 4641 21683 4675
rect 29837 4641 29871 4675
rect 1685 4573 1719 4607
rect 8585 4573 8619 4607
rect 9137 4573 9171 4607
rect 14289 4573 14323 4607
rect 15025 4573 15059 4607
rect 17969 4573 18003 4607
rect 19441 4573 19475 4607
rect 25329 4573 25363 4607
rect 26065 4573 26099 4607
rect 26709 4573 26743 4607
rect 27353 4573 27387 4607
rect 27997 4573 28031 4607
rect 28641 4573 28675 4607
rect 29745 4573 29779 4607
rect 30389 4573 30423 4607
rect 31033 4573 31067 4607
rect 31677 4573 31711 4607
rect 32505 4573 32539 4607
rect 33149 4573 33183 4607
rect 33793 4573 33827 4607
rect 38025 4573 38059 4607
rect 4261 4505 4295 4539
rect 6469 4505 6503 4539
rect 10057 4505 10091 4539
rect 12265 4505 12299 4539
rect 19717 4505 19751 4539
rect 21925 4505 21959 4539
rect 24685 4505 24719 4539
rect 24777 4505 24811 4539
rect 31125 4505 31159 4539
rect 5733 4437 5767 4471
rect 9229 4437 9263 4471
rect 14473 4437 14507 4471
rect 23397 4437 23431 4471
rect 23857 4437 23891 4471
rect 26157 4437 26191 4471
rect 26801 4437 26835 4471
rect 28089 4437 28123 4471
rect 30481 4437 30515 4471
rect 32965 4437 32999 4471
rect 38209 4437 38243 4471
rect 33609 4233 33643 4267
rect 4537 4165 4571 4199
rect 14841 4165 14875 4199
rect 17141 4165 17175 4199
rect 19441 4165 19475 4199
rect 22477 4165 22511 4199
rect 24041 4165 24075 4199
rect 9413 4097 9447 4131
rect 11713 4097 11747 4131
rect 19165 4097 19199 4131
rect 24593 4097 24627 4131
rect 25053 4097 25087 4131
rect 25789 4097 25823 4131
rect 26433 4097 26467 4131
rect 27169 4097 27203 4131
rect 27813 4097 27847 4131
rect 28457 4097 28491 4131
rect 29101 4097 29135 4131
rect 29745 4097 29779 4131
rect 30389 4097 30423 4131
rect 30481 4097 30515 4131
rect 31033 4097 31067 4131
rect 32321 4097 32355 4131
rect 32965 4097 32999 4131
rect 33793 4097 33827 4131
rect 34253 4097 34287 4131
rect 38301 4097 38335 4131
rect 1685 4029 1719 4063
rect 1961 4029 1995 4063
rect 4261 4029 4295 4063
rect 6561 4029 6595 4063
rect 6837 4029 6871 4063
rect 9689 4029 9723 4063
rect 11989 4029 12023 4063
rect 13737 4029 13771 4063
rect 14565 4029 14599 4063
rect 16865 4029 16899 4063
rect 20913 4029 20947 4063
rect 22385 4029 22419 4063
rect 23397 4029 23431 4063
rect 23949 4029 23983 4063
rect 27905 4029 27939 4063
rect 25145 3961 25179 3995
rect 29193 3961 29227 3995
rect 32413 3961 32447 3995
rect 38117 3961 38151 3995
rect 3433 3893 3467 3927
rect 6009 3893 6043 3927
rect 8309 3893 8343 3927
rect 11161 3893 11195 3927
rect 16313 3893 16347 3927
rect 18613 3893 18647 3927
rect 25881 3893 25915 3927
rect 26525 3893 26559 3927
rect 27261 3893 27295 3927
rect 28549 3893 28583 3927
rect 29837 3893 29871 3927
rect 31125 3893 31159 3927
rect 33057 3893 33091 3927
rect 34345 3893 34379 3927
rect 3433 3689 3467 3723
rect 6377 3689 6411 3723
rect 29837 3689 29871 3723
rect 31769 3689 31803 3723
rect 36737 3689 36771 3723
rect 17601 3621 17635 3655
rect 21189 3621 21223 3655
rect 32321 3621 32355 3655
rect 1961 3553 1995 3587
rect 4629 3553 4663 3587
rect 6837 3553 6871 3587
rect 9781 3553 9815 3587
rect 10057 3553 10091 3587
rect 11989 3553 12023 3587
rect 15209 3553 15243 3587
rect 15853 3553 15887 3587
rect 18061 3553 18095 3587
rect 19441 3553 19475 3587
rect 22845 3553 22879 3587
rect 30481 3553 30515 3587
rect 1685 3485 1719 3519
rect 3985 3485 4019 3519
rect 9321 3485 9355 3519
rect 14473 3485 14507 3519
rect 18337 3485 18371 3519
rect 21741 3485 21775 3519
rect 26341 3485 26375 3519
rect 26801 3485 26835 3519
rect 27905 3485 27939 3519
rect 28181 3485 28215 3519
rect 28641 3485 28675 3519
rect 29745 3485 29779 3519
rect 30389 3485 30423 3519
rect 31033 3485 31067 3519
rect 31677 3485 31711 3519
rect 32505 3485 32539 3519
rect 32965 3485 32999 3519
rect 35081 3485 35115 3519
rect 35725 3485 35759 3519
rect 36921 3485 36955 3519
rect 38025 3485 38059 3519
rect 4905 3417 4939 3451
rect 7113 3417 7147 3451
rect 12265 3417 12299 3451
rect 16129 3417 16163 3451
rect 19717 3417 19751 3451
rect 22937 3417 22971 3451
rect 23489 3417 23523 3451
rect 24685 3417 24719 3451
rect 24777 3417 24811 3451
rect 25697 3417 25731 3451
rect 33057 3417 33091 3451
rect 4077 3349 4111 3383
rect 8585 3349 8619 3383
rect 9137 3349 9171 3383
rect 11529 3349 11563 3383
rect 13737 3349 13771 3383
rect 21925 3349 21959 3383
rect 26157 3349 26191 3383
rect 26893 3349 26927 3383
rect 28733 3349 28767 3383
rect 31125 3349 31159 3383
rect 33609 3349 33643 3383
rect 34897 3349 34931 3383
rect 35541 3349 35575 3383
rect 38209 3349 38243 3383
rect 6009 3145 6043 3179
rect 34345 3145 34379 3179
rect 35633 3145 35667 3179
rect 2329 3077 2363 3111
rect 8585 3077 8619 3111
rect 9689 3077 9723 3111
rect 12633 3077 12667 3111
rect 14841 3077 14875 3111
rect 22477 3077 22511 3111
rect 25605 3077 25639 3111
rect 25697 3077 25731 3111
rect 26617 3077 26651 3111
rect 27353 3077 27387 3111
rect 6561 3009 6595 3043
rect 9413 3009 9447 3043
rect 11713 3009 11747 3043
rect 14565 3009 14599 3043
rect 17141 3009 17175 3043
rect 19349 3009 19383 3043
rect 23857 3009 23891 3043
rect 24685 3009 24719 3043
rect 28549 3009 28583 3043
rect 29193 3009 29227 3043
rect 29653 3009 29687 3043
rect 30297 3009 30331 3043
rect 30941 3009 30975 3043
rect 31585 3009 31619 3043
rect 32321 3009 32355 3043
rect 32965 3009 32999 3043
rect 33609 3009 33643 3043
rect 34253 3009 34287 3043
rect 34897 3009 34931 3043
rect 35541 3009 35575 3043
rect 36369 3009 36403 3043
rect 38025 3009 38059 3043
rect 2053 2941 2087 2975
rect 4261 2941 4295 2975
rect 4537 2941 4571 2975
rect 6837 2941 6871 2975
rect 12357 2941 12391 2975
rect 16313 2941 16347 2975
rect 17417 2941 17451 2975
rect 19625 2941 19659 2975
rect 22385 2941 22419 2975
rect 22661 2941 22695 2975
rect 27261 2941 27295 2975
rect 29745 2941 29779 2975
rect 3801 2873 3835 2907
rect 11161 2873 11195 2907
rect 21097 2873 21131 2907
rect 23949 2873 23983 2907
rect 24501 2873 24535 2907
rect 27813 2873 27847 2907
rect 28365 2873 28399 2907
rect 29009 2873 29043 2907
rect 30389 2873 30423 2907
rect 31033 2873 31067 2907
rect 33701 2873 33735 2907
rect 11805 2805 11839 2839
rect 14105 2805 14139 2839
rect 18889 2805 18923 2839
rect 31677 2805 31711 2839
rect 32413 2805 32447 2839
rect 33057 2805 33091 2839
rect 34989 2805 35023 2839
rect 36185 2805 36219 2839
rect 38209 2805 38243 2839
rect 3433 2601 3467 2635
rect 13737 2601 13771 2635
rect 18889 2601 18923 2635
rect 21189 2601 21223 2635
rect 23857 2601 23891 2635
rect 27169 2601 27203 2635
rect 11161 2533 11195 2567
rect 25329 2533 25363 2567
rect 36093 2533 36127 2567
rect 1685 2465 1719 2499
rect 1961 2465 1995 2499
rect 4261 2465 4295 2499
rect 6837 2465 6871 2499
rect 9413 2465 9447 2499
rect 11989 2465 12023 2499
rect 14565 2465 14599 2499
rect 14841 2465 14875 2499
rect 17141 2465 17175 2499
rect 19441 2465 19475 2499
rect 19717 2465 19751 2499
rect 22385 2465 22419 2499
rect 22661 2465 22695 2499
rect 28089 2465 28123 2499
rect 30021 2465 30055 2499
rect 37749 2465 37783 2499
rect 24041 2397 24075 2431
rect 24777 2397 24811 2431
rect 25237 2397 25271 2431
rect 25881 2397 25915 2431
rect 27353 2397 27387 2431
rect 27813 2397 27847 2431
rect 29745 2397 29779 2431
rect 31033 2397 31067 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 35909 2397 35943 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 4537 2329 4571 2363
rect 7113 2329 7147 2363
rect 9689 2329 9723 2363
rect 12265 2329 12299 2363
rect 17417 2329 17451 2363
rect 22477 2329 22511 2363
rect 6009 2261 6043 2295
rect 8585 2261 8619 2295
rect 16313 2261 16347 2295
rect 24593 2261 24627 2295
rect 26065 2261 26099 2295
rect 31217 2261 31251 2295
rect 32505 2261 32539 2295
rect 33793 2261 33827 2295
rect 35081 2261 35115 2295
rect 36829 2261 36863 2295
<< metal1 >>
rect 16574 37612 16580 37664
rect 16632 37652 16638 37664
rect 19150 37652 19156 37664
rect 16632 37624 19156 37652
rect 16632 37612 16638 37624
rect 19150 37612 19156 37624
rect 19208 37612 19214 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 3145 37383 3203 37389
rect 3145 37349 3157 37383
rect 3191 37380 3203 37383
rect 16574 37380 16580 37392
rect 3191 37352 16580 37380
rect 3191 37349 3203 37352
rect 3145 37343 3203 37349
rect 16574 37340 16580 37352
rect 16632 37340 16638 37392
rect 17129 37383 17187 37389
rect 17129 37349 17141 37383
rect 17175 37380 17187 37383
rect 23566 37380 23572 37392
rect 17175 37352 23572 37380
rect 17175 37349 17187 37352
rect 17129 37343 17187 37349
rect 1578 37312 1584 37324
rect 1539 37284 1584 37312
rect 1578 37272 1584 37284
rect 1636 37272 1642 37324
rect 3878 37272 3884 37324
rect 3936 37312 3942 37324
rect 3973 37315 4031 37321
rect 3973 37312 3985 37315
rect 3936 37284 3985 37312
rect 3936 37272 3942 37284
rect 3973 37281 3985 37284
rect 4019 37281 4031 37315
rect 3973 37275 4031 37281
rect 5810 37272 5816 37324
rect 5868 37312 5874 37324
rect 6549 37315 6607 37321
rect 6549 37312 6561 37315
rect 5868 37284 6561 37312
rect 5868 37272 5874 37284
rect 6549 37281 6561 37284
rect 6595 37281 6607 37315
rect 6549 37275 6607 37281
rect 8386 37272 8392 37324
rect 8444 37312 8450 37324
rect 9125 37315 9183 37321
rect 9125 37312 9137 37315
rect 8444 37284 9137 37312
rect 8444 37272 8450 37284
rect 9125 37281 9137 37284
rect 9171 37281 9183 37315
rect 9125 37275 9183 37281
rect 16114 37272 16120 37324
rect 16172 37312 16178 37324
rect 17144 37312 17172 37343
rect 23566 37340 23572 37352
rect 23624 37340 23630 37392
rect 16172 37284 17172 37312
rect 16172 37272 16178 37284
rect 22554 37272 22560 37324
rect 22612 37312 22618 37324
rect 22649 37315 22707 37321
rect 22649 37312 22661 37315
rect 22612 37284 22661 37312
rect 22612 37272 22618 37284
rect 22649 37281 22661 37284
rect 22695 37281 22707 37315
rect 24854 37312 24860 37324
rect 24815 37284 24860 37312
rect 22649 37275 22707 37281
rect 24854 37272 24860 37284
rect 24912 37272 24918 37324
rect 27706 37272 27712 37324
rect 27764 37312 27770 37324
rect 27801 37315 27859 37321
rect 27801 37312 27813 37315
rect 27764 37284 27813 37312
rect 27764 37272 27770 37284
rect 27801 37281 27813 37284
rect 27847 37281 27859 37315
rect 27801 37275 27859 37281
rect 29638 37272 29644 37324
rect 29696 37312 29702 37324
rect 29696 37284 30236 37312
rect 29696 37272 29702 37284
rect 1854 37244 1860 37256
rect 1815 37216 1860 37244
rect 1854 37204 1860 37216
rect 1912 37204 1918 37256
rect 2774 37204 2780 37256
rect 2832 37244 2838 37256
rect 2961 37247 3019 37253
rect 2961 37244 2973 37247
rect 2832 37216 2973 37244
rect 2832 37204 2838 37216
rect 2961 37213 2973 37216
rect 3007 37213 3019 37247
rect 4246 37244 4252 37256
rect 4207 37216 4252 37244
rect 2961 37207 3019 37213
rect 4246 37204 4252 37216
rect 4304 37204 4310 37256
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5445 37247 5503 37253
rect 5445 37244 5457 37247
rect 5224 37216 5457 37244
rect 5224 37204 5230 37216
rect 5445 37213 5457 37216
rect 5491 37213 5503 37247
rect 6822 37244 6828 37256
rect 6783 37216 6828 37244
rect 5445 37207 5503 37213
rect 6822 37204 6828 37216
rect 6880 37204 6886 37256
rect 7098 37204 7104 37256
rect 7156 37244 7162 37256
rect 8021 37247 8079 37253
rect 8021 37244 8033 37247
rect 7156 37216 8033 37244
rect 7156 37204 7162 37216
rect 8021 37213 8033 37216
rect 8067 37213 8079 37247
rect 9398 37244 9404 37256
rect 9359 37216 9404 37244
rect 8021 37207 8079 37213
rect 9398 37204 9404 37216
rect 9456 37204 9462 37256
rect 10413 37247 10471 37253
rect 10413 37213 10425 37247
rect 10459 37244 10471 37247
rect 10459 37216 11468 37244
rect 10459 37213 10471 37216
rect 10413 37207 10471 37213
rect 11054 37176 11060 37188
rect 7852 37148 11060 37176
rect 5258 37108 5264 37120
rect 5219 37080 5264 37108
rect 5258 37068 5264 37080
rect 5316 37068 5322 37120
rect 7852 37117 7880 37148
rect 11054 37136 11060 37148
rect 11112 37136 11118 37188
rect 11440 37176 11468 37216
rect 11606 37204 11612 37256
rect 11664 37244 11670 37256
rect 11885 37247 11943 37253
rect 11885 37244 11897 37247
rect 11664 37216 11897 37244
rect 11664 37204 11670 37216
rect 11885 37213 11897 37216
rect 11931 37213 11943 37247
rect 11885 37207 11943 37213
rect 12434 37204 12440 37256
rect 12492 37244 12498 37256
rect 12529 37247 12587 37253
rect 12529 37244 12541 37247
rect 12492 37216 12541 37244
rect 12492 37204 12498 37216
rect 12529 37213 12541 37216
rect 12575 37213 12587 37247
rect 12529 37207 12587 37213
rect 13538 37204 13544 37256
rect 13596 37244 13602 37256
rect 14277 37247 14335 37253
rect 14277 37244 14289 37247
rect 13596 37216 14289 37244
rect 13596 37204 13602 37216
rect 14277 37213 14289 37216
rect 14323 37213 14335 37247
rect 14277 37207 14335 37213
rect 14645 37247 14703 37253
rect 14645 37213 14657 37247
rect 14691 37244 14703 37247
rect 14918 37244 14924 37256
rect 14691 37216 14924 37244
rect 14691 37213 14703 37216
rect 14645 37207 14703 37213
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18414 37204 18420 37256
rect 18472 37244 18478 37256
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 18472 37216 20085 37244
rect 18472 37204 18478 37216
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 20073 37207 20131 37213
rect 21266 37204 21272 37256
rect 21324 37244 21330 37256
rect 22189 37247 22247 37253
rect 22189 37244 22201 37247
rect 21324 37216 22201 37244
rect 21324 37204 21330 37216
rect 22189 37213 22201 37216
rect 22235 37213 22247 37247
rect 22189 37207 22247 37213
rect 22925 37247 22983 37253
rect 22925 37213 22937 37247
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 11440 37148 12572 37176
rect 12544 37120 12572 37148
rect 16574 37136 16580 37188
rect 16632 37176 16638 37188
rect 16945 37179 17003 37185
rect 16945 37176 16957 37179
rect 16632 37148 16957 37176
rect 16632 37136 16638 37148
rect 16945 37145 16957 37148
rect 16991 37145 17003 37179
rect 16945 37139 17003 37145
rect 21082 37136 21088 37188
rect 21140 37176 21146 37188
rect 22940 37176 22968 37207
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24673 37247 24731 37253
rect 24673 37244 24685 37247
rect 24544 37216 24685 37244
rect 24544 37204 24550 37216
rect 24673 37213 24685 37216
rect 24719 37213 24731 37247
rect 24673 37207 24731 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25832 37216 25881 37244
rect 25832 37204 25838 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 26326 37244 26332 37256
rect 26287 37216 26332 37244
rect 25869 37207 25927 37213
rect 26326 37204 26332 37216
rect 26384 37204 26390 37256
rect 28074 37244 28080 37256
rect 28035 37216 28080 37244
rect 28074 37204 28080 37216
rect 28132 37204 28138 37256
rect 28994 37204 29000 37256
rect 29052 37244 29058 37256
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29052 37216 29929 37244
rect 29052 37204 29058 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 30208 37244 30236 37284
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30208 37216 30573 37244
rect 29917 37207 29975 37213
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 31018 37244 31024 37256
rect 30979 37216 31024 37244
rect 30561 37207 30619 37213
rect 31018 37204 31024 37216
rect 31076 37204 31082 37256
rect 32122 37204 32128 37256
rect 32180 37244 32186 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 32180 37216 32321 37244
rect 32180 37204 32186 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 32309 37207 32367 37213
rect 32398 37204 32404 37256
rect 32456 37244 32462 37256
rect 33045 37247 33103 37253
rect 33045 37244 33057 37247
rect 32456 37216 33057 37244
rect 32456 37204 32462 37216
rect 33045 37213 33057 37216
rect 33091 37213 33103 37247
rect 34882 37244 34888 37256
rect 34843 37216 34888 37244
rect 33045 37207 33103 37213
rect 34882 37204 34888 37216
rect 34940 37204 34946 37256
rect 35526 37204 35532 37256
rect 35584 37244 35590 37256
rect 36173 37247 36231 37253
rect 36173 37244 36185 37247
rect 35584 37216 36185 37244
rect 35584 37204 35590 37216
rect 36173 37213 36185 37216
rect 36219 37213 36231 37247
rect 37458 37244 37464 37256
rect 37419 37216 37464 37244
rect 36173 37207 36231 37213
rect 37458 37204 37464 37216
rect 37516 37204 37522 37256
rect 21140 37148 22968 37176
rect 21140 37136 21146 37148
rect 7837 37111 7895 37117
rect 7837 37077 7849 37111
rect 7883 37077 7895 37111
rect 7837 37071 7895 37077
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10376 37080 10609 37108
rect 10376 37068 10382 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 11698 37108 11704 37120
rect 11659 37080 11704 37108
rect 10597 37071 10655 37077
rect 11698 37068 11704 37080
rect 11756 37068 11762 37120
rect 12342 37108 12348 37120
rect 12303 37080 12348 37108
rect 12342 37068 12348 37080
rect 12400 37068 12406 37120
rect 12526 37068 12532 37120
rect 12584 37068 12590 37120
rect 14090 37108 14096 37120
rect 14051 37080 14096 37108
rect 14090 37068 14096 37080
rect 14148 37068 14154 37120
rect 14826 37068 14832 37120
rect 14884 37108 14890 37120
rect 15105 37111 15163 37117
rect 15105 37108 15117 37111
rect 14884 37080 15117 37108
rect 14884 37068 14890 37080
rect 15105 37077 15117 37080
rect 15151 37077 15163 37111
rect 15105 37071 15163 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 18104 37080 18153 37108
rect 18104 37068 18110 37080
rect 18141 37077 18153 37080
rect 18187 37077 18199 37111
rect 18141 37071 18199 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 20346 37068 20352 37120
rect 20404 37108 20410 37120
rect 22005 37111 22063 37117
rect 22005 37108 22017 37111
rect 20404 37080 22017 37108
rect 20404 37068 20410 37080
rect 22005 37077 22017 37080
rect 22051 37077 22063 37111
rect 22005 37071 22063 37077
rect 23014 37068 23020 37120
rect 23072 37108 23078 37120
rect 25685 37111 25743 37117
rect 25685 37108 25697 37111
rect 23072 37080 25697 37108
rect 23072 37068 23078 37080
rect 25685 37077 25697 37080
rect 25731 37077 25743 37111
rect 25685 37071 25743 37077
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 26513 37111 26571 37117
rect 26513 37108 26525 37111
rect 26476 37080 26525 37108
rect 26476 37068 26482 37080
rect 26513 37077 26525 37080
rect 26559 37077 26571 37111
rect 26513 37071 26571 37077
rect 27154 37068 27160 37120
rect 27212 37108 27218 37120
rect 29733 37111 29791 37117
rect 29733 37108 29745 37111
rect 27212 37080 29745 37108
rect 27212 37068 27218 37080
rect 29733 37077 29745 37080
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 29822 37068 29828 37120
rect 29880 37108 29886 37120
rect 30377 37111 30435 37117
rect 30377 37108 30389 37111
rect 29880 37080 30389 37108
rect 29880 37068 29886 37080
rect 30377 37077 30389 37080
rect 30423 37077 30435 37111
rect 30377 37071 30435 37077
rect 30926 37068 30932 37120
rect 30984 37108 30990 37120
rect 31205 37111 31263 37117
rect 31205 37108 31217 37111
rect 30984 37080 31217 37108
rect 30984 37068 30990 37080
rect 31205 37077 31217 37080
rect 31251 37077 31263 37111
rect 31205 37071 31263 37077
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 32272 37080 32505 37108
rect 32272 37068 32278 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33134 37068 33140 37120
rect 33192 37108 33198 37120
rect 33229 37111 33287 37117
rect 33229 37108 33241 37111
rect 33192 37080 33241 37108
rect 33192 37068 33198 37080
rect 33229 37077 33241 37080
rect 33275 37077 33287 37111
rect 33229 37071 33287 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35069 37071 35127 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 36136 37080 36369 37108
rect 36136 37068 36142 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 36357 37071 36415 37077
rect 37366 37068 37372 37120
rect 37424 37108 37430 37120
rect 37645 37111 37703 37117
rect 37645 37108 37657 37111
rect 37424 37080 37657 37108
rect 37424 37068 37430 37080
rect 37645 37077 37657 37080
rect 37691 37077 37703 37111
rect 37645 37071 37703 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1762 36904 1768 36916
rect 1723 36876 1768 36904
rect 1762 36864 1768 36876
rect 1820 36864 1826 36916
rect 4246 36864 4252 36916
rect 4304 36904 4310 36916
rect 11790 36904 11796 36916
rect 4304 36876 11796 36904
rect 4304 36864 4310 36876
rect 11790 36864 11796 36876
rect 11848 36864 11854 36916
rect 17681 36907 17739 36913
rect 17681 36873 17693 36907
rect 17727 36904 17739 36907
rect 18414 36904 18420 36916
rect 17727 36876 18420 36904
rect 17727 36873 17739 36876
rect 17681 36867 17739 36873
rect 18414 36864 18420 36876
rect 18472 36864 18478 36916
rect 19334 36864 19340 36916
rect 19392 36904 19398 36916
rect 19613 36907 19671 36913
rect 19613 36904 19625 36907
rect 19392 36876 19625 36904
rect 19392 36864 19398 36876
rect 19613 36873 19625 36876
rect 19659 36873 19671 36907
rect 19613 36867 19671 36873
rect 29181 36907 29239 36913
rect 29181 36873 29193 36907
rect 29227 36904 29239 36907
rect 31018 36904 31024 36916
rect 29227 36876 31024 36904
rect 29227 36873 29239 36876
rect 29181 36867 29239 36873
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 31389 36907 31447 36913
rect 31389 36873 31401 36907
rect 31435 36904 31447 36907
rect 37458 36904 37464 36916
rect 31435 36876 37464 36904
rect 31435 36873 31447 36876
rect 31389 36867 31447 36873
rect 37458 36864 37464 36876
rect 37516 36864 37522 36916
rect 9398 36796 9404 36848
rect 9456 36836 9462 36848
rect 15562 36836 15568 36848
rect 9456 36808 15568 36836
rect 9456 36796 9462 36808
rect 15562 36796 15568 36808
rect 15620 36836 15626 36848
rect 15620 36808 17908 36836
rect 15620 36796 15626 36808
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36737 1639 36771
rect 1581 36731 1639 36737
rect 1596 36700 1624 36731
rect 1946 36728 1952 36780
rect 2004 36768 2010 36780
rect 2501 36771 2559 36777
rect 2501 36768 2513 36771
rect 2004 36740 2513 36768
rect 2004 36728 2010 36740
rect 2501 36737 2513 36740
rect 2547 36737 2559 36771
rect 3142 36768 3148 36780
rect 3103 36740 3148 36768
rect 2501 36731 2559 36737
rect 3142 36728 3148 36740
rect 3200 36728 3206 36780
rect 9030 36728 9036 36780
rect 9088 36768 9094 36780
rect 9309 36771 9367 36777
rect 9309 36768 9321 36771
rect 9088 36740 9321 36768
rect 9088 36728 9094 36740
rect 9309 36737 9321 36740
rect 9355 36737 9367 36771
rect 9309 36731 9367 36737
rect 11790 36728 11796 36780
rect 11848 36768 11854 36780
rect 13173 36771 13231 36777
rect 13173 36768 13185 36771
rect 11848 36740 13185 36768
rect 11848 36728 11854 36740
rect 13173 36737 13185 36740
rect 13219 36737 13231 36771
rect 13173 36731 13231 36737
rect 16758 36728 16764 36780
rect 16816 36768 16822 36780
rect 17880 36777 17908 36808
rect 28074 36796 28080 36848
rect 28132 36836 28138 36848
rect 38102 36836 38108 36848
rect 28132 36808 31616 36836
rect 38063 36808 38108 36836
rect 28132 36796 28138 36808
rect 17037 36771 17095 36777
rect 17037 36768 17049 36771
rect 16816 36740 17049 36768
rect 16816 36728 16822 36740
rect 17037 36737 17049 36740
rect 17083 36737 17095 36771
rect 17037 36731 17095 36737
rect 17865 36771 17923 36777
rect 17865 36737 17877 36771
rect 17911 36737 17923 36771
rect 19426 36768 19432 36780
rect 19387 36740 19432 36768
rect 17865 36731 17923 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 23474 36768 23480 36780
rect 23435 36740 23480 36768
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 28442 36768 28448 36780
rect 28403 36740 28448 36768
rect 28442 36728 28448 36740
rect 28500 36728 28506 36780
rect 31588 36777 31616 36808
rect 38102 36796 38108 36808
rect 38160 36796 38166 36848
rect 28721 36771 28779 36777
rect 28721 36737 28733 36771
rect 28767 36768 28779 36771
rect 29365 36771 29423 36777
rect 29365 36768 29377 36771
rect 28767 36740 29377 36768
rect 28767 36737 28779 36740
rect 28721 36731 28779 36737
rect 29365 36737 29377 36740
rect 29411 36737 29423 36771
rect 29365 36731 29423 36737
rect 31573 36771 31631 36777
rect 31573 36737 31585 36771
rect 31619 36737 31631 36771
rect 31573 36731 31631 36737
rect 35434 36728 35440 36780
rect 35492 36768 35498 36780
rect 35713 36771 35771 36777
rect 35713 36768 35725 36771
rect 35492 36740 35725 36768
rect 35492 36728 35498 36740
rect 35713 36737 35725 36740
rect 35759 36737 35771 36771
rect 36354 36768 36360 36780
rect 36315 36740 36360 36768
rect 35713 36731 35771 36737
rect 36354 36728 36360 36740
rect 36412 36728 36418 36780
rect 4614 36700 4620 36712
rect 1596 36672 4620 36700
rect 4614 36660 4620 36672
rect 4672 36660 4678 36712
rect 2317 36635 2375 36641
rect 2317 36601 2329 36635
rect 2363 36632 2375 36635
rect 6730 36632 6736 36644
rect 2363 36604 6736 36632
rect 2363 36601 2375 36604
rect 2317 36595 2375 36601
rect 6730 36592 6736 36604
rect 6788 36592 6794 36644
rect 12989 36635 13047 36641
rect 12989 36601 13001 36635
rect 13035 36632 13047 36635
rect 34882 36632 34888 36644
rect 13035 36604 34888 36632
rect 13035 36601 13047 36604
rect 12989 36595 13047 36601
rect 34882 36592 34888 36604
rect 34940 36592 34946 36644
rect 2961 36567 3019 36573
rect 2961 36533 2973 36567
rect 3007 36564 3019 36567
rect 5810 36564 5816 36576
rect 3007 36536 5816 36564
rect 3007 36533 3019 36536
rect 2961 36527 3019 36533
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 8018 36524 8024 36576
rect 8076 36564 8082 36576
rect 9125 36567 9183 36573
rect 9125 36564 9137 36567
rect 8076 36536 9137 36564
rect 8076 36524 8082 36536
rect 9125 36533 9137 36536
rect 9171 36533 9183 36567
rect 9125 36527 9183 36533
rect 15470 36524 15476 36576
rect 15528 36564 15534 36576
rect 16853 36567 16911 36573
rect 16853 36564 16865 36567
rect 15528 36536 16865 36564
rect 15528 36524 15534 36536
rect 16853 36533 16865 36536
rect 16899 36533 16911 36567
rect 16853 36527 16911 36533
rect 21634 36524 21640 36576
rect 21692 36564 21698 36576
rect 23293 36567 23351 36573
rect 23293 36564 23305 36567
rect 21692 36536 23305 36564
rect 21692 36524 21698 36536
rect 23293 36533 23305 36536
rect 23339 36533 23351 36567
rect 23293 36527 23351 36533
rect 33134 36524 33140 36576
rect 33192 36564 33198 36576
rect 35529 36567 35587 36573
rect 35529 36564 35541 36567
rect 33192 36536 35541 36564
rect 33192 36524 33198 36536
rect 35529 36533 35541 36536
rect 35575 36533 35587 36567
rect 35529 36527 35587 36533
rect 36449 36567 36507 36573
rect 36449 36533 36461 36567
rect 36495 36564 36507 36567
rect 36814 36564 36820 36576
rect 36495 36536 36820 36564
rect 36495 36533 36507 36536
rect 36449 36527 36507 36533
rect 36814 36524 36820 36536
rect 36872 36524 36878 36576
rect 37274 36524 37280 36576
rect 37332 36564 37338 36576
rect 38197 36567 38255 36573
rect 38197 36564 38209 36567
rect 37332 36536 38209 36564
rect 37332 36524 37338 36536
rect 38197 36533 38209 36536
rect 38243 36533 38255 36567
rect 38197 36527 38255 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 37461 36363 37519 36369
rect 37461 36329 37473 36363
rect 37507 36360 37519 36363
rect 39298 36360 39304 36372
rect 37507 36332 39304 36360
rect 37507 36329 37519 36332
rect 37461 36323 37519 36329
rect 39298 36320 39304 36332
rect 39356 36320 39362 36372
rect 36633 36295 36691 36301
rect 36633 36261 36645 36295
rect 36679 36261 36691 36295
rect 36633 36255 36691 36261
rect 36648 36224 36676 36255
rect 36648 36196 37320 36224
rect 1762 36156 1768 36168
rect 1723 36128 1768 36156
rect 1762 36116 1768 36128
rect 1820 36116 1826 36168
rect 36814 36156 36820 36168
rect 36775 36128 36820 36156
rect 36814 36116 36820 36128
rect 36872 36116 36878 36168
rect 37292 36165 37320 36196
rect 37277 36159 37335 36165
rect 37277 36125 37289 36159
rect 37323 36125 37335 36159
rect 37277 36119 37335 36125
rect 38013 36159 38071 36165
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 33318 36048 33324 36100
rect 33376 36088 33382 36100
rect 38028 36088 38056 36119
rect 33376 36060 38056 36088
rect 33376 36048 33382 36060
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 2682 36020 2688 36032
rect 1627 35992 2688 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 2682 35980 2688 35992
rect 2740 35980 2746 36032
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 12526 35816 12532 35828
rect 12487 35788 12532 35816
rect 12526 35776 12532 35788
rect 12584 35776 12590 35828
rect 38654 35748 38660 35760
rect 36924 35720 38660 35748
rect 658 35640 664 35692
rect 716 35680 722 35692
rect 1765 35683 1823 35689
rect 1765 35680 1777 35683
rect 716 35652 1777 35680
rect 716 35640 722 35652
rect 1765 35649 1777 35652
rect 1811 35649 1823 35683
rect 1765 35643 1823 35649
rect 12713 35683 12771 35689
rect 12713 35649 12725 35683
rect 12759 35680 12771 35683
rect 13906 35680 13912 35692
rect 12759 35652 13912 35680
rect 12759 35649 12771 35652
rect 12713 35643 12771 35649
rect 13906 35640 13912 35652
rect 13964 35640 13970 35692
rect 36924 35689 36952 35720
rect 38654 35708 38660 35720
rect 38712 35708 38718 35760
rect 36909 35683 36967 35689
rect 36909 35649 36921 35683
rect 36955 35649 36967 35683
rect 38010 35680 38016 35692
rect 37971 35652 38016 35680
rect 36909 35643 36967 35649
rect 38010 35640 38016 35652
rect 38068 35640 38074 35692
rect 1581 35479 1639 35485
rect 1581 35445 1593 35479
rect 1627 35476 1639 35479
rect 5718 35476 5724 35488
rect 1627 35448 5724 35476
rect 1627 35445 1639 35448
rect 1581 35439 1639 35445
rect 5718 35436 5724 35448
rect 5776 35436 5782 35488
rect 34514 35436 34520 35488
rect 34572 35476 34578 35488
rect 36725 35479 36783 35485
rect 36725 35476 36737 35479
rect 34572 35448 36737 35476
rect 34572 35436 34578 35448
rect 36725 35445 36737 35448
rect 36771 35445 36783 35479
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 36725 35439 36783 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 38286 35068 38292 35080
rect 38247 35040 38292 35068
rect 38286 35028 38292 35040
rect 38344 35028 38350 35080
rect 20622 34892 20628 34944
rect 20680 34932 20686 34944
rect 38105 34935 38163 34941
rect 38105 34932 38117 34935
rect 20680 34904 38117 34932
rect 20680 34892 20686 34904
rect 38105 34901 38117 34904
rect 38151 34901 38163 34935
rect 38105 34895 38163 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 33778 34552 33784 34604
rect 33836 34592 33842 34604
rect 38013 34595 38071 34601
rect 38013 34592 38025 34595
rect 33836 34564 38025 34592
rect 33836 34552 33842 34564
rect 38013 34561 38025 34564
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 19978 33804 19984 33856
rect 20036 33844 20042 33856
rect 37274 33844 37280 33856
rect 20036 33816 37280 33844
rect 20036 33804 20042 33816
rect 37274 33804 37280 33816
rect 37332 33804 37338 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 4525 33643 4583 33649
rect 4525 33609 4537 33643
rect 4571 33640 4583 33643
rect 4614 33640 4620 33652
rect 4571 33612 4620 33640
rect 4571 33609 4583 33612
rect 4525 33603 4583 33609
rect 4614 33600 4620 33612
rect 4672 33600 4678 33652
rect 4709 33507 4767 33513
rect 4709 33473 4721 33507
rect 4755 33504 4767 33507
rect 6638 33504 6644 33516
rect 4755 33476 6644 33504
rect 4755 33473 4767 33476
rect 4709 33467 4767 33473
rect 6638 33464 6644 33476
rect 6696 33464 6702 33516
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 28169 33099 28227 33105
rect 28169 33065 28181 33099
rect 28215 33096 28227 33099
rect 32398 33096 32404 33108
rect 28215 33068 32404 33096
rect 28215 33065 28227 33068
rect 28169 33059 28227 33065
rect 32398 33056 32404 33068
rect 32456 33056 32462 33108
rect 37369 33099 37427 33105
rect 37369 33065 37381 33099
rect 37415 33096 37427 33099
rect 38010 33096 38016 33108
rect 37415 33068 38016 33096
rect 37415 33065 37427 33068
rect 37369 33059 37427 33065
rect 38010 33056 38016 33068
rect 38068 33056 38074 33108
rect 1581 32895 1639 32901
rect 1581 32861 1593 32895
rect 1627 32892 1639 32895
rect 4157 32895 4215 32901
rect 1627 32864 4016 32892
rect 1627 32861 1639 32864
rect 1581 32855 1639 32861
rect 1762 32756 1768 32768
rect 1723 32728 1768 32756
rect 1762 32716 1768 32728
rect 1820 32716 1826 32768
rect 3988 32765 4016 32864
rect 4157 32861 4169 32895
rect 4203 32892 4215 32895
rect 5534 32892 5540 32904
rect 4203 32864 5540 32892
rect 4203 32861 4215 32864
rect 4157 32855 4215 32861
rect 5534 32852 5540 32864
rect 5592 32892 5598 32904
rect 6822 32892 6828 32904
rect 5592 32864 6828 32892
rect 5592 32852 5598 32864
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 28350 32892 28356 32904
rect 28311 32864 28356 32892
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 36814 32852 36820 32904
rect 36872 32892 36878 32904
rect 37553 32895 37611 32901
rect 37553 32892 37565 32895
rect 36872 32864 37565 32892
rect 36872 32852 36878 32864
rect 37553 32861 37565 32864
rect 37599 32861 37611 32895
rect 37553 32855 37611 32861
rect 38102 32824 38108 32836
rect 38063 32796 38108 32824
rect 38102 32784 38108 32796
rect 38160 32784 38166 32836
rect 3973 32759 4031 32765
rect 3973 32725 3985 32759
rect 4019 32725 4031 32759
rect 3973 32719 4031 32725
rect 37826 32716 37832 32768
rect 37884 32756 37890 32768
rect 38197 32759 38255 32765
rect 38197 32756 38209 32759
rect 37884 32728 38209 32756
rect 37884 32716 37890 32728
rect 38197 32725 38209 32728
rect 38243 32725 38255 32759
rect 38197 32719 38255 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 13906 32552 13912 32564
rect 13867 32524 13912 32552
rect 13906 32512 13912 32524
rect 13964 32512 13970 32564
rect 36814 32552 36820 32564
rect 36775 32524 36820 32552
rect 36814 32512 36820 32524
rect 36872 32512 36878 32564
rect 12342 32444 12348 32496
rect 12400 32484 12406 32496
rect 12400 32456 15332 32484
rect 12400 32444 12406 32456
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 2590 32416 2596 32428
rect 1627 32388 2596 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 2590 32376 2596 32388
rect 2648 32376 2654 32428
rect 13817 32419 13875 32425
rect 13817 32385 13829 32419
rect 13863 32416 13875 32419
rect 15010 32416 15016 32428
rect 13863 32388 15016 32416
rect 13863 32385 13875 32388
rect 13817 32379 13875 32385
rect 15010 32376 15016 32388
rect 15068 32376 15074 32428
rect 15304 32425 15332 32456
rect 15289 32419 15347 32425
rect 15289 32385 15301 32419
rect 15335 32385 15347 32419
rect 36722 32416 36728 32428
rect 36683 32388 36728 32416
rect 15289 32379 15347 32385
rect 36722 32376 36728 32388
rect 36780 32376 36786 32428
rect 38102 32416 38108 32428
rect 38063 32388 38108 32416
rect 38102 32376 38108 32388
rect 38160 32376 38166 32428
rect 3418 32240 3424 32292
rect 3476 32280 3482 32292
rect 20806 32280 20812 32292
rect 3476 32252 20812 32280
rect 3476 32240 3482 32252
rect 20806 32240 20812 32252
rect 20864 32240 20870 32292
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 15378 32212 15384 32224
rect 15339 32184 15384 32212
rect 15378 32172 15384 32184
rect 15436 32172 15442 32224
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 17034 31968 17040 32020
rect 17092 32008 17098 32020
rect 23017 32011 23075 32017
rect 23017 32008 23029 32011
rect 17092 31980 23029 32008
rect 17092 31968 17098 31980
rect 23017 31977 23029 31980
rect 23063 31977 23075 32011
rect 23017 31971 23075 31977
rect 23106 31968 23112 32020
rect 23164 32008 23170 32020
rect 23164 31980 35894 32008
rect 23164 31968 23170 31980
rect 11698 31900 11704 31952
rect 11756 31940 11762 31952
rect 35866 31940 35894 31980
rect 38194 31940 38200 31952
rect 11756 31912 26234 31940
rect 35866 31912 38200 31940
rect 11756 31900 11762 31912
rect 5905 31875 5963 31881
rect 5905 31841 5917 31875
rect 5951 31872 5963 31875
rect 10410 31872 10416 31884
rect 5951 31844 10416 31872
rect 5951 31841 5963 31844
rect 5905 31835 5963 31841
rect 10410 31832 10416 31844
rect 10468 31832 10474 31884
rect 18230 31832 18236 31884
rect 18288 31872 18294 31884
rect 19613 31875 19671 31881
rect 19613 31872 19625 31875
rect 18288 31844 19625 31872
rect 18288 31832 18294 31844
rect 19613 31841 19625 31844
rect 19659 31841 19671 31875
rect 19613 31835 19671 31841
rect 20070 31832 20076 31884
rect 20128 31872 20134 31884
rect 21729 31875 21787 31881
rect 21729 31872 21741 31875
rect 20128 31844 21741 31872
rect 20128 31832 20134 31844
rect 21729 31841 21741 31844
rect 21775 31841 21787 31875
rect 21729 31835 21787 31841
rect 5810 31804 5816 31816
rect 5771 31776 5816 31804
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 19521 31807 19579 31813
rect 19521 31773 19533 31807
rect 19567 31804 19579 31807
rect 20346 31804 20352 31816
rect 19567 31776 20352 31804
rect 19567 31773 19579 31776
rect 19521 31767 19579 31773
rect 20346 31764 20352 31776
rect 20404 31764 20410 31816
rect 20622 31804 20628 31816
rect 20583 31776 20628 31804
rect 20622 31764 20628 31776
rect 20680 31764 20686 31816
rect 20806 31804 20812 31816
rect 20767 31776 20812 31804
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 21634 31804 21640 31816
rect 21595 31776 21640 31804
rect 21634 31764 21640 31776
rect 21692 31764 21698 31816
rect 22925 31807 22983 31813
rect 22925 31773 22937 31807
rect 22971 31804 22983 31807
rect 23014 31804 23020 31816
rect 22971 31776 23020 31804
rect 22971 31773 22983 31776
rect 22925 31767 22983 31773
rect 23014 31764 23020 31776
rect 23072 31764 23078 31816
rect 26206 31804 26234 31912
rect 38194 31900 38200 31912
rect 38252 31900 38258 31952
rect 26697 31807 26755 31813
rect 26697 31804 26709 31807
rect 26206 31776 26709 31804
rect 26697 31773 26709 31776
rect 26743 31773 26755 31807
rect 26697 31767 26755 31773
rect 26510 31668 26516 31680
rect 26471 31640 26516 31668
rect 26510 31628 26516 31640
rect 26568 31628 26574 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 33318 31464 33324 31476
rect 33279 31436 33324 31464
rect 33318 31424 33324 31436
rect 33376 31424 33382 31476
rect 5718 31328 5724 31340
rect 5679 31300 5724 31328
rect 5718 31288 5724 31300
rect 5776 31288 5782 31340
rect 25685 31331 25743 31337
rect 25685 31297 25697 31331
rect 25731 31328 25743 31331
rect 29822 31328 29828 31340
rect 25731 31300 29828 31328
rect 25731 31297 25743 31300
rect 25685 31291 25743 31297
rect 29822 31288 29828 31300
rect 29880 31288 29886 31340
rect 32398 31288 32404 31340
rect 32456 31328 32462 31340
rect 33505 31331 33563 31337
rect 33505 31328 33517 31331
rect 32456 31300 33517 31328
rect 32456 31288 32462 31300
rect 33505 31297 33517 31300
rect 33551 31297 33563 31331
rect 33505 31291 33563 31297
rect 5813 31127 5871 31133
rect 5813 31093 5825 31127
rect 5859 31124 5871 31127
rect 6086 31124 6092 31136
rect 5859 31096 6092 31124
rect 5859 31093 5871 31096
rect 5813 31087 5871 31093
rect 6086 31084 6092 31096
rect 6144 31084 6150 31136
rect 24026 31084 24032 31136
rect 24084 31124 24090 31136
rect 25777 31127 25835 31133
rect 25777 31124 25789 31127
rect 24084 31096 25789 31124
rect 24084 31084 24090 31096
rect 25777 31093 25789 31096
rect 25823 31093 25835 31127
rect 25777 31087 25835 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 11146 30784 11152 30796
rect 1596 30756 11152 30784
rect 1596 30725 1624 30756
rect 11146 30744 11152 30756
rect 11204 30744 11210 30796
rect 33134 30784 33140 30796
rect 29748 30756 33140 30784
rect 1581 30719 1639 30725
rect 1581 30685 1593 30719
rect 1627 30685 1639 30719
rect 1581 30679 1639 30685
rect 2682 30676 2688 30728
rect 2740 30716 2746 30728
rect 6825 30719 6883 30725
rect 6825 30716 6837 30719
rect 2740 30688 6837 30716
rect 2740 30676 2746 30688
rect 6825 30685 6837 30688
rect 6871 30685 6883 30719
rect 8018 30716 8024 30728
rect 7979 30688 8024 30716
rect 6825 30679 6883 30685
rect 8018 30676 8024 30688
rect 8076 30676 8082 30728
rect 11054 30716 11060 30728
rect 11015 30688 11060 30716
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 29748 30725 29776 30756
rect 33134 30744 33140 30756
rect 33192 30744 33198 30796
rect 29733 30719 29791 30725
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 30469 30719 30527 30725
rect 30469 30685 30481 30719
rect 30515 30716 30527 30719
rect 34514 30716 34520 30728
rect 30515 30688 34520 30716
rect 30515 30685 30527 30688
rect 30469 30679 30527 30685
rect 34514 30676 34520 30688
rect 34572 30676 34578 30728
rect 38010 30716 38016 30728
rect 37971 30688 38016 30716
rect 38010 30676 38016 30688
rect 38068 30676 38074 30728
rect 6917 30651 6975 30657
rect 6917 30617 6929 30651
rect 6963 30648 6975 30651
rect 10962 30648 10968 30660
rect 6963 30620 10968 30648
rect 6963 30617 6975 30620
rect 6917 30611 6975 30617
rect 10962 30608 10968 30620
rect 11020 30608 11026 30660
rect 30561 30651 30619 30657
rect 30561 30648 30573 30651
rect 26206 30620 30573 30648
rect 1762 30580 1768 30592
rect 1723 30552 1768 30580
rect 1762 30540 1768 30552
rect 1820 30540 1826 30592
rect 8113 30583 8171 30589
rect 8113 30549 8125 30583
rect 8159 30580 8171 30583
rect 8202 30580 8208 30592
rect 8159 30552 8208 30580
rect 8159 30549 8171 30552
rect 8113 30543 8171 30549
rect 8202 30540 8208 30552
rect 8260 30540 8266 30592
rect 11149 30583 11207 30589
rect 11149 30549 11161 30583
rect 11195 30580 11207 30583
rect 13354 30580 13360 30592
rect 11195 30552 13360 30580
rect 11195 30549 11207 30552
rect 11149 30543 11207 30549
rect 13354 30540 13360 30552
rect 13412 30540 13418 30592
rect 24946 30540 24952 30592
rect 25004 30580 25010 30592
rect 26206 30580 26234 30620
rect 30561 30617 30573 30620
rect 30607 30617 30619 30651
rect 30561 30611 30619 30617
rect 29822 30580 29828 30592
rect 25004 30552 26234 30580
rect 29783 30552 29828 30580
rect 25004 30540 25010 30552
rect 29822 30540 29828 30552
rect 29880 30540 29886 30592
rect 38194 30580 38200 30592
rect 38155 30552 38200 30580
rect 38194 30540 38200 30552
rect 38252 30540 38258 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 23566 30336 23572 30388
rect 23624 30376 23630 30388
rect 23624 30348 25452 30376
rect 23624 30336 23630 30348
rect 6638 30308 6644 30320
rect 6599 30280 6644 30308
rect 6638 30268 6644 30280
rect 6696 30268 6702 30320
rect 3881 30243 3939 30249
rect 3881 30209 3893 30243
rect 3927 30240 3939 30243
rect 5994 30240 6000 30252
rect 3927 30212 6000 30240
rect 3927 30209 3939 30212
rect 3881 30203 3939 30209
rect 5994 30200 6000 30212
rect 6052 30200 6058 30252
rect 6549 30243 6607 30249
rect 6549 30209 6561 30243
rect 6595 30240 6607 30243
rect 10502 30240 10508 30252
rect 6595 30212 10508 30240
rect 6595 30209 6607 30212
rect 6549 30203 6607 30209
rect 10502 30200 10508 30212
rect 10560 30200 10566 30252
rect 13265 30243 13323 30249
rect 13265 30209 13277 30243
rect 13311 30240 13323 30243
rect 17862 30240 17868 30252
rect 13311 30212 17868 30240
rect 13311 30209 13323 30212
rect 13265 30203 13323 30209
rect 17862 30200 17868 30212
rect 17920 30240 17926 30252
rect 24854 30240 24860 30252
rect 17920 30212 24860 30240
rect 17920 30200 17926 30212
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 25424 30249 25452 30348
rect 25409 30243 25467 30249
rect 25409 30209 25421 30243
rect 25455 30209 25467 30243
rect 27154 30240 27160 30252
rect 27115 30212 27160 30240
rect 25409 30203 25467 30209
rect 27154 30200 27160 30212
rect 27212 30200 27218 30252
rect 1578 30064 1584 30116
rect 1636 30104 1642 30116
rect 3697 30107 3755 30113
rect 3697 30104 3709 30107
rect 1636 30076 3709 30104
rect 1636 30064 1642 30076
rect 3697 30073 3709 30076
rect 3743 30073 3755 30107
rect 3697 30067 3755 30073
rect 11146 30064 11152 30116
rect 11204 30104 11210 30116
rect 13081 30107 13139 30113
rect 13081 30104 13093 30107
rect 11204 30076 13093 30104
rect 11204 30064 11210 30076
rect 13081 30073 13093 30076
rect 13127 30073 13139 30107
rect 13081 30067 13139 30073
rect 25225 30107 25283 30113
rect 25225 30073 25237 30107
rect 25271 30104 25283 30107
rect 38010 30104 38016 30116
rect 25271 30076 38016 30104
rect 25271 30073 25283 30076
rect 25225 30067 25283 30073
rect 38010 30064 38016 30076
rect 38068 30064 38074 30116
rect 25958 29996 25964 30048
rect 26016 30036 26022 30048
rect 27249 30039 27307 30045
rect 27249 30036 27261 30039
rect 26016 30008 27261 30036
rect 26016 29996 26022 30008
rect 27249 30005 27261 30008
rect 27295 30005 27307 30039
rect 27249 29999 27307 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 33778 29832 33784 29844
rect 33739 29804 33784 29832
rect 33778 29792 33784 29804
rect 33836 29792 33842 29844
rect 5258 29656 5264 29708
rect 5316 29696 5322 29708
rect 5316 29668 10640 29696
rect 5316 29656 5322 29668
rect 1762 29628 1768 29640
rect 1723 29600 1768 29628
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 6730 29588 6736 29640
rect 6788 29628 6794 29640
rect 10612 29637 10640 29668
rect 7837 29631 7895 29637
rect 7837 29628 7849 29631
rect 6788 29600 7849 29628
rect 6788 29588 6794 29600
rect 7837 29597 7849 29600
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 16574 29588 16580 29640
rect 16632 29628 16638 29640
rect 26326 29628 26332 29640
rect 16632 29600 26332 29628
rect 16632 29588 16638 29600
rect 26326 29588 26332 29600
rect 26384 29588 26390 29640
rect 32490 29588 32496 29640
rect 32548 29628 32554 29640
rect 33965 29631 34023 29637
rect 33965 29628 33977 29631
rect 32548 29600 33977 29628
rect 32548 29588 32554 29600
rect 33965 29597 33977 29600
rect 34011 29597 34023 29631
rect 33965 29591 34023 29597
rect 35434 29588 35440 29640
rect 35492 29628 35498 29640
rect 38013 29631 38071 29637
rect 38013 29628 38025 29631
rect 35492 29600 38025 29628
rect 35492 29588 35498 29600
rect 38013 29597 38025 29600
rect 38059 29597 38071 29631
rect 38013 29591 38071 29597
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 5626 29492 5632 29504
rect 1627 29464 5632 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 5626 29452 5632 29464
rect 5684 29452 5690 29504
rect 7006 29452 7012 29504
rect 7064 29492 7070 29504
rect 7929 29495 7987 29501
rect 7929 29492 7941 29495
rect 7064 29464 7941 29492
rect 7064 29452 7070 29464
rect 7929 29461 7941 29464
rect 7975 29461 7987 29495
rect 10686 29492 10692 29504
rect 10647 29464 10692 29492
rect 7929 29455 7987 29461
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 38194 29492 38200 29504
rect 38155 29464 38200 29492
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29152 1639 29155
rect 2314 29152 2320 29164
rect 1627 29124 2320 29152
rect 1627 29121 1639 29124
rect 1581 29115 1639 29121
rect 2314 29112 2320 29124
rect 2372 29112 2378 29164
rect 14090 29112 14096 29164
rect 14148 29152 14154 29164
rect 14553 29155 14611 29161
rect 14553 29152 14565 29155
rect 14148 29124 14565 29152
rect 14148 29112 14154 29124
rect 14553 29121 14565 29124
rect 14599 29121 14611 29155
rect 15470 29152 15476 29164
rect 15431 29124 15476 29152
rect 14553 29115 14611 29121
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 36262 29112 36268 29164
rect 36320 29152 36326 29164
rect 38013 29155 38071 29161
rect 38013 29152 38025 29155
rect 36320 29124 38025 29152
rect 36320 29112 36326 29124
rect 38013 29121 38025 29124
rect 38059 29121 38071 29155
rect 38013 29115 38071 29121
rect 14645 29087 14703 29093
rect 14645 29053 14657 29087
rect 14691 29084 14703 29087
rect 15930 29084 15936 29096
rect 14691 29056 15936 29084
rect 14691 29053 14703 29056
rect 14645 29047 14703 29053
rect 15930 29044 15936 29056
rect 15988 29044 15994 29096
rect 1762 29016 1768 29028
rect 1723 28988 1768 29016
rect 1762 28976 1768 28988
rect 1820 28976 1826 29028
rect 15194 28976 15200 29028
rect 15252 29016 15258 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 15252 28988 15577 29016
rect 15252 28976 15258 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 38194 29016 38200 29028
rect 38155 28988 38200 29016
rect 15565 28979 15623 28985
rect 38194 28976 38200 28988
rect 38252 28976 38258 29028
rect 17310 28908 17316 28960
rect 17368 28948 17374 28960
rect 23106 28948 23112 28960
rect 17368 28920 23112 28948
rect 17368 28908 17374 28920
rect 23106 28908 23112 28920
rect 23164 28908 23170 28960
rect 27706 28908 27712 28960
rect 27764 28948 27770 28960
rect 35526 28948 35532 28960
rect 27764 28920 35532 28948
rect 27764 28908 27770 28920
rect 35526 28908 35532 28920
rect 35584 28908 35590 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 11790 28500 11796 28552
rect 11848 28540 11854 28552
rect 11885 28543 11943 28549
rect 11885 28540 11897 28543
rect 11848 28512 11897 28540
rect 11848 28500 11854 28512
rect 11885 28509 11897 28512
rect 11931 28509 11943 28543
rect 18046 28540 18052 28552
rect 18007 28512 18052 28540
rect 11885 28503 11943 28509
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 11977 28407 12035 28413
rect 11977 28373 11989 28407
rect 12023 28404 12035 28407
rect 14090 28404 14096 28416
rect 12023 28376 14096 28404
rect 12023 28373 12035 28376
rect 11977 28367 12035 28373
rect 14090 28364 14096 28376
rect 14148 28364 14154 28416
rect 18138 28404 18144 28416
rect 18099 28376 18144 28404
rect 18138 28364 18144 28376
rect 18196 28364 18202 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 35069 28203 35127 28209
rect 35069 28169 35081 28203
rect 35115 28200 35127 28203
rect 36262 28200 36268 28212
rect 35115 28172 36268 28200
rect 35115 28169 35127 28172
rect 35069 28163 35127 28169
rect 36262 28160 36268 28172
rect 36320 28160 36326 28212
rect 15197 28067 15255 28073
rect 15197 28033 15209 28067
rect 15243 28064 15255 28067
rect 15562 28064 15568 28076
rect 15243 28036 15568 28064
rect 15243 28033 15255 28036
rect 15197 28027 15255 28033
rect 15562 28024 15568 28036
rect 15620 28024 15626 28076
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28064 23719 28067
rect 28074 28064 28080 28076
rect 23707 28036 28080 28064
rect 23707 28033 23719 28036
rect 23661 28027 23719 28033
rect 28074 28024 28080 28036
rect 28132 28024 28138 28076
rect 35253 28067 35311 28073
rect 35253 28033 35265 28067
rect 35299 28064 35311 28067
rect 35342 28064 35348 28076
rect 35299 28036 35348 28064
rect 35299 28033 35311 28036
rect 35253 28027 35311 28033
rect 35342 28024 35348 28036
rect 35400 28024 35406 28076
rect 14550 27820 14556 27872
rect 14608 27860 14614 27872
rect 15289 27863 15347 27869
rect 15289 27860 15301 27863
rect 14608 27832 15301 27860
rect 14608 27820 14614 27832
rect 15289 27829 15301 27832
rect 15335 27829 15347 27863
rect 15289 27823 15347 27829
rect 22094 27820 22100 27872
rect 22152 27860 22158 27872
rect 23753 27863 23811 27869
rect 23753 27860 23765 27863
rect 22152 27832 23765 27860
rect 22152 27820 22158 27832
rect 23753 27829 23765 27832
rect 23799 27829 23811 27863
rect 23753 27823 23811 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1762 27452 1768 27464
rect 1723 27424 1768 27452
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 38286 27452 38292 27464
rect 38247 27424 38292 27452
rect 38286 27412 38292 27424
rect 38344 27412 38350 27464
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 4062 27316 4068 27328
rect 1627 27288 4068 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 37366 27276 37372 27328
rect 37424 27316 37430 27328
rect 38105 27319 38163 27325
rect 38105 27316 38117 27319
rect 37424 27288 38117 27316
rect 37424 27276 37430 27288
rect 38105 27285 38117 27288
rect 38151 27285 38163 27319
rect 38105 27279 38163 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 5994 27072 6000 27124
rect 6052 27112 6058 27124
rect 6825 27115 6883 27121
rect 6825 27112 6837 27115
rect 6052 27084 6837 27112
rect 6052 27072 6058 27084
rect 6825 27081 6837 27084
rect 6871 27081 6883 27115
rect 6825 27075 6883 27081
rect 22462 27072 22468 27124
rect 22520 27112 22526 27124
rect 29822 27112 29828 27124
rect 22520 27084 29828 27112
rect 22520 27072 22526 27084
rect 29822 27072 29828 27084
rect 29880 27072 29886 27124
rect 35342 27112 35348 27124
rect 35303 27084 35348 27112
rect 35342 27072 35348 27084
rect 35400 27072 35406 27124
rect 16298 27004 16304 27056
rect 16356 27044 16362 27056
rect 28442 27044 28448 27056
rect 16356 27016 28448 27044
rect 16356 27004 16362 27016
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 37734 27044 37740 27056
rect 31036 27016 37740 27044
rect 6733 26979 6791 26985
rect 6733 26945 6745 26979
rect 6779 26976 6791 26979
rect 7098 26976 7104 26988
rect 6779 26948 7104 26976
rect 6779 26945 6791 26948
rect 6733 26939 6791 26945
rect 7098 26936 7104 26948
rect 7156 26936 7162 26988
rect 12434 26936 12440 26988
rect 12492 26976 12498 26988
rect 12989 26979 13047 26985
rect 12989 26976 13001 26979
rect 12492 26948 13001 26976
rect 12492 26936 12498 26948
rect 12989 26945 13001 26948
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26976 13691 26979
rect 15102 26976 15108 26988
rect 13679 26948 15108 26976
rect 13679 26945 13691 26948
rect 13633 26939 13691 26945
rect 15102 26936 15108 26948
rect 15160 26936 15166 26988
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26976 22155 26979
rect 31036 26976 31064 27016
rect 37734 27004 37740 27016
rect 37792 27004 37798 27056
rect 22143 26948 31064 26976
rect 35253 26979 35311 26985
rect 22143 26945 22155 26948
rect 22097 26939 22155 26945
rect 35253 26945 35265 26979
rect 35299 26945 35311 26979
rect 35253 26939 35311 26945
rect 20530 26868 20536 26920
rect 20588 26908 20594 26920
rect 35268 26908 35296 26939
rect 20588 26880 35296 26908
rect 20588 26868 20594 26880
rect 2590 26800 2596 26852
rect 2648 26840 2654 26852
rect 22281 26843 22339 26849
rect 22281 26840 22293 26843
rect 2648 26812 22293 26840
rect 2648 26800 2654 26812
rect 22281 26809 22293 26812
rect 22327 26809 22339 26843
rect 22281 26803 22339 26809
rect 12802 26772 12808 26784
rect 12763 26744 12808 26772
rect 12802 26732 12808 26744
rect 12860 26732 12866 26784
rect 13449 26775 13507 26781
rect 13449 26741 13461 26775
rect 13495 26772 13507 26775
rect 13722 26772 13728 26784
rect 13495 26744 13728 26772
rect 13495 26741 13507 26744
rect 13449 26735 13507 26741
rect 13722 26732 13728 26744
rect 13780 26732 13786 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 20346 26568 20352 26580
rect 12268 26540 20352 26568
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 5534 26500 5540 26512
rect 1627 26472 5540 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 5534 26460 5540 26472
rect 5592 26460 5598 26512
rect 1762 26364 1768 26376
rect 1723 26336 1768 26364
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 5718 26324 5724 26376
rect 5776 26364 5782 26376
rect 12161 26367 12219 26373
rect 12161 26364 12173 26367
rect 5776 26336 12173 26364
rect 5776 26324 5782 26336
rect 12161 26333 12173 26336
rect 12207 26333 12219 26367
rect 12161 26327 12219 26333
rect 11514 26256 11520 26308
rect 11572 26296 11578 26308
rect 12268 26305 12296 26540
rect 20346 26528 20352 26540
rect 20404 26528 20410 26580
rect 34885 26571 34943 26577
rect 34885 26537 34897 26571
rect 34931 26568 34943 26571
rect 35434 26568 35440 26580
rect 34931 26540 35440 26568
rect 34931 26537 34943 26540
rect 34885 26531 34943 26537
rect 35434 26528 35440 26540
rect 35492 26528 35498 26580
rect 13541 26503 13599 26509
rect 13541 26469 13553 26503
rect 13587 26500 13599 26503
rect 13998 26500 14004 26512
rect 13587 26472 14004 26500
rect 13587 26469 13599 26472
rect 13541 26463 13599 26469
rect 13998 26460 14004 26472
rect 14056 26460 14062 26512
rect 15013 26503 15071 26509
rect 15013 26469 15025 26503
rect 15059 26500 15071 26503
rect 15562 26500 15568 26512
rect 15059 26472 15568 26500
rect 15059 26469 15071 26472
rect 15013 26463 15071 26469
rect 15562 26460 15568 26472
rect 15620 26460 15626 26512
rect 15657 26503 15715 26509
rect 15657 26469 15669 26503
rect 15703 26469 15715 26503
rect 15657 26463 15715 26469
rect 12434 26392 12440 26444
rect 12492 26432 12498 26444
rect 12492 26404 14320 26432
rect 12492 26392 12498 26404
rect 13722 26364 13728 26376
rect 13683 26336 13728 26364
rect 13722 26324 13728 26336
rect 13780 26324 13786 26376
rect 14292 26373 14320 26404
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 15197 26367 15255 26373
rect 15197 26333 15209 26367
rect 15243 26364 15255 26367
rect 15672 26364 15700 26463
rect 15243 26336 15700 26364
rect 15841 26367 15899 26373
rect 15243 26333 15255 26336
rect 15197 26327 15255 26333
rect 15841 26333 15853 26367
rect 15887 26333 15899 26367
rect 15841 26327 15899 26333
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26364 18107 26367
rect 19058 26364 19064 26376
rect 18095 26336 19064 26364
rect 18095 26333 18107 26336
rect 18049 26327 18107 26333
rect 12253 26299 12311 26305
rect 12253 26296 12265 26299
rect 11572 26268 12265 26296
rect 11572 26256 11578 26268
rect 12253 26265 12265 26268
rect 12299 26265 12311 26299
rect 14366 26296 14372 26308
rect 14327 26268 14372 26296
rect 12253 26259 12311 26265
rect 14366 26256 14372 26268
rect 14424 26256 14430 26308
rect 15102 26256 15108 26308
rect 15160 26296 15166 26308
rect 15856 26296 15884 26327
rect 19058 26324 19064 26336
rect 19116 26324 19122 26376
rect 29178 26324 29184 26376
rect 29236 26364 29242 26376
rect 35069 26367 35127 26373
rect 35069 26364 35081 26367
rect 29236 26336 35081 26364
rect 29236 26324 29242 26336
rect 35069 26333 35081 26336
rect 35115 26333 35127 26367
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 35069 26327 35127 26333
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 15160 26268 15884 26296
rect 15160 26256 15166 26268
rect 17218 26188 17224 26240
rect 17276 26228 17282 26240
rect 17865 26231 17923 26237
rect 17865 26228 17877 26231
rect 17276 26200 17877 26228
rect 17276 26188 17282 26200
rect 17865 26197 17877 26200
rect 17911 26197 17923 26231
rect 38102 26228 38108 26240
rect 38063 26200 38108 26228
rect 17865 26191 17923 26197
rect 38102 26188 38108 26200
rect 38160 26188 38166 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 28077 26027 28135 26033
rect 28077 25993 28089 26027
rect 28123 26024 28135 26027
rect 32398 26024 32404 26036
rect 28123 25996 32404 26024
rect 28123 25993 28135 25996
rect 28077 25987 28135 25993
rect 32398 25984 32404 25996
rect 32456 25984 32462 26036
rect 12802 25848 12808 25900
rect 12860 25888 12866 25900
rect 13725 25891 13783 25897
rect 13725 25888 13737 25891
rect 12860 25860 13737 25888
rect 12860 25848 12866 25860
rect 13725 25857 13737 25860
rect 13771 25857 13783 25891
rect 17862 25888 17868 25900
rect 17823 25860 17868 25888
rect 13725 25851 13783 25857
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 18877 25891 18935 25897
rect 18877 25857 18889 25891
rect 18923 25888 18935 25891
rect 19058 25888 19064 25900
rect 18923 25860 19064 25888
rect 18923 25857 18935 25860
rect 18877 25851 18935 25857
rect 19058 25848 19064 25860
rect 19116 25848 19122 25900
rect 27062 25848 27068 25900
rect 27120 25888 27126 25900
rect 27985 25891 28043 25897
rect 27985 25888 27997 25891
rect 27120 25860 27997 25888
rect 27120 25848 27126 25860
rect 27985 25857 27997 25860
rect 28031 25857 28043 25891
rect 27985 25851 28043 25857
rect 13541 25687 13599 25693
rect 13541 25653 13553 25687
rect 13587 25684 13599 25687
rect 14458 25684 14464 25696
rect 13587 25656 14464 25684
rect 13587 25653 13599 25656
rect 13541 25647 13599 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 17957 25687 18015 25693
rect 17957 25653 17969 25687
rect 18003 25684 18015 25687
rect 18046 25684 18052 25696
rect 18003 25656 18052 25684
rect 18003 25653 18015 25656
rect 17957 25647 18015 25653
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 18322 25644 18328 25696
rect 18380 25684 18386 25696
rect 18969 25687 19027 25693
rect 18969 25684 18981 25687
rect 18380 25656 18981 25684
rect 18380 25644 18386 25656
rect 18969 25653 18981 25656
rect 19015 25653 19027 25687
rect 18969 25647 19027 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 28077 25483 28135 25489
rect 28077 25449 28089 25483
rect 28123 25480 28135 25483
rect 32490 25480 32496 25492
rect 28123 25452 32496 25480
rect 28123 25449 28135 25452
rect 28077 25443 28135 25449
rect 32490 25440 32496 25452
rect 32548 25440 32554 25492
rect 2682 25372 2688 25424
rect 2740 25412 2746 25424
rect 3418 25412 3424 25424
rect 2740 25384 3424 25412
rect 2740 25372 2746 25384
rect 3418 25372 3424 25384
rect 3476 25372 3482 25424
rect 21634 25344 21640 25356
rect 15488 25316 21640 25344
rect 14182 25236 14188 25288
rect 14240 25276 14246 25288
rect 15488 25285 15516 25316
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 14240 25248 14289 25276
rect 14240 25236 14246 25248
rect 14277 25245 14289 25248
rect 14323 25245 14335 25279
rect 14277 25239 14335 25245
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25245 16175 25279
rect 17218 25276 17224 25288
rect 17179 25248 17224 25276
rect 16117 25239 16175 25245
rect 11238 25168 11244 25220
rect 11296 25208 11302 25220
rect 13078 25208 13084 25220
rect 11296 25180 13084 25208
rect 11296 25168 11302 25180
rect 13078 25168 13084 25180
rect 13136 25208 13142 25220
rect 16132 25208 16160 25239
rect 17218 25236 17224 25248
rect 17276 25236 17282 25288
rect 27982 25276 27988 25288
rect 27943 25248 27988 25276
rect 27982 25236 27988 25248
rect 28040 25236 28046 25288
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 13136 25180 16160 25208
rect 13136 25168 13142 25180
rect 18046 25168 18052 25220
rect 18104 25208 18110 25220
rect 18233 25211 18291 25217
rect 18233 25208 18245 25211
rect 18104 25180 18245 25208
rect 18104 25168 18110 25180
rect 18233 25177 18245 25180
rect 18279 25177 18291 25211
rect 18233 25171 18291 25177
rect 18322 25168 18328 25220
rect 18380 25208 18386 25220
rect 18877 25211 18935 25217
rect 18380 25180 18425 25208
rect 18380 25168 18386 25180
rect 18877 25177 18889 25211
rect 18923 25208 18935 25211
rect 19334 25208 19340 25220
rect 18923 25180 19340 25208
rect 18923 25177 18935 25180
rect 18877 25171 18935 25177
rect 19334 25168 19340 25180
rect 19392 25168 19398 25220
rect 13906 25100 13912 25152
rect 13964 25140 13970 25152
rect 14369 25143 14427 25149
rect 14369 25140 14381 25143
rect 13964 25112 14381 25140
rect 13964 25100 13970 25112
rect 14369 25109 14381 25112
rect 14415 25109 14427 25143
rect 14369 25103 14427 25109
rect 15286 25100 15292 25152
rect 15344 25140 15350 25152
rect 15565 25143 15623 25149
rect 15565 25140 15577 25143
rect 15344 25112 15577 25140
rect 15344 25100 15350 25112
rect 15565 25109 15577 25112
rect 15611 25109 15623 25143
rect 15565 25103 15623 25109
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16942 25140 16948 25152
rect 16255 25112 16948 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 17037 25143 17095 25149
rect 17037 25109 17049 25143
rect 17083 25140 17095 25143
rect 17126 25140 17132 25152
rect 17083 25112 17132 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17126 25100 17132 25112
rect 17184 25100 17190 25152
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 14366 24868 14372 24880
rect 14327 24840 14372 24868
rect 14366 24828 14372 24840
rect 14424 24828 14430 24880
rect 16942 24828 16948 24880
rect 17000 24868 17006 24880
rect 17037 24871 17095 24877
rect 17037 24868 17049 24871
rect 17000 24840 17049 24868
rect 17000 24828 17006 24840
rect 17037 24837 17049 24840
rect 17083 24837 17095 24871
rect 17037 24831 17095 24837
rect 1578 24800 1584 24812
rect 1539 24772 1584 24800
rect 1578 24760 1584 24772
rect 1636 24760 1642 24812
rect 5626 24760 5632 24812
rect 5684 24800 5690 24812
rect 7377 24803 7435 24809
rect 7377 24800 7389 24803
rect 5684 24772 7389 24800
rect 5684 24760 5690 24772
rect 7377 24769 7389 24772
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 9030 24760 9036 24812
rect 9088 24800 9094 24812
rect 9217 24803 9275 24809
rect 9217 24800 9229 24803
rect 9088 24772 9229 24800
rect 9088 24760 9094 24772
rect 9217 24769 9229 24772
rect 9263 24769 9275 24803
rect 9217 24763 9275 24769
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24800 14979 24803
rect 15010 24800 15016 24812
rect 14967 24772 15016 24800
rect 14967 24769 14979 24772
rect 14921 24763 14979 24769
rect 15010 24760 15016 24772
rect 15068 24760 15074 24812
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 15473 24803 15531 24809
rect 15473 24800 15485 24803
rect 15436 24772 15485 24800
rect 15436 24760 15442 24772
rect 15473 24769 15485 24772
rect 15519 24769 15531 24803
rect 15473 24763 15531 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 22738 24800 22744 24812
rect 22699 24772 22744 24800
rect 16117 24763 16175 24769
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24732 13599 24735
rect 13814 24732 13820 24744
rect 13587 24704 13820 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 13814 24692 13820 24704
rect 13872 24692 13878 24744
rect 14277 24735 14335 24741
rect 14277 24701 14289 24735
rect 14323 24732 14335 24735
rect 15838 24732 15844 24744
rect 14323 24704 15844 24732
rect 14323 24701 14335 24704
rect 14277 24695 14335 24701
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 7469 24667 7527 24673
rect 7469 24633 7481 24667
rect 7515 24664 7527 24667
rect 9582 24664 9588 24676
rect 7515 24636 9588 24664
rect 7515 24633 7527 24636
rect 7469 24627 7527 24633
rect 9582 24624 9588 24636
rect 9640 24624 9646 24676
rect 14182 24624 14188 24676
rect 14240 24664 14246 24676
rect 15102 24664 15108 24676
rect 14240 24636 15108 24664
rect 14240 24624 14246 24636
rect 15102 24624 15108 24636
rect 15160 24664 15166 24676
rect 16132 24664 16160 24763
rect 22738 24760 22744 24772
rect 22796 24760 22802 24812
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24769 23443 24803
rect 23385 24763 23443 24769
rect 16945 24735 17003 24741
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 18046 24732 18052 24744
rect 16991 24704 18052 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 23400 24732 23428 24763
rect 22572 24704 23428 24732
rect 15160 24636 16160 24664
rect 17497 24667 17555 24673
rect 15160 24624 15166 24636
rect 17497 24633 17509 24667
rect 17543 24664 17555 24667
rect 17954 24664 17960 24676
rect 17543 24636 17960 24664
rect 17543 24633 17555 24636
rect 17497 24627 17555 24633
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 22572 24673 22600 24704
rect 22557 24667 22615 24673
rect 22557 24633 22569 24667
rect 22603 24633 22615 24667
rect 22557 24627 22615 24633
rect 1762 24596 1768 24608
rect 1723 24568 1768 24596
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 9033 24599 9091 24605
rect 9033 24565 9045 24599
rect 9079 24596 9091 24599
rect 10134 24596 10140 24608
rect 9079 24568 10140 24596
rect 9079 24565 9091 24568
rect 9033 24559 9091 24565
rect 10134 24556 10140 24568
rect 10192 24556 10198 24608
rect 10226 24556 10232 24608
rect 10284 24596 10290 24608
rect 10686 24596 10692 24608
rect 10284 24568 10692 24596
rect 10284 24556 10290 24568
rect 10686 24556 10692 24568
rect 10744 24596 10750 24608
rect 15470 24596 15476 24608
rect 10744 24568 15476 24596
rect 10744 24556 10750 24568
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 15565 24599 15623 24605
rect 15565 24565 15577 24599
rect 15611 24596 15623 24599
rect 15746 24596 15752 24608
rect 15611 24568 15752 24596
rect 15611 24565 15623 24568
rect 15565 24559 15623 24565
rect 15746 24556 15752 24568
rect 15804 24556 15810 24608
rect 16209 24599 16267 24605
rect 16209 24565 16221 24599
rect 16255 24596 16267 24599
rect 16942 24596 16948 24608
rect 16255 24568 16948 24596
rect 16255 24565 16267 24568
rect 16209 24559 16267 24565
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 22830 24556 22836 24608
rect 22888 24596 22894 24608
rect 23201 24599 23259 24605
rect 23201 24596 23213 24599
rect 22888 24568 23213 24596
rect 22888 24556 22894 24568
rect 23201 24565 23213 24568
rect 23247 24565 23259 24599
rect 23201 24559 23259 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1578 24352 1584 24404
rect 1636 24392 1642 24404
rect 30742 24392 30748 24404
rect 1636 24364 30748 24392
rect 1636 24352 1642 24364
rect 30742 24352 30748 24364
rect 30800 24352 30806 24404
rect 10689 24327 10747 24333
rect 10689 24293 10701 24327
rect 10735 24324 10747 24327
rect 12158 24324 12164 24336
rect 10735 24296 12164 24324
rect 10735 24293 10747 24296
rect 10689 24287 10747 24293
rect 12158 24284 12164 24296
rect 12216 24284 12222 24336
rect 12802 24284 12808 24336
rect 12860 24324 12866 24336
rect 15838 24324 15844 24336
rect 12860 24296 15148 24324
rect 15799 24296 15844 24324
rect 12860 24284 12866 24296
rect 8478 24216 8484 24268
rect 8536 24256 8542 24268
rect 10870 24256 10876 24268
rect 8536 24228 10876 24256
rect 8536 24216 8542 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 10962 24216 10968 24268
rect 11020 24256 11026 24268
rect 12253 24259 12311 24265
rect 12253 24256 12265 24259
rect 11020 24228 12265 24256
rect 11020 24216 11026 24228
rect 12253 24225 12265 24228
rect 12299 24225 12311 24259
rect 15010 24256 15016 24268
rect 14971 24228 15016 24256
rect 12253 24219 12311 24225
rect 15010 24216 15016 24228
rect 15068 24216 15074 24268
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 2682 24188 2688 24200
rect 1627 24160 2688 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 2682 24148 2688 24160
rect 2740 24148 2746 24200
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 9088 24160 9321 24188
rect 9088 24148 9094 24160
rect 9309 24157 9321 24160
rect 9355 24157 9367 24191
rect 10134 24188 10140 24200
rect 10095 24160 10140 24188
rect 9309 24151 9367 24157
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 10597 24191 10655 24197
rect 10597 24157 10609 24191
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 9490 24080 9496 24132
rect 9548 24120 9554 24132
rect 10612 24120 10640 24151
rect 11238 24148 11244 24200
rect 11296 24188 11302 24200
rect 11296 24160 11341 24188
rect 11296 24148 11302 24160
rect 12342 24120 12348 24132
rect 9548 24092 10640 24120
rect 12303 24092 12348 24120
rect 9548 24080 9554 24092
rect 12342 24080 12348 24092
rect 12400 24080 12406 24132
rect 13265 24123 13323 24129
rect 13265 24089 13277 24123
rect 13311 24089 13323 24123
rect 14366 24120 14372 24132
rect 14327 24092 14372 24120
rect 13265 24083 13323 24089
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 9398 24052 9404 24064
rect 9359 24024 9404 24052
rect 9398 24012 9404 24024
rect 9456 24012 9462 24064
rect 9953 24055 10011 24061
rect 9953 24021 9965 24055
rect 9999 24052 10011 24055
rect 11146 24052 11152 24064
rect 9999 24024 11152 24052
rect 9999 24021 10011 24024
rect 9953 24015 10011 24021
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 11330 24052 11336 24064
rect 11291 24024 11336 24052
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 13280 24052 13308 24083
rect 14366 24080 14372 24092
rect 14424 24080 14430 24132
rect 14458 24080 14464 24132
rect 14516 24120 14522 24132
rect 15120 24120 15148 24296
rect 15838 24284 15844 24296
rect 15896 24284 15902 24336
rect 23382 24324 23388 24336
rect 16776 24296 23388 24324
rect 15470 24256 15476 24268
rect 15431 24228 15476 24256
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 15562 24216 15568 24268
rect 15620 24256 15626 24268
rect 15657 24259 15715 24265
rect 15657 24256 15669 24259
rect 15620 24228 15669 24256
rect 15620 24216 15626 24228
rect 15657 24225 15669 24228
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 15856 24188 15884 24284
rect 16776 24265 16804 24296
rect 23382 24284 23388 24296
rect 23440 24284 23446 24336
rect 16761 24259 16819 24265
rect 16761 24225 16773 24259
rect 16807 24225 16819 24259
rect 16942 24256 16948 24268
rect 16903 24228 16948 24256
rect 16761 24219 16819 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 19610 24256 19616 24268
rect 17512 24228 19616 24256
rect 17405 24191 17463 24197
rect 17405 24188 17417 24191
rect 15856 24160 17417 24188
rect 17405 24157 17417 24160
rect 17451 24157 17463 24191
rect 17405 24151 17463 24157
rect 17512 24120 17540 24228
rect 19610 24216 19616 24228
rect 19668 24216 19674 24268
rect 20162 24216 20168 24268
rect 20220 24256 20226 24268
rect 20530 24256 20536 24268
rect 20220 24228 20536 24256
rect 20220 24216 20226 24228
rect 20530 24216 20536 24228
rect 20588 24216 20594 24268
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24188 18475 24191
rect 18874 24188 18880 24200
rect 18463 24160 18880 24188
rect 18463 24157 18475 24160
rect 18417 24151 18475 24157
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 37458 24188 37464 24200
rect 37419 24160 37464 24188
rect 37458 24148 37464 24160
rect 37516 24148 37522 24200
rect 37737 24191 37795 24197
rect 37737 24157 37749 24191
rect 37783 24188 37795 24191
rect 37918 24188 37924 24200
rect 37783 24160 37924 24188
rect 37783 24157 37795 24160
rect 37737 24151 37795 24157
rect 37918 24148 37924 24160
rect 37976 24148 37982 24200
rect 14516 24092 14561 24120
rect 15120 24092 17540 24120
rect 14516 24080 14522 24092
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 19521 24123 19579 24129
rect 19521 24120 19533 24123
rect 18012 24092 19533 24120
rect 18012 24080 18018 24092
rect 19521 24089 19533 24092
rect 19567 24089 19579 24123
rect 19521 24083 19579 24089
rect 19610 24080 19616 24132
rect 19668 24120 19674 24132
rect 19668 24092 19713 24120
rect 19668 24080 19674 24092
rect 16298 24052 16304 24064
rect 13280 24024 16304 24052
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 18322 24012 18328 24064
rect 18380 24052 18386 24064
rect 18509 24055 18567 24061
rect 18509 24052 18521 24055
rect 18380 24024 18521 24052
rect 18380 24012 18386 24024
rect 18509 24021 18521 24024
rect 18555 24021 18567 24055
rect 22646 24052 22652 24064
rect 22607 24024 22652 24052
rect 18509 24015 18567 24021
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 10870 23808 10876 23860
rect 10928 23808 10934 23860
rect 15562 23808 15568 23860
rect 15620 23848 15626 23860
rect 22097 23851 22155 23857
rect 15620 23820 22048 23848
rect 15620 23808 15626 23820
rect 9398 23740 9404 23792
rect 9456 23780 9462 23792
rect 10413 23783 10471 23789
rect 10413 23780 10425 23783
rect 9456 23752 10425 23780
rect 9456 23740 9462 23752
rect 10413 23749 10425 23752
rect 10459 23749 10471 23783
rect 10413 23743 10471 23749
rect 10502 23740 10508 23792
rect 10560 23780 10566 23792
rect 10888 23780 10916 23808
rect 10965 23783 11023 23789
rect 10965 23780 10977 23783
rect 10560 23752 10977 23780
rect 10560 23740 10566 23752
rect 10965 23749 10977 23752
rect 11011 23749 11023 23783
rect 15102 23780 15108 23792
rect 15063 23752 15108 23780
rect 10965 23743 11023 23749
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 17129 23783 17187 23789
rect 17129 23749 17141 23783
rect 17175 23780 17187 23783
rect 17865 23783 17923 23789
rect 17865 23780 17877 23783
rect 17175 23752 17877 23780
rect 17175 23749 17187 23752
rect 17129 23743 17187 23749
rect 17865 23749 17877 23752
rect 17911 23749 17923 23783
rect 17865 23743 17923 23749
rect 5534 23672 5540 23724
rect 5592 23712 5598 23724
rect 7561 23715 7619 23721
rect 7561 23712 7573 23715
rect 5592 23684 7573 23712
rect 5592 23672 5598 23684
rect 7561 23681 7573 23684
rect 7607 23681 7619 23715
rect 7561 23675 7619 23681
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23712 8447 23715
rect 9490 23712 9496 23724
rect 8435 23684 9496 23712
rect 8435 23681 8447 23684
rect 8389 23675 8447 23681
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 13814 23712 13820 23724
rect 13775 23684 13820 23712
rect 13814 23672 13820 23684
rect 13872 23672 13878 23724
rect 13998 23712 14004 23724
rect 13959 23684 14004 23712
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 16114 23712 16120 23724
rect 16075 23684 16120 23712
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 18874 23712 18880 23724
rect 18835 23684 18880 23712
rect 17037 23675 17095 23681
rect 10321 23647 10379 23653
rect 10321 23613 10333 23647
rect 10367 23644 10379 23647
rect 11054 23644 11060 23656
rect 10367 23616 11060 23644
rect 10367 23613 10379 23616
rect 10321 23607 10379 23613
rect 11054 23604 11060 23616
rect 11112 23604 11118 23656
rect 12710 23644 12716 23656
rect 12671 23616 12716 23644
rect 12710 23604 12716 23616
rect 12768 23604 12774 23656
rect 12897 23647 12955 23653
rect 12897 23613 12909 23647
rect 12943 23644 12955 23647
rect 13906 23644 13912 23656
rect 12943 23616 13912 23644
rect 12943 23613 12955 23616
rect 12897 23607 12955 23613
rect 13906 23604 13912 23616
rect 13964 23604 13970 23656
rect 15013 23647 15071 23653
rect 15013 23613 15025 23647
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 7653 23579 7711 23585
rect 7653 23545 7665 23579
rect 7699 23576 7711 23579
rect 9398 23576 9404 23588
rect 7699 23548 9404 23576
rect 7699 23545 7711 23548
rect 7653 23539 7711 23545
rect 9398 23536 9404 23548
rect 9456 23536 9462 23588
rect 13357 23579 13415 23585
rect 13357 23545 13369 23579
rect 13403 23576 13415 23579
rect 14185 23579 14243 23585
rect 14185 23576 14197 23579
rect 13403 23548 14197 23576
rect 13403 23545 13415 23548
rect 13357 23539 13415 23545
rect 14185 23545 14197 23548
rect 14231 23576 14243 23579
rect 14366 23576 14372 23588
rect 14231 23548 14372 23576
rect 14231 23545 14243 23548
rect 14185 23539 14243 23545
rect 14366 23536 14372 23548
rect 14424 23536 14430 23588
rect 8205 23511 8263 23517
rect 8205 23477 8217 23511
rect 8251 23508 8263 23511
rect 8570 23508 8576 23520
rect 8251 23480 8576 23508
rect 8251 23477 8263 23480
rect 8205 23471 8263 23477
rect 8570 23468 8576 23480
rect 8628 23468 8634 23520
rect 13722 23468 13728 23520
rect 13780 23508 13786 23520
rect 15028 23508 15056 23607
rect 15378 23604 15384 23656
rect 15436 23644 15442 23656
rect 17052 23644 17080 23675
rect 18874 23672 18880 23684
rect 18932 23672 18938 23724
rect 22020 23721 22048 23820
rect 22097 23817 22109 23851
rect 22143 23848 22155 23851
rect 28350 23848 28356 23860
rect 22143 23820 28356 23848
rect 22143 23817 22155 23820
rect 22097 23811 22155 23817
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 30742 23848 30748 23860
rect 30703 23820 30748 23848
rect 30742 23808 30748 23820
rect 30800 23808 30806 23860
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 22646 23712 22652 23724
rect 22607 23684 22652 23712
rect 22005 23675 22063 23681
rect 22646 23672 22652 23684
rect 22704 23672 22710 23724
rect 22830 23712 22836 23724
rect 22791 23684 22836 23712
rect 22830 23672 22836 23684
rect 22888 23672 22894 23724
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23681 25835 23715
rect 25777 23675 25835 23681
rect 15436 23616 17080 23644
rect 17773 23647 17831 23653
rect 15436 23604 15442 23616
rect 17773 23613 17785 23647
rect 17819 23644 17831 23647
rect 17862 23644 17868 23656
rect 17819 23616 17868 23644
rect 17819 23613 17831 23616
rect 17773 23607 17831 23613
rect 17862 23604 17868 23616
rect 17920 23604 17926 23656
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 15565 23579 15623 23585
rect 15565 23545 15577 23579
rect 15611 23576 15623 23579
rect 17954 23576 17960 23588
rect 15611 23548 17960 23576
rect 15611 23545 15623 23548
rect 15565 23539 15623 23545
rect 17954 23536 17960 23548
rect 18012 23576 18018 23588
rect 18064 23576 18092 23607
rect 20438 23604 20444 23656
rect 20496 23644 20502 23656
rect 25792 23644 25820 23675
rect 30098 23672 30104 23724
rect 30156 23712 30162 23724
rect 30653 23715 30711 23721
rect 30653 23712 30665 23715
rect 30156 23684 30665 23712
rect 30156 23672 30162 23684
rect 30653 23681 30665 23684
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 20496 23616 25820 23644
rect 20496 23604 20502 23616
rect 18506 23576 18512 23588
rect 18012 23548 18512 23576
rect 18012 23536 18018 23548
rect 18506 23536 18512 23548
rect 18564 23536 18570 23588
rect 26206 23548 35894 23576
rect 16209 23511 16267 23517
rect 16209 23508 16221 23511
rect 13780 23480 16221 23508
rect 13780 23468 13786 23480
rect 16209 23477 16221 23480
rect 16255 23477 16267 23511
rect 16209 23471 16267 23477
rect 18414 23468 18420 23520
rect 18472 23508 18478 23520
rect 18969 23511 19027 23517
rect 18969 23508 18981 23511
rect 18472 23480 18981 23508
rect 18472 23468 18478 23480
rect 18969 23477 18981 23480
rect 19015 23477 19027 23511
rect 23014 23508 23020 23520
rect 22975 23480 23020 23508
rect 18969 23471 19027 23477
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 25593 23511 25651 23517
rect 25593 23477 25605 23511
rect 25639 23508 25651 23511
rect 26206 23508 26234 23548
rect 25639 23480 26234 23508
rect 35866 23508 35894 23548
rect 38010 23508 38016 23520
rect 35866 23480 38016 23508
rect 25639 23477 25651 23480
rect 25593 23471 25651 23477
rect 38010 23468 38016 23480
rect 38068 23468 38074 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 17494 23264 17500 23316
rect 17552 23304 17558 23316
rect 19426 23304 19432 23316
rect 17552 23276 19432 23304
rect 17552 23264 17558 23276
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 8389 23239 8447 23245
rect 8389 23205 8401 23239
rect 8435 23236 8447 23239
rect 10318 23236 10324 23248
rect 8435 23208 10324 23236
rect 8435 23205 8447 23208
rect 8389 23199 8447 23205
rect 10318 23196 10324 23208
rect 10376 23196 10382 23248
rect 12066 23236 12072 23248
rect 10704 23208 12072 23236
rect 10226 23128 10232 23180
rect 10284 23168 10290 23180
rect 10704 23168 10732 23208
rect 12066 23196 12072 23208
rect 12124 23196 12130 23248
rect 16025 23239 16083 23245
rect 16025 23205 16037 23239
rect 16071 23236 16083 23239
rect 16574 23236 16580 23248
rect 16071 23208 16580 23236
rect 16071 23205 16083 23208
rect 16025 23199 16083 23205
rect 16574 23196 16580 23208
rect 16632 23196 16638 23248
rect 24946 23236 24952 23248
rect 18248 23208 24952 23236
rect 18248 23177 18276 23208
rect 24946 23196 24952 23208
rect 25004 23196 25010 23248
rect 10284 23140 10732 23168
rect 10781 23171 10839 23177
rect 10284 23128 10290 23140
rect 10781 23137 10793 23171
rect 10827 23168 10839 23171
rect 12253 23171 12311 23177
rect 12253 23168 12265 23171
rect 10827 23140 12265 23168
rect 10827 23137 10839 23140
rect 10781 23131 10839 23137
rect 12253 23137 12265 23140
rect 12299 23137 12311 23171
rect 12253 23131 12311 23137
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23137 18291 23171
rect 18506 23168 18512 23180
rect 18467 23140 18512 23168
rect 18233 23131 18291 23137
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 20622 23168 20628 23180
rect 20180 23140 20628 23168
rect 1946 23060 1952 23112
rect 2004 23100 2010 23112
rect 7745 23103 7803 23109
rect 7745 23100 7757 23103
rect 2004 23072 7757 23100
rect 2004 23060 2010 23072
rect 7745 23069 7757 23072
rect 7791 23069 7803 23103
rect 8570 23100 8576 23112
rect 8531 23072 8576 23100
rect 7745 23063 7803 23069
rect 8570 23060 8576 23072
rect 8628 23060 8634 23112
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9306 23100 9312 23112
rect 9171 23072 9312 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 10686 23100 10692 23112
rect 10647 23072 10692 23100
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 12069 23103 12127 23109
rect 12069 23069 12081 23103
rect 12115 23100 12127 23103
rect 12710 23100 12716 23112
rect 12115 23072 12716 23100
rect 12115 23069 12127 23072
rect 12069 23063 12127 23069
rect 7837 23035 7895 23041
rect 7837 23001 7849 23035
rect 7883 23032 7895 23035
rect 12084 23032 12112 23063
rect 12710 23060 12716 23072
rect 12768 23060 12774 23112
rect 20180 23109 20208 23140
rect 20622 23128 20628 23140
rect 20680 23168 20686 23180
rect 22738 23168 22744 23180
rect 20680 23140 22744 23168
rect 20680 23128 20686 23140
rect 22738 23128 22744 23140
rect 22796 23128 22802 23180
rect 20165 23103 20223 23109
rect 20165 23069 20177 23103
rect 20211 23069 20223 23103
rect 20165 23063 20223 23069
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21085 23103 21143 23109
rect 21085 23100 21097 23103
rect 20864 23072 21097 23100
rect 20864 23060 20870 23072
rect 21085 23069 21097 23072
rect 21131 23069 21143 23103
rect 21634 23100 21640 23112
rect 21595 23072 21640 23100
rect 21085 23063 21143 23069
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 7883 23004 12112 23032
rect 7883 23001 7895 23004
rect 7837 22995 7895 23001
rect 12526 22992 12532 23044
rect 12584 23032 12590 23044
rect 15841 23035 15899 23041
rect 15841 23032 15853 23035
rect 12584 23004 15853 23032
rect 12584 22992 12590 23004
rect 15841 23001 15853 23004
rect 15887 23001 15899 23035
rect 15841 22995 15899 23001
rect 18322 22992 18328 23044
rect 18380 23032 18386 23044
rect 18380 23004 18425 23032
rect 18380 22992 18386 23004
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 10778 22964 10784 22976
rect 9263 22936 10784 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 12710 22964 12716 22976
rect 12671 22936 12716 22964
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 13170 22964 13176 22976
rect 13131 22936 13176 22964
rect 13170 22924 13176 22936
rect 13228 22924 13234 22976
rect 14734 22964 14740 22976
rect 14695 22936 14740 22964
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 20254 22964 20260 22976
rect 20215 22936 20260 22964
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 20901 22967 20959 22973
rect 20901 22933 20913 22967
rect 20947 22964 20959 22967
rect 21450 22964 21456 22976
rect 20947 22936 21456 22964
rect 20947 22933 20959 22936
rect 20901 22927 20959 22933
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 21729 22967 21787 22973
rect 21729 22933 21741 22967
rect 21775 22964 21787 22967
rect 23474 22964 23480 22976
rect 21775 22936 23480 22964
rect 21775 22933 21787 22936
rect 21729 22927 21787 22933
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 2314 22760 2320 22772
rect 2275 22732 2320 22760
rect 2314 22720 2320 22732
rect 2372 22720 2378 22772
rect 8389 22763 8447 22769
rect 8389 22729 8401 22763
rect 8435 22760 8447 22763
rect 10226 22760 10232 22772
rect 8435 22732 10232 22760
rect 8435 22729 8447 22732
rect 8389 22723 8447 22729
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 10686 22760 10692 22772
rect 10336 22732 10692 22760
rect 4062 22652 4068 22704
rect 4120 22692 4126 22704
rect 4120 22664 8340 22692
rect 4120 22652 4126 22664
rect 1670 22624 1676 22636
rect 1631 22596 1676 22624
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 2498 22624 2504 22636
rect 2459 22596 2504 22624
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 7190 22624 7196 22636
rect 7151 22596 7196 22624
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 8312 22633 8340 22664
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22593 8355 22627
rect 8297 22587 8355 22593
rect 9125 22627 9183 22633
rect 9125 22593 9137 22627
rect 9171 22624 9183 22627
rect 9306 22624 9312 22636
rect 9171 22596 9312 22624
rect 9171 22593 9183 22596
rect 9125 22587 9183 22593
rect 9306 22584 9312 22596
rect 9364 22584 9370 22636
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 10336 22624 10364 22732
rect 10686 22720 10692 22732
rect 10744 22720 10750 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 11422 22760 11428 22772
rect 11112 22732 11428 22760
rect 11112 22720 11118 22732
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 14369 22763 14427 22769
rect 14369 22729 14381 22763
rect 14415 22760 14427 22763
rect 15102 22760 15108 22772
rect 14415 22732 15108 22760
rect 14415 22729 14427 22732
rect 14369 22723 14427 22729
rect 15102 22720 15108 22732
rect 15160 22720 15166 22772
rect 15654 22720 15660 22772
rect 15712 22760 15718 22772
rect 20257 22763 20315 22769
rect 15712 22732 16344 22760
rect 15712 22720 15718 22732
rect 10597 22695 10655 22701
rect 10597 22661 10609 22695
rect 10643 22692 10655 22695
rect 11330 22692 11336 22704
rect 10643 22664 11336 22692
rect 10643 22661 10655 22664
rect 10597 22655 10655 22661
rect 11330 22652 11336 22664
rect 11388 22652 11394 22704
rect 15746 22692 15752 22704
rect 13648 22664 14964 22692
rect 15707 22664 15752 22692
rect 13648 22636 13676 22664
rect 11882 22624 11888 22636
rect 9815 22596 10364 22624
rect 11164 22596 11888 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 9398 22516 9404 22568
rect 9456 22556 9462 22568
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 9456 22528 10517 22556
rect 9456 22516 9462 22528
rect 10505 22525 10517 22528
rect 10551 22556 10563 22559
rect 11164 22556 11192 22596
rect 11882 22584 11888 22596
rect 11940 22584 11946 22636
rect 12069 22627 12127 22633
rect 12069 22593 12081 22627
rect 12115 22624 12127 22627
rect 13630 22624 13636 22636
rect 12115 22596 12434 22624
rect 13543 22596 13636 22624
rect 12115 22593 12127 22596
rect 12069 22587 12127 22593
rect 10551 22528 11192 22556
rect 10551 22525 10563 22528
rect 10505 22519 10563 22525
rect 12158 22516 12164 22568
rect 12216 22556 12222 22568
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 12216 22528 12265 22556
rect 12216 22516 12222 22528
rect 12253 22525 12265 22528
rect 12299 22525 12311 22559
rect 12406 22556 12434 22596
rect 13630 22584 13636 22596
rect 13688 22584 13694 22636
rect 14277 22627 14335 22633
rect 14277 22593 14289 22627
rect 14323 22624 14335 22627
rect 14642 22624 14648 22636
rect 14323 22596 14648 22624
rect 14323 22593 14335 22596
rect 14277 22587 14335 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 14936 22633 14964 22664
rect 15746 22652 15752 22664
rect 15804 22652 15810 22704
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22593 14979 22627
rect 14921 22587 14979 22593
rect 13722 22556 13728 22568
rect 12406 22528 13728 22556
rect 12253 22519 12311 22525
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 15657 22559 15715 22565
rect 15657 22525 15669 22559
rect 15703 22556 15715 22559
rect 15838 22556 15844 22568
rect 15703 22528 15844 22556
rect 15703 22525 15715 22528
rect 15657 22519 15715 22525
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 15933 22559 15991 22565
rect 15933 22525 15945 22559
rect 15979 22525 15991 22559
rect 16316 22556 16344 22732
rect 20257 22729 20269 22763
rect 20303 22760 20315 22763
rect 23014 22760 23020 22772
rect 20303 22732 23020 22760
rect 20303 22729 20315 22732
rect 20257 22723 20315 22729
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 29178 22760 29184 22772
rect 29139 22732 29184 22760
rect 29178 22720 29184 22732
rect 29236 22720 29242 22772
rect 17126 22692 17132 22704
rect 17087 22664 17132 22692
rect 17126 22652 17132 22664
rect 17184 22652 17190 22704
rect 17681 22695 17739 22701
rect 17681 22661 17693 22695
rect 17727 22692 17739 22695
rect 19334 22692 19340 22704
rect 17727 22664 19340 22692
rect 17727 22661 17739 22664
rect 17681 22655 17739 22661
rect 19334 22652 19340 22664
rect 19392 22692 19398 22704
rect 20530 22692 20536 22704
rect 19392 22664 20536 22692
rect 19392 22652 19398 22664
rect 20530 22652 20536 22664
rect 20588 22652 20594 22704
rect 23474 22692 23480 22704
rect 23435 22664 23480 22692
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 25038 22692 25044 22704
rect 24999 22664 25044 22692
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 26510 22652 26516 22704
rect 26568 22692 26574 22704
rect 26568 22664 35894 22692
rect 26568 22652 26574 22664
rect 19797 22627 19855 22633
rect 19797 22593 19809 22627
rect 19843 22624 19855 22627
rect 20254 22624 20260 22636
rect 19843 22596 20260 22624
rect 19843 22593 19855 22596
rect 19797 22587 19855 22593
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 20622 22584 20628 22636
rect 20680 22624 20686 22636
rect 20901 22627 20959 22633
rect 20901 22624 20913 22627
rect 20680 22596 20913 22624
rect 20680 22584 20686 22596
rect 20901 22593 20913 22596
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 22189 22627 22247 22633
rect 22189 22624 22201 22627
rect 21508 22596 22201 22624
rect 21508 22584 21514 22596
rect 22189 22593 22201 22596
rect 22235 22593 22247 22627
rect 29086 22624 29092 22636
rect 29047 22596 29092 22624
rect 22189 22587 22247 22593
rect 29086 22584 29092 22596
rect 29144 22584 29150 22636
rect 35866 22624 35894 22664
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 35866 22596 38025 22624
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 17037 22559 17095 22565
rect 17037 22556 17049 22559
rect 16316 22528 17049 22556
rect 15933 22519 15991 22525
rect 17037 22525 17049 22528
rect 17083 22525 17095 22559
rect 17037 22519 17095 22525
rect 19613 22559 19671 22565
rect 19613 22525 19625 22559
rect 19659 22556 19671 22559
rect 20346 22556 20352 22568
rect 19659 22528 20352 22556
rect 19659 22525 19671 22528
rect 19613 22519 19671 22525
rect 2498 22448 2504 22500
rect 2556 22488 2562 22500
rect 9122 22488 9128 22500
rect 2556 22460 9128 22488
rect 2556 22448 2562 22460
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 9217 22491 9275 22497
rect 9217 22457 9229 22491
rect 9263 22488 9275 22491
rect 11057 22491 11115 22497
rect 9263 22460 10548 22488
rect 9263 22457 9275 22460
rect 9217 22451 9275 22457
rect 10520 22432 10548 22460
rect 11057 22457 11069 22491
rect 11103 22488 11115 22491
rect 11238 22488 11244 22500
rect 11103 22460 11244 22488
rect 11103 22457 11115 22460
rect 11057 22451 11115 22457
rect 11238 22448 11244 22460
rect 11296 22448 11302 22500
rect 11422 22448 11428 22500
rect 11480 22488 11486 22500
rect 12437 22491 12495 22497
rect 12437 22488 12449 22491
rect 11480 22460 12449 22488
rect 11480 22448 11486 22460
rect 12437 22457 12449 22460
rect 12483 22457 12495 22491
rect 15948 22488 15976 22519
rect 20346 22516 20352 22528
rect 20404 22516 20410 22568
rect 23385 22559 23443 22565
rect 23385 22525 23397 22559
rect 23431 22556 23443 22559
rect 24026 22556 24032 22568
rect 23431 22528 24032 22556
rect 23431 22525 23443 22528
rect 23385 22519 23443 22525
rect 24026 22516 24032 22528
rect 24084 22516 24090 22568
rect 24302 22556 24308 22568
rect 24263 22528 24308 22556
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 24946 22556 24952 22568
rect 24907 22528 24952 22556
rect 24946 22516 24952 22528
rect 25004 22516 25010 22568
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22525 25283 22559
rect 25225 22519 25283 22525
rect 17402 22488 17408 22500
rect 12437 22451 12495 22457
rect 13556 22460 17408 22488
rect 1762 22420 1768 22432
rect 1723 22392 1768 22420
rect 1762 22380 1768 22392
rect 1820 22380 1826 22432
rect 7009 22423 7067 22429
rect 7009 22389 7021 22423
rect 7055 22420 7067 22423
rect 7282 22420 7288 22432
rect 7055 22392 7288 22420
rect 7055 22389 7067 22392
rect 7009 22383 7067 22389
rect 7282 22380 7288 22392
rect 7340 22380 7346 22432
rect 9766 22380 9772 22432
rect 9824 22420 9830 22432
rect 9861 22423 9919 22429
rect 9861 22420 9873 22423
rect 9824 22392 9873 22420
rect 9824 22380 9830 22392
rect 9861 22389 9873 22392
rect 9907 22389 9919 22423
rect 9861 22383 9919 22389
rect 10502 22380 10508 22432
rect 10560 22380 10566 22432
rect 11256 22420 11284 22448
rect 13556 22420 13584 22460
rect 17402 22448 17408 22460
rect 17460 22448 17466 22500
rect 25240 22488 25268 22519
rect 38194 22488 38200 22500
rect 19306 22460 25268 22488
rect 38155 22460 38200 22488
rect 13722 22420 13728 22432
rect 11256 22392 13584 22420
rect 13683 22392 13728 22420
rect 13722 22380 13728 22392
rect 13780 22380 13786 22432
rect 15010 22420 15016 22432
rect 14971 22392 15016 22420
rect 15010 22380 15016 22392
rect 15068 22380 15074 22432
rect 16850 22380 16856 22432
rect 16908 22420 16914 22432
rect 18322 22420 18328 22432
rect 16908 22392 18328 22420
rect 16908 22380 16914 22392
rect 18322 22380 18328 22392
rect 18380 22420 18386 22432
rect 19306 22420 19334 22460
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 20990 22420 20996 22432
rect 18380 22392 19334 22420
rect 20951 22392 20996 22420
rect 18380 22380 18386 22392
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 22738 22420 22744 22432
rect 22051 22392 22744 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 22738 22380 22744 22392
rect 22796 22380 22802 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1762 22176 1768 22228
rect 1820 22216 1826 22228
rect 1820 22188 12434 22216
rect 1820 22176 1826 22188
rect 12406 22148 12434 22188
rect 12710 22176 12716 22228
rect 12768 22216 12774 22228
rect 13173 22219 13231 22225
rect 13173 22216 13185 22219
rect 12768 22188 13185 22216
rect 12768 22176 12774 22188
rect 13173 22185 13185 22188
rect 13219 22216 13231 22219
rect 13262 22216 13268 22228
rect 13219 22188 13268 22216
rect 13219 22185 13231 22188
rect 13173 22179 13231 22185
rect 13262 22176 13268 22188
rect 13320 22176 13326 22228
rect 17678 22216 17684 22228
rect 13372 22188 17684 22216
rect 13372 22148 13400 22188
rect 17678 22176 17684 22188
rect 17736 22176 17742 22228
rect 12406 22120 13400 22148
rect 17402 22108 17408 22160
rect 17460 22148 17466 22160
rect 17460 22120 18552 22148
rect 17460 22108 17466 22120
rect 9950 22040 9956 22092
rect 10008 22080 10014 22092
rect 10008 22052 12204 22080
rect 10008 22040 10014 22052
rect 1946 22012 1952 22024
rect 1907 21984 1952 22012
rect 1946 21972 1952 21984
rect 2004 21972 2010 22024
rect 7282 22012 7288 22024
rect 7243 21984 7288 22012
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 12176 22021 12204 22052
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12618 22080 12624 22092
rect 12308 22052 12624 22080
rect 12308 22040 12314 22052
rect 12618 22040 12624 22052
rect 12676 22040 12682 22092
rect 12805 22083 12863 22089
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 13170 22080 13176 22092
rect 12851 22052 13176 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 14734 22080 14740 22092
rect 14695 22052 14740 22080
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 14918 22040 14924 22092
rect 14976 22080 14982 22092
rect 15749 22083 15807 22089
rect 15749 22080 15761 22083
rect 14976 22052 15761 22080
rect 14976 22040 14982 22052
rect 15749 22049 15761 22052
rect 15795 22080 15807 22083
rect 16298 22080 16304 22092
rect 15795 22052 16304 22080
rect 15795 22049 15807 22052
rect 15749 22043 15807 22049
rect 16298 22040 16304 22052
rect 16356 22040 16362 22092
rect 18230 22080 18236 22092
rect 18191 22052 18236 22080
rect 18230 22040 18236 22052
rect 18288 22040 18294 22092
rect 18524 22089 18552 22120
rect 18509 22083 18567 22089
rect 18509 22049 18521 22083
rect 18555 22049 18567 22083
rect 18509 22043 18567 22049
rect 19521 22083 19579 22089
rect 19521 22049 19533 22083
rect 19567 22080 19579 22083
rect 20070 22080 20076 22092
rect 19567 22052 20076 22080
rect 19567 22049 19579 22052
rect 19521 22043 19579 22049
rect 20070 22040 20076 22052
rect 20128 22040 20134 22092
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 21361 22083 21419 22089
rect 21361 22080 21373 22083
rect 20220 22052 21373 22080
rect 20220 22040 20226 22052
rect 21361 22049 21373 22052
rect 21407 22049 21419 22083
rect 23290 22080 23296 22092
rect 23203 22052 23296 22080
rect 21361 22043 21419 22049
rect 23290 22040 23296 22052
rect 23348 22080 23354 22092
rect 27982 22080 27988 22092
rect 23348 22052 27988 22080
rect 23348 22040 23354 22052
rect 27982 22040 27988 22052
rect 28040 22040 28046 22092
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12526 22012 12532 22024
rect 12207 21984 12532 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 12986 22012 12992 22024
rect 12947 21984 12992 22012
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 22012 23995 22015
rect 24578 22012 24584 22024
rect 23983 21984 24584 22012
rect 23983 21981 23995 21984
rect 23937 21975 23995 21981
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 31481 22015 31539 22021
rect 31481 21981 31493 22015
rect 31527 22012 31539 22015
rect 38102 22012 38108 22024
rect 31527 21984 38108 22012
rect 31527 21981 31539 21984
rect 31481 21975 31539 21981
rect 38102 21972 38108 21984
rect 38160 21972 38166 22024
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 7190 21904 7196 21956
rect 7248 21944 7254 21956
rect 10689 21947 10747 21953
rect 7248 21916 7420 21944
rect 7248 21904 7254 21916
rect 7392 21888 7420 21916
rect 10689 21913 10701 21947
rect 10735 21913 10747 21947
rect 10689 21907 10747 21913
rect 1578 21836 1584 21888
rect 1636 21876 1642 21888
rect 1765 21879 1823 21885
rect 1765 21876 1777 21879
rect 1636 21848 1777 21876
rect 1636 21836 1642 21848
rect 1765 21845 1777 21848
rect 1811 21845 1823 21879
rect 1765 21839 1823 21845
rect 7101 21879 7159 21885
rect 7101 21845 7113 21879
rect 7147 21876 7159 21879
rect 7282 21876 7288 21888
rect 7147 21848 7288 21876
rect 7147 21845 7159 21848
rect 7101 21839 7159 21845
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 10594 21876 10600 21888
rect 7432 21848 10600 21876
rect 7432 21836 7438 21848
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 10704 21876 10732 21907
rect 10778 21904 10784 21956
rect 10836 21944 10842 21956
rect 11698 21944 11704 21956
rect 10836 21916 10881 21944
rect 11659 21916 11704 21944
rect 10836 21904 10842 21916
rect 11698 21904 11704 21916
rect 11756 21904 11762 21956
rect 14826 21944 14832 21956
rect 14787 21916 14832 21944
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 16022 21904 16028 21956
rect 16080 21944 16086 21956
rect 16301 21947 16359 21953
rect 16301 21944 16313 21947
rect 16080 21916 16313 21944
rect 16080 21904 16086 21916
rect 16301 21913 16313 21916
rect 16347 21913 16359 21947
rect 16301 21907 16359 21913
rect 16393 21947 16451 21953
rect 16393 21913 16405 21947
rect 16439 21913 16451 21947
rect 16393 21907 16451 21913
rect 12250 21876 12256 21888
rect 10704 21848 12256 21876
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 12342 21836 12348 21888
rect 12400 21876 12406 21888
rect 16408 21876 16436 21907
rect 16666 21904 16672 21956
rect 16724 21944 16730 21956
rect 16945 21947 17003 21953
rect 16945 21944 16957 21947
rect 16724 21916 16957 21944
rect 16724 21904 16730 21916
rect 16945 21913 16957 21916
rect 16991 21944 17003 21947
rect 17770 21944 17776 21956
rect 16991 21916 17776 21944
rect 16991 21913 17003 21916
rect 16945 21907 17003 21913
rect 17770 21904 17776 21916
rect 17828 21904 17834 21956
rect 18325 21947 18383 21953
rect 18325 21913 18337 21947
rect 18371 21944 18383 21947
rect 18414 21944 18420 21956
rect 18371 21916 18420 21944
rect 18371 21913 18383 21916
rect 18325 21907 18383 21913
rect 18414 21904 18420 21916
rect 18472 21904 18478 21956
rect 19606 21947 19664 21953
rect 19606 21913 19618 21947
rect 19652 21913 19664 21947
rect 21082 21944 21088 21956
rect 21043 21916 21088 21944
rect 19606 21907 19664 21913
rect 12400 21848 16436 21876
rect 12400 21836 12406 21848
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19628 21876 19656 21907
rect 21082 21904 21088 21916
rect 21140 21904 21146 21956
rect 21174 21904 21180 21956
rect 21232 21944 21238 21956
rect 22646 21944 22652 21956
rect 21232 21916 21277 21944
rect 22607 21916 22652 21944
rect 21232 21904 21238 21916
rect 22646 21904 22652 21916
rect 22704 21904 22710 21956
rect 22738 21904 22744 21956
rect 22796 21944 22802 21956
rect 22796 21916 22841 21944
rect 22796 21904 22802 21916
rect 23750 21876 23756 21888
rect 19484 21848 19656 21876
rect 23711 21848 23756 21876
rect 19484 21836 19490 21848
rect 23750 21836 23756 21848
rect 23808 21836 23814 21888
rect 27522 21836 27528 21888
rect 27580 21876 27586 21888
rect 31573 21879 31631 21885
rect 31573 21876 31585 21879
rect 27580 21848 31585 21876
rect 27580 21836 27586 21848
rect 31573 21845 31585 21848
rect 31619 21845 31631 21879
rect 31573 21839 31631 21845
rect 34698 21836 34704 21888
rect 34756 21876 34762 21888
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 34756 21848 38117 21876
rect 34756 21836 34762 21848
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 8386 21632 8392 21684
rect 8444 21672 8450 21684
rect 10962 21672 10968 21684
rect 8444 21644 10968 21672
rect 8444 21632 8450 21644
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 11149 21675 11207 21681
rect 11149 21672 11161 21675
rect 11112 21644 11161 21672
rect 11112 21632 11118 21644
rect 11149 21641 11161 21644
rect 11195 21641 11207 21675
rect 11698 21672 11704 21684
rect 11149 21635 11207 21641
rect 11256 21644 11704 21672
rect 8846 21564 8852 21616
rect 8904 21604 8910 21616
rect 11256 21604 11284 21644
rect 11698 21632 11704 21644
rect 11756 21672 11762 21684
rect 17494 21672 17500 21684
rect 11756 21644 16252 21672
rect 17455 21644 17500 21672
rect 11756 21632 11762 21644
rect 12345 21607 12403 21613
rect 12345 21604 12357 21607
rect 8904 21576 11284 21604
rect 11440 21576 12357 21604
rect 8904 21564 8910 21576
rect 1578 21536 1584 21548
rect 1539 21508 1584 21536
rect 1578 21496 1584 21508
rect 1636 21496 1642 21548
rect 7193 21539 7251 21545
rect 7193 21505 7205 21539
rect 7239 21536 7251 21539
rect 7374 21536 7380 21548
rect 7239 21508 7380 21536
rect 7239 21505 7251 21508
rect 7193 21499 7251 21505
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 9122 21536 9128 21548
rect 9083 21508 9128 21536
rect 8481 21499 8539 21505
rect 8496 21400 8524 21499
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 10376 21508 10701 21536
rect 10376 21496 10382 21508
rect 10689 21505 10701 21508
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 9217 21471 9275 21477
rect 9217 21437 9229 21471
rect 9263 21468 9275 21471
rect 10505 21471 10563 21477
rect 10505 21468 10517 21471
rect 9263 21440 10517 21468
rect 9263 21437 9275 21440
rect 9217 21431 9275 21437
rect 10505 21437 10517 21440
rect 10551 21468 10563 21471
rect 10551 21440 10732 21468
rect 10551 21437 10563 21440
rect 10505 21431 10563 21437
rect 9858 21400 9864 21412
rect 8496 21372 9864 21400
rect 9858 21360 9864 21372
rect 9916 21360 9922 21412
rect 1762 21332 1768 21344
rect 1723 21304 1768 21332
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7285 21335 7343 21341
rect 7285 21332 7297 21335
rect 6972 21304 7297 21332
rect 6972 21292 6978 21304
rect 7285 21301 7297 21304
rect 7331 21301 7343 21335
rect 7285 21295 7343 21301
rect 8573 21335 8631 21341
rect 8573 21301 8585 21335
rect 8619 21332 8631 21335
rect 8662 21332 8668 21344
rect 8619 21304 8668 21332
rect 8619 21301 8631 21304
rect 8573 21295 8631 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 10704 21332 10732 21440
rect 11146 21428 11152 21480
rect 11204 21468 11210 21480
rect 11440 21468 11468 21576
rect 12345 21573 12357 21576
rect 12391 21573 12403 21607
rect 12345 21567 12403 21573
rect 13262 21564 13268 21616
rect 13320 21604 13326 21616
rect 13725 21607 13783 21613
rect 13725 21604 13737 21607
rect 13320 21576 13737 21604
rect 13320 21564 13326 21576
rect 13725 21573 13737 21576
rect 13771 21573 13783 21607
rect 13725 21567 13783 21573
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 13872 21576 13917 21604
rect 13872 21564 13878 21576
rect 15194 21564 15200 21616
rect 15252 21604 15258 21616
rect 16224 21613 16252 21644
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 17862 21632 17868 21684
rect 17920 21672 17926 21684
rect 17920 21644 20208 21672
rect 17920 21632 17926 21644
rect 15289 21607 15347 21613
rect 15289 21604 15301 21607
rect 15252 21576 15301 21604
rect 15252 21564 15258 21576
rect 15289 21573 15301 21576
rect 15335 21573 15347 21607
rect 15289 21567 15347 21573
rect 16209 21607 16267 21613
rect 16209 21573 16221 21607
rect 16255 21573 16267 21607
rect 16209 21567 16267 21573
rect 19334 21564 19340 21616
rect 19392 21604 19398 21616
rect 20073 21607 20131 21613
rect 20073 21604 20085 21607
rect 19392 21576 20085 21604
rect 19392 21564 19398 21576
rect 20073 21573 20085 21576
rect 20119 21573 20131 21607
rect 20180 21604 20208 21644
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 21140 21644 22017 21672
rect 21140 21632 21146 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22646 21672 22652 21684
rect 22607 21644 22652 21672
rect 22005 21635 22063 21641
rect 22646 21632 22652 21644
rect 22704 21632 22710 21684
rect 21177 21607 21235 21613
rect 21177 21604 21189 21607
rect 20180 21576 21189 21604
rect 20073 21567 20131 21573
rect 21177 21573 21189 21576
rect 21223 21573 21235 21607
rect 27522 21604 27528 21616
rect 21177 21567 21235 21573
rect 22066 21576 27200 21604
rect 27483 21576 27528 21604
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 16845 21537 16903 21543
rect 16356 21534 16804 21536
rect 16845 21534 16857 21537
rect 16356 21508 16857 21534
rect 16356 21496 16362 21508
rect 16776 21506 16857 21508
rect 16845 21503 16857 21506
rect 16891 21503 16903 21537
rect 16845 21497 16903 21503
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 18598 21536 18604 21548
rect 18559 21508 18604 21536
rect 17681 21499 17739 21505
rect 11204 21440 11468 21468
rect 12253 21471 12311 21477
rect 11204 21428 11210 21440
rect 12253 21437 12265 21471
rect 12299 21468 12311 21471
rect 12342 21468 12348 21480
rect 12299 21440 12348 21468
rect 12299 21437 12311 21440
rect 12253 21431 12311 21437
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21437 12587 21471
rect 12529 21431 12587 21437
rect 11054 21360 11060 21412
rect 11112 21400 11118 21412
rect 12544 21400 12572 21431
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 13814 21468 13820 21480
rect 12768 21440 13820 21468
rect 12768 21428 12774 21440
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 15194 21468 15200 21480
rect 15155 21440 15200 21468
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 11112 21372 12572 21400
rect 14277 21403 14335 21409
rect 11112 21360 11118 21372
rect 14277 21369 14289 21403
rect 14323 21369 14335 21403
rect 14277 21363 14335 21369
rect 10778 21332 10784 21344
rect 10704 21304 10784 21332
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 14292 21332 14320 21363
rect 14366 21360 14372 21412
rect 14424 21400 14430 21412
rect 17696 21400 17724 21499
rect 18598 21496 18604 21508
rect 18656 21536 18662 21548
rect 19702 21536 19708 21548
rect 18656 21508 19708 21536
rect 18656 21496 18662 21508
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 21082 21536 21088 21548
rect 20956 21508 21088 21536
rect 20956 21496 20962 21508
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 22066 21536 22094 21576
rect 21324 21508 22094 21536
rect 21324 21496 21330 21508
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23072 21508 23397 21536
rect 23072 21496 23078 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 23750 21536 23756 21548
rect 23615 21508 23756 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 23842 21496 23848 21548
rect 23900 21536 23906 21548
rect 24581 21539 24639 21545
rect 24581 21536 24593 21539
rect 23900 21508 24593 21536
rect 23900 21496 23906 21508
rect 24581 21505 24593 21508
rect 24627 21505 24639 21539
rect 25498 21536 25504 21548
rect 25459 21508 25504 21536
rect 24581 21499 24639 21505
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 19245 21471 19303 21477
rect 19245 21437 19257 21471
rect 19291 21468 19303 21471
rect 19981 21471 20039 21477
rect 19981 21468 19993 21471
rect 19291 21440 19993 21468
rect 19291 21437 19303 21440
rect 19245 21431 19303 21437
rect 19981 21437 19993 21440
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21468 20315 21471
rect 27062 21468 27068 21480
rect 20303 21440 27068 21468
rect 20303 21437 20315 21440
rect 20257 21431 20315 21437
rect 14424 21372 17724 21400
rect 14424 21360 14430 21372
rect 17770 21360 17776 21412
rect 17828 21400 17834 21412
rect 20272 21400 20300 21431
rect 27062 21428 27068 21440
rect 27120 21428 27126 21480
rect 27172 21468 27200 21576
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 27614 21564 27620 21616
rect 27672 21604 27678 21616
rect 27672 21576 27717 21604
rect 27672 21564 27678 21576
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 37366 21536 37372 21548
rect 31251 21508 37372 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 37366 21496 37372 21508
rect 37424 21496 37430 21548
rect 28537 21471 28595 21477
rect 28537 21468 28549 21471
rect 27172 21440 28549 21468
rect 28537 21437 28549 21440
rect 28583 21468 28595 21471
rect 30834 21468 30840 21480
rect 28583 21440 30840 21468
rect 28583 21437 28595 21440
rect 28537 21431 28595 21437
rect 30834 21428 30840 21440
rect 30892 21428 30898 21480
rect 17828 21372 20300 21400
rect 17828 21360 17834 21372
rect 20714 21360 20720 21412
rect 20772 21400 20778 21412
rect 25593 21403 25651 21409
rect 25593 21400 25605 21403
rect 20772 21372 25605 21400
rect 20772 21360 20778 21372
rect 25593 21369 25605 21372
rect 25639 21369 25651 21403
rect 25593 21363 25651 21369
rect 15562 21332 15568 21344
rect 14292 21304 15568 21332
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 16574 21332 16580 21344
rect 16080 21304 16580 21332
rect 16080 21292 16086 21304
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 16942 21332 16948 21344
rect 16903 21304 16948 21332
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 18693 21335 18751 21341
rect 18693 21301 18705 21335
rect 18739 21332 18751 21335
rect 19610 21332 19616 21344
rect 18739 21304 19616 21332
rect 18739 21301 18751 21304
rect 18693 21295 18751 21301
rect 19610 21292 19616 21304
rect 19668 21292 19674 21344
rect 19702 21292 19708 21344
rect 19760 21332 19766 21344
rect 20806 21332 20812 21344
rect 19760 21304 20812 21332
rect 19760 21292 19766 21304
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 24026 21332 24032 21344
rect 23987 21304 24032 21332
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24670 21332 24676 21344
rect 24631 21304 24676 21332
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 29454 21292 29460 21344
rect 29512 21332 29518 21344
rect 31297 21335 31355 21341
rect 31297 21332 31309 21335
rect 29512 21304 31309 21332
rect 29512 21292 29518 21304
rect 31297 21301 31309 21304
rect 31343 21301 31355 21335
rect 31297 21295 31355 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1581 21131 1639 21137
rect 1581 21097 1593 21131
rect 1627 21128 1639 21131
rect 8294 21128 8300 21140
rect 1627 21100 8300 21128
rect 1627 21097 1639 21100
rect 1581 21091 1639 21097
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 8478 21128 8484 21140
rect 8439 21100 8484 21128
rect 8478 21088 8484 21100
rect 8536 21088 8542 21140
rect 8938 21088 8944 21140
rect 8996 21128 9002 21140
rect 11146 21128 11152 21140
rect 8996 21100 11152 21128
rect 8996 21088 9002 21100
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 12406 21100 17540 21128
rect 6641 21063 6699 21069
rect 6641 21029 6653 21063
rect 6687 21060 6699 21063
rect 11054 21060 11060 21072
rect 6687 21032 9444 21060
rect 6687 21029 6699 21032
rect 6641 21023 6699 21029
rect 5166 20952 5172 21004
rect 5224 20992 5230 21004
rect 9416 20992 9444 21032
rect 9600 21032 11060 21060
rect 9600 20992 9628 21032
rect 11054 21020 11060 21032
rect 11112 21060 11118 21072
rect 12406 21060 12434 21100
rect 11112 21032 12434 21060
rect 13633 21063 13691 21069
rect 11112 21020 11118 21032
rect 13633 21029 13645 21063
rect 13679 21060 13691 21063
rect 16022 21060 16028 21072
rect 13679 21032 16028 21060
rect 13679 21029 13691 21032
rect 13633 21023 13691 21029
rect 16022 21020 16028 21032
rect 16080 21020 16086 21072
rect 16114 21020 16120 21072
rect 16172 21060 16178 21072
rect 17034 21060 17040 21072
rect 16172 21032 17040 21060
rect 16172 21020 16178 21032
rect 17034 21020 17040 21032
rect 17092 21020 17098 21072
rect 5224 20964 7512 20992
rect 9416 20964 9628 20992
rect 5224 20952 5230 20964
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 7374 20924 7380 20936
rect 7335 20896 7380 20924
rect 7374 20884 7380 20896
rect 7432 20884 7438 20936
rect 5258 20816 5264 20868
rect 5316 20856 5322 20868
rect 6089 20859 6147 20865
rect 6089 20856 6101 20859
rect 5316 20828 6101 20856
rect 5316 20816 5322 20828
rect 6089 20825 6101 20828
rect 6135 20825 6147 20859
rect 6089 20819 6147 20825
rect 6181 20859 6239 20865
rect 6181 20825 6193 20859
rect 6227 20825 6239 20859
rect 6181 20819 6239 20825
rect 6196 20788 6224 20819
rect 7193 20791 7251 20797
rect 7193 20788 7205 20791
rect 6196 20760 7205 20788
rect 7193 20757 7205 20760
rect 7239 20757 7251 20791
rect 7484 20788 7512 20964
rect 12342 20952 12348 21004
rect 12400 20992 12406 21004
rect 12400 20964 12445 20992
rect 12400 20952 12406 20964
rect 12618 20952 12624 21004
rect 12676 20992 12682 21004
rect 13081 20995 13139 21001
rect 13081 20992 13093 20995
rect 12676 20964 13093 20992
rect 12676 20952 12682 20964
rect 13081 20961 13093 20964
rect 13127 20961 13139 20995
rect 13081 20955 13139 20961
rect 13265 20995 13323 21001
rect 13265 20961 13277 20995
rect 13311 20992 13323 20995
rect 13722 20992 13728 21004
rect 13311 20964 13728 20992
rect 13311 20961 13323 20964
rect 13265 20955 13323 20961
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 14550 20992 14556 21004
rect 14511 20964 14556 20992
rect 14550 20952 14556 20964
rect 14608 20952 14614 21004
rect 14737 20995 14795 21001
rect 14737 20961 14749 20995
rect 14783 20992 14795 20995
rect 15010 20992 15016 21004
rect 14783 20964 15016 20992
rect 14783 20961 14795 20964
rect 14737 20955 14795 20961
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 15838 20992 15844 21004
rect 15799 20964 15844 20992
rect 15838 20952 15844 20964
rect 15896 20952 15902 21004
rect 16850 20992 16856 21004
rect 16811 20964 16856 20992
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 17402 20992 17408 21004
rect 17363 20964 17408 20992
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 17512 20992 17540 21100
rect 17586 21088 17592 21140
rect 17644 21128 17650 21140
rect 21266 21128 21272 21140
rect 17644 21100 21272 21128
rect 17644 21088 17650 21100
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 24578 21128 24584 21140
rect 24539 21100 24584 21128
rect 24578 21088 24584 21100
rect 24636 21088 24642 21140
rect 25498 21088 25504 21140
rect 25556 21128 25562 21140
rect 33962 21128 33968 21140
rect 25556 21100 33968 21128
rect 25556 21088 25562 21100
rect 33962 21088 33968 21100
rect 34020 21088 34026 21140
rect 20073 21063 20131 21069
rect 20073 21029 20085 21063
rect 20119 21060 20131 21063
rect 23290 21060 23296 21072
rect 20119 21032 23296 21060
rect 20119 21029 20131 21032
rect 20073 21023 20131 21029
rect 23290 21020 23296 21032
rect 23348 21020 23354 21072
rect 27706 21060 27712 21072
rect 27667 21032 27712 21060
rect 27706 21020 27712 21032
rect 27764 21020 27770 21072
rect 19521 20995 19579 21001
rect 19521 20992 19533 20995
rect 17512 20964 19533 20992
rect 19521 20961 19533 20964
rect 19567 20961 19579 20995
rect 20714 20992 20720 21004
rect 20675 20964 20720 20992
rect 19521 20955 19579 20961
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 20990 20992 20996 21004
rect 20947 20964 20996 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 20990 20952 20996 20964
rect 21048 20952 21054 21004
rect 24670 20952 24676 21004
rect 24728 20992 24734 21004
rect 34790 20992 34796 21004
rect 24728 20964 34796 20992
rect 24728 20952 24734 20964
rect 34790 20952 34796 20964
rect 34848 20952 34854 21004
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20924 8447 20927
rect 8938 20924 8944 20936
rect 8435 20896 8944 20924
rect 8435 20893 8447 20896
rect 8389 20887 8447 20893
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 9732 20896 9777 20924
rect 9732 20884 9738 20896
rect 10226 20884 10232 20936
rect 10284 20884 10290 20936
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20924 15255 20927
rect 15378 20924 15384 20936
rect 15243 20896 15384 20924
rect 15243 20893 15255 20896
rect 15197 20887 15255 20893
rect 15378 20884 15384 20896
rect 15436 20884 15442 20936
rect 22925 20927 22983 20933
rect 22925 20924 22937 20927
rect 22066 20896 22937 20924
rect 8570 20816 8576 20868
rect 8628 20856 8634 20868
rect 10244 20856 10272 20884
rect 10413 20859 10471 20865
rect 10413 20856 10425 20859
rect 8628 20828 10180 20856
rect 10244 20828 10425 20856
rect 8628 20816 8634 20828
rect 9674 20788 9680 20800
rect 7484 20760 9680 20788
rect 7193 20751 7251 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 9769 20791 9827 20797
rect 9769 20757 9781 20791
rect 9815 20788 9827 20791
rect 10042 20788 10048 20800
rect 9815 20760 10048 20788
rect 9815 20757 9827 20760
rect 9769 20751 9827 20757
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10152 20788 10180 20828
rect 10413 20825 10425 20828
rect 10459 20825 10471 20859
rect 10413 20819 10471 20825
rect 10502 20816 10508 20868
rect 10560 20856 10566 20868
rect 10560 20828 10605 20856
rect 10560 20816 10566 20828
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 11425 20859 11483 20865
rect 11425 20856 11437 20859
rect 10928 20828 11437 20856
rect 10928 20816 10934 20828
rect 11425 20825 11437 20828
rect 11471 20825 11483 20859
rect 11425 20819 11483 20825
rect 15933 20859 15991 20865
rect 15933 20825 15945 20859
rect 15979 20856 15991 20859
rect 16758 20856 16764 20868
rect 15979 20828 16764 20856
rect 15979 20825 15991 20828
rect 15933 20819 15991 20825
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 17494 20816 17500 20868
rect 17552 20856 17558 20868
rect 18417 20859 18475 20865
rect 17552 20828 17597 20856
rect 17552 20816 17558 20828
rect 18417 20825 18429 20859
rect 18463 20825 18475 20859
rect 18417 20819 18475 20825
rect 12250 20788 12256 20800
rect 10152 20760 12256 20788
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 18432 20788 18460 20819
rect 19610 20816 19616 20868
rect 19668 20856 19674 20868
rect 19668 20828 19713 20856
rect 19668 20816 19674 20828
rect 20162 20788 20168 20800
rect 18432 20760 20168 20788
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 21361 20791 21419 20797
rect 21361 20788 21373 20791
rect 20864 20760 21373 20788
rect 20864 20748 20870 20760
rect 21361 20757 21373 20760
rect 21407 20788 21419 20791
rect 22066 20788 22094 20896
rect 22925 20893 22937 20896
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 24118 20924 24124 20936
rect 23155 20896 24124 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 24118 20884 24124 20896
rect 24176 20884 24182 20936
rect 24762 20924 24768 20936
rect 24723 20896 24768 20924
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 26789 20927 26847 20933
rect 26789 20893 26801 20927
rect 26835 20893 26847 20927
rect 26789 20887 26847 20893
rect 26881 20927 26939 20933
rect 26881 20893 26893 20927
rect 26927 20924 26939 20927
rect 33965 20927 34023 20933
rect 33965 20924 33977 20927
rect 26927 20896 33977 20924
rect 26927 20893 26939 20896
rect 26881 20887 26939 20893
rect 33965 20893 33977 20896
rect 34011 20893 34023 20927
rect 38013 20927 38071 20933
rect 38013 20924 38025 20927
rect 33965 20887 34023 20893
rect 35866 20896 38025 20924
rect 23569 20859 23627 20865
rect 23569 20825 23581 20859
rect 23615 20856 23627 20859
rect 24026 20856 24032 20868
rect 23615 20828 24032 20856
rect 23615 20825 23627 20828
rect 23569 20819 23627 20825
rect 24026 20816 24032 20828
rect 24084 20856 24090 20868
rect 26804 20856 26832 20887
rect 24084 20828 26832 20856
rect 27525 20859 27583 20865
rect 24084 20816 24090 20828
rect 27525 20825 27537 20859
rect 27571 20856 27583 20859
rect 27798 20856 27804 20868
rect 27571 20828 27804 20856
rect 27571 20825 27583 20828
rect 27525 20819 27583 20825
rect 27798 20816 27804 20828
rect 27856 20816 27862 20868
rect 21407 20760 22094 20788
rect 33781 20791 33839 20797
rect 21407 20757 21419 20760
rect 21361 20751 21419 20757
rect 33781 20757 33793 20791
rect 33827 20788 33839 20791
rect 35866 20788 35894 20896
rect 38013 20893 38025 20896
rect 38059 20893 38071 20927
rect 38013 20887 38071 20893
rect 38194 20788 38200 20800
rect 33827 20760 35894 20788
rect 38155 20760 38200 20788
rect 33827 20757 33839 20760
rect 33781 20751 33839 20757
rect 38194 20748 38200 20760
rect 38252 20748 38258 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 8846 20584 8852 20596
rect 8128 20556 8852 20584
rect 7006 20516 7012 20528
rect 6967 20488 7012 20516
rect 7006 20476 7012 20488
rect 7064 20476 7070 20528
rect 7101 20519 7159 20525
rect 7101 20485 7113 20519
rect 7147 20516 7159 20519
rect 8018 20516 8024 20528
rect 7147 20488 8024 20516
rect 7147 20485 7159 20488
rect 7101 20479 7159 20485
rect 8018 20476 8024 20488
rect 8076 20476 8082 20528
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20380 8079 20383
rect 8128 20380 8156 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 12161 20587 12219 20593
rect 8996 20556 11376 20584
rect 8996 20544 9002 20556
rect 8662 20516 8668 20528
rect 8623 20488 8668 20516
rect 8662 20476 8668 20488
rect 8720 20476 8726 20528
rect 8864 20516 8892 20544
rect 9674 20516 9680 20528
rect 8864 20488 9680 20516
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 10042 20476 10048 20528
rect 10100 20516 10106 20528
rect 10321 20519 10379 20525
rect 10321 20516 10333 20519
rect 10100 20488 10333 20516
rect 10100 20476 10106 20488
rect 10321 20485 10333 20488
rect 10367 20485 10379 20519
rect 10321 20479 10379 20485
rect 10873 20519 10931 20525
rect 10873 20485 10885 20519
rect 10919 20516 10931 20519
rect 11238 20516 11244 20528
rect 10919 20488 11244 20516
rect 10919 20485 10931 20488
rect 10873 20479 10931 20485
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 11348 20516 11376 20556
rect 12161 20553 12173 20587
rect 12207 20584 12219 20587
rect 12710 20584 12716 20596
rect 12207 20556 12716 20584
rect 12207 20553 12219 20556
rect 12161 20547 12219 20553
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12805 20587 12863 20593
rect 12805 20553 12817 20587
rect 12851 20584 12863 20587
rect 12986 20584 12992 20596
rect 12851 20556 12992 20584
rect 12851 20553 12863 20556
rect 12805 20547 12863 20553
rect 12986 20544 12992 20556
rect 13044 20544 13050 20596
rect 16758 20544 16764 20596
rect 16816 20584 16822 20596
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 16816 20556 17049 20584
rect 16816 20544 16822 20556
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 18598 20584 18604 20596
rect 17037 20547 17095 20553
rect 17144 20556 18604 20584
rect 14737 20519 14795 20525
rect 14737 20516 14749 20519
rect 11348 20488 14749 20516
rect 14737 20485 14749 20488
rect 14783 20485 14795 20519
rect 14737 20479 14795 20485
rect 15289 20519 15347 20525
rect 15289 20485 15301 20519
rect 15335 20516 15347 20519
rect 16666 20516 16672 20528
rect 15335 20488 16672 20516
rect 15335 20485 15347 20488
rect 15289 20479 15347 20485
rect 16666 20476 16672 20488
rect 16724 20476 16730 20528
rect 12069 20451 12127 20457
rect 12069 20417 12081 20451
rect 12115 20448 12127 20451
rect 12618 20448 12624 20460
rect 12115 20420 12624 20448
rect 12115 20417 12127 20420
rect 12069 20411 12127 20417
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 12713 20451 12771 20457
rect 12713 20417 12725 20451
rect 12759 20448 12771 20451
rect 13170 20448 13176 20460
rect 12759 20420 13176 20448
rect 12759 20417 12771 20420
rect 12713 20411 12771 20417
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 15746 20448 15752 20460
rect 15659 20420 15752 20448
rect 15746 20408 15752 20420
rect 15804 20448 15810 20460
rect 16298 20448 16304 20460
rect 15804 20420 16304 20448
rect 15804 20408 15810 20420
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16816 20420 16957 20448
rect 16816 20408 16822 20420
rect 16945 20417 16957 20420
rect 16991 20448 17003 20451
rect 17144 20448 17172 20556
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 19150 20544 19156 20596
rect 19208 20584 19214 20596
rect 23842 20584 23848 20596
rect 19208 20556 23848 20584
rect 19208 20544 19214 20556
rect 23842 20544 23848 20556
rect 23900 20544 23906 20596
rect 24118 20584 24124 20596
rect 24079 20556 24124 20584
rect 24118 20544 24124 20556
rect 24176 20544 24182 20596
rect 17681 20519 17739 20525
rect 17681 20485 17693 20519
rect 17727 20516 17739 20519
rect 20073 20519 20131 20525
rect 20073 20516 20085 20519
rect 17727 20488 20085 20516
rect 17727 20485 17739 20488
rect 17681 20479 17739 20485
rect 20073 20485 20085 20488
rect 20119 20485 20131 20519
rect 20073 20479 20131 20485
rect 21082 20476 21088 20528
rect 21140 20516 21146 20528
rect 23385 20519 23443 20525
rect 23385 20516 23397 20519
rect 21140 20488 23397 20516
rect 21140 20476 21146 20488
rect 23385 20485 23397 20488
rect 23431 20485 23443 20519
rect 23385 20479 23443 20485
rect 16991 20420 17172 20448
rect 17589 20451 17647 20457
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17589 20417 17601 20451
rect 17635 20417 17647 20451
rect 19150 20448 19156 20460
rect 19111 20420 19156 20448
rect 17589 20411 17647 20417
rect 8067 20352 8156 20380
rect 8573 20383 8631 20389
rect 8067 20349 8079 20352
rect 8021 20343 8079 20349
rect 8573 20349 8585 20383
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20349 8907 20383
rect 10226 20380 10232 20392
rect 10187 20352 10232 20380
rect 8849 20343 8907 20349
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 8588 20312 8616 20343
rect 7064 20284 8616 20312
rect 7064 20272 7070 20284
rect 6178 20204 6184 20256
rect 6236 20244 6242 20256
rect 8864 20244 8892 20343
rect 10226 20340 10232 20352
rect 10284 20340 10290 20392
rect 11974 20340 11980 20392
rect 12032 20380 12038 20392
rect 14366 20380 14372 20392
rect 12032 20352 14372 20380
rect 12032 20340 12038 20352
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 15378 20380 15384 20392
rect 14691 20352 15384 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 15378 20340 15384 20352
rect 15436 20340 15442 20392
rect 9122 20272 9128 20324
rect 9180 20312 9186 20324
rect 9180 20284 13952 20312
rect 9180 20272 9186 20284
rect 13262 20244 13268 20256
rect 6236 20216 13268 20244
rect 6236 20204 6242 20216
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13538 20244 13544 20256
rect 13499 20216 13544 20244
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 13924 20244 13952 20284
rect 15010 20272 15016 20324
rect 15068 20312 15074 20324
rect 17604 20312 17632 20411
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 20680 20420 21281 20448
rect 20680 20408 20686 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 24029 20451 24087 20457
rect 24029 20448 24041 20451
rect 21692 20420 24041 20448
rect 21692 20408 21698 20420
rect 24029 20417 24041 20420
rect 24075 20448 24087 20451
rect 24762 20448 24768 20460
rect 24075 20420 24768 20448
rect 24075 20417 24087 20420
rect 24029 20411 24087 20417
rect 24762 20408 24768 20420
rect 24820 20408 24826 20460
rect 29178 20448 29184 20460
rect 29139 20420 29184 20448
rect 29178 20408 29184 20420
rect 29236 20408 29242 20460
rect 33962 20448 33968 20460
rect 33923 20420 33968 20448
rect 33962 20408 33968 20420
rect 34020 20448 34026 20460
rect 37826 20448 37832 20460
rect 34020 20420 37832 20448
rect 34020 20408 34026 20420
rect 37826 20408 37832 20420
rect 37884 20408 37890 20460
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20714 20380 20720 20392
rect 20027 20352 20720 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 15068 20284 17632 20312
rect 15068 20272 15074 20284
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 20162 20312 20168 20324
rect 17736 20284 20168 20312
rect 17736 20272 17742 20284
rect 20162 20272 20168 20284
rect 20220 20272 20226 20324
rect 20533 20315 20591 20321
rect 20533 20312 20545 20315
rect 20456 20284 20545 20312
rect 14458 20244 14464 20256
rect 13924 20216 14464 20244
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 15838 20244 15844 20256
rect 15799 20216 15844 20244
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 17770 20204 17776 20256
rect 17828 20244 17834 20256
rect 19245 20247 19303 20253
rect 19245 20244 19257 20247
rect 17828 20216 19257 20244
rect 17828 20204 17834 20216
rect 19245 20213 19257 20216
rect 19291 20213 19303 20247
rect 19245 20207 19303 20213
rect 20346 20204 20352 20256
rect 20404 20244 20410 20256
rect 20456 20244 20484 20284
rect 20533 20281 20545 20284
rect 20579 20281 20591 20315
rect 20533 20275 20591 20281
rect 23569 20315 23627 20321
rect 23569 20281 23581 20315
rect 23615 20312 23627 20315
rect 27522 20312 27528 20324
rect 23615 20284 27528 20312
rect 23615 20281 23627 20284
rect 23569 20275 23627 20281
rect 27522 20272 27528 20284
rect 27580 20272 27586 20324
rect 20404 20216 20484 20244
rect 21085 20247 21143 20253
rect 20404 20204 20410 20216
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 21450 20244 21456 20256
rect 21131 20216 21456 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 28718 20204 28724 20256
rect 28776 20244 28782 20256
rect 28997 20247 29055 20253
rect 28997 20244 29009 20247
rect 28776 20216 29009 20244
rect 28776 20204 28782 20216
rect 28997 20213 29009 20216
rect 29043 20213 29055 20247
rect 28997 20207 29055 20213
rect 33502 20204 33508 20256
rect 33560 20244 33566 20256
rect 33781 20247 33839 20253
rect 33781 20244 33793 20247
rect 33560 20216 33793 20244
rect 33560 20204 33566 20216
rect 33781 20213 33793 20216
rect 33827 20213 33839 20247
rect 33781 20207 33839 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 12342 20040 12348 20052
rect 10100 20012 12348 20040
rect 10100 20000 10106 20012
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 12986 20040 12992 20052
rect 12820 20012 12992 20040
rect 9217 19975 9275 19981
rect 9217 19941 9229 19975
rect 9263 19972 9275 19975
rect 11790 19972 11796 19984
rect 9263 19944 11796 19972
rect 9263 19941 9275 19944
rect 9217 19935 9275 19941
rect 11790 19932 11796 19944
rect 11848 19932 11854 19984
rect 12069 19975 12127 19981
rect 12069 19941 12081 19975
rect 12115 19972 12127 19975
rect 12820 19972 12848 20012
rect 12986 20000 12992 20012
rect 13044 20040 13050 20052
rect 15654 20040 15660 20052
rect 13044 20012 15660 20040
rect 13044 20000 13050 20012
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16574 20040 16580 20052
rect 16535 20012 16580 20040
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 19484 20012 19533 20040
rect 19484 20000 19490 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 20346 20040 20352 20052
rect 19521 20003 19579 20009
rect 20272 20012 20352 20040
rect 12115 19944 12848 19972
rect 12115 19941 12127 19944
rect 12069 19935 12127 19941
rect 12894 19932 12900 19984
rect 12952 19972 12958 19984
rect 12952 19944 20208 19972
rect 12952 19932 12958 19944
rect 10229 19907 10287 19913
rect 10229 19873 10241 19907
rect 10275 19904 10287 19907
rect 12526 19904 12532 19916
rect 10275 19876 12532 19904
rect 10275 19873 10287 19876
rect 10229 19867 10287 19873
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 12713 19907 12771 19913
rect 12713 19873 12725 19907
rect 12759 19904 12771 19907
rect 13354 19904 13360 19916
rect 12759 19876 13360 19904
rect 12759 19873 12771 19876
rect 12713 19867 12771 19873
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 13722 19904 13728 19916
rect 13683 19876 13728 19904
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 14550 19864 14556 19916
rect 14608 19904 14614 19916
rect 15013 19907 15071 19913
rect 15013 19904 15025 19907
rect 14608 19876 15025 19904
rect 14608 19864 14614 19876
rect 15013 19873 15025 19876
rect 15059 19873 15071 19907
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 15013 19867 15071 19873
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 16301 19907 16359 19913
rect 16301 19873 16313 19907
rect 16347 19904 16359 19907
rect 16942 19904 16948 19916
rect 16347 19876 16948 19904
rect 16347 19873 16359 19876
rect 16301 19867 16359 19873
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 20180 19913 20208 19944
rect 20165 19907 20223 19913
rect 19306 19876 20116 19904
rect 7558 19796 7564 19848
rect 7616 19836 7622 19848
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 7616 19808 7941 19836
rect 7616 19796 7622 19808
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 8352 19808 9137 19836
rect 8352 19796 8358 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 9214 19796 9220 19848
rect 9272 19836 9278 19848
rect 10137 19839 10195 19845
rect 10137 19836 10149 19839
rect 9272 19808 10149 19836
rect 9272 19796 9278 19808
rect 10137 19805 10149 19808
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19836 10839 19839
rect 10962 19836 10968 19848
rect 10827 19808 10968 19836
rect 10827 19805 10839 19808
rect 10781 19799 10839 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 14274 19836 14280 19848
rect 14235 19808 14280 19836
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 19306 19836 19334 19876
rect 15712 19808 19334 19836
rect 19429 19839 19487 19845
rect 15712 19796 15718 19808
rect 19429 19805 19441 19839
rect 19475 19805 19487 19839
rect 20088 19836 20116 19876
rect 20165 19873 20177 19907
rect 20211 19873 20223 19907
rect 20165 19867 20223 19873
rect 20272 19836 20300 20012
rect 20346 20000 20352 20012
rect 20404 20040 20410 20052
rect 20622 20040 20628 20052
rect 20404 20012 20628 20040
rect 20404 20000 20410 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 20806 20040 20812 20052
rect 20767 20012 20812 20040
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 22664 20012 28672 20040
rect 21269 19975 21327 19981
rect 21269 19941 21281 19975
rect 21315 19941 21327 19975
rect 21269 19935 21327 19941
rect 20349 19907 20407 19913
rect 20349 19873 20361 19907
rect 20395 19904 20407 19907
rect 21284 19904 21312 19935
rect 20395 19876 21312 19904
rect 20395 19873 20407 19876
rect 20349 19867 20407 19873
rect 21450 19836 21456 19848
rect 20088 19808 20300 19836
rect 21411 19808 21456 19836
rect 19429 19799 19487 19805
rect 6825 19771 6883 19777
rect 6825 19737 6837 19771
rect 6871 19737 6883 19771
rect 6825 19731 6883 19737
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 6840 19700 6868 19731
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 6972 19740 7017 19768
rect 6972 19728 6978 19740
rect 7098 19728 7104 19780
rect 7156 19768 7162 19780
rect 7466 19768 7472 19780
rect 7156 19740 7472 19768
rect 7156 19728 7162 19740
rect 7466 19728 7472 19740
rect 7524 19728 7530 19780
rect 10410 19728 10416 19780
rect 10468 19768 10474 19780
rect 11517 19771 11575 19777
rect 11517 19768 11529 19771
rect 10468 19740 11529 19768
rect 10468 19728 10474 19740
rect 11517 19737 11529 19740
rect 11563 19737 11575 19771
rect 11517 19731 11575 19737
rect 11606 19728 11612 19780
rect 11664 19768 11670 19780
rect 12805 19771 12863 19777
rect 11664 19740 11709 19768
rect 11664 19728 11670 19740
rect 12805 19737 12817 19771
rect 12851 19768 12863 19771
rect 13538 19768 13544 19780
rect 12851 19740 13544 19768
rect 12851 19737 12863 19740
rect 12805 19731 12863 19737
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 15102 19728 15108 19780
rect 15160 19768 15166 19780
rect 15160 19740 15205 19768
rect 15160 19728 15166 19740
rect 17218 19728 17224 19780
rect 17276 19768 17282 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 17276 19740 17325 19768
rect 17276 19728 17282 19740
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17494 19768 17500 19780
rect 17455 19740 17500 19768
rect 17313 19731 17371 19737
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 17586 19728 17592 19780
rect 17644 19768 17650 19780
rect 19444 19768 19472 19799
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 22664 19845 22692 20012
rect 26234 19932 26240 19984
rect 26292 19972 26298 19984
rect 27065 19975 27123 19981
rect 27065 19972 27077 19975
rect 26292 19944 27077 19972
rect 26292 19932 26298 19944
rect 27065 19941 27077 19944
rect 27111 19941 27123 19975
rect 27065 19935 27123 19941
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19904 26939 19907
rect 28537 19907 28595 19913
rect 28537 19904 28549 19907
rect 26927 19876 28549 19904
rect 26927 19873 26939 19876
rect 26881 19867 26939 19873
rect 28537 19873 28549 19876
rect 28583 19873 28595 19907
rect 28537 19867 28595 19873
rect 22649 19839 22707 19845
rect 22649 19836 22661 19839
rect 22066 19808 22661 19836
rect 21818 19768 21824 19780
rect 17644 19740 19380 19768
rect 19444 19740 21824 19768
rect 17644 19728 17650 19740
rect 10870 19700 10876 19712
rect 6788 19672 6868 19700
rect 10831 19672 10876 19700
rect 6788 19660 6794 19672
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 13354 19660 13360 19712
rect 13412 19700 13418 19712
rect 14274 19700 14280 19712
rect 13412 19672 14280 19700
rect 13412 19660 13418 19672
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 14369 19703 14427 19709
rect 14369 19669 14381 19703
rect 14415 19700 14427 19703
rect 14642 19700 14648 19712
rect 14415 19672 14648 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 19352 19700 19380 19740
rect 21818 19728 21824 19740
rect 21876 19728 21882 19780
rect 22066 19700 22094 19808
rect 22649 19805 22661 19808
rect 22695 19805 22707 19839
rect 22649 19799 22707 19805
rect 26697 19839 26755 19845
rect 26697 19805 26709 19839
rect 26743 19805 26755 19839
rect 27798 19836 27804 19848
rect 27711 19808 27804 19836
rect 26697 19799 26755 19805
rect 26712 19768 26740 19799
rect 27798 19796 27804 19808
rect 27856 19836 27862 19848
rect 28445 19839 28503 19845
rect 27856 19808 28028 19836
rect 27856 19796 27862 19808
rect 27246 19768 27252 19780
rect 26712 19740 27252 19768
rect 27246 19728 27252 19740
rect 27304 19768 27310 19780
rect 27893 19771 27951 19777
rect 27893 19768 27905 19771
rect 27304 19740 27905 19768
rect 27304 19728 27310 19740
rect 27893 19737 27905 19740
rect 27939 19737 27951 19771
rect 28000 19768 28028 19808
rect 28445 19805 28457 19839
rect 28491 19836 28503 19839
rect 28644 19836 28672 20012
rect 29178 19836 29184 19848
rect 28491 19808 29184 19836
rect 28491 19805 28503 19808
rect 28445 19799 28503 19805
rect 29178 19796 29184 19808
rect 29236 19796 29242 19848
rect 30837 19839 30895 19845
rect 30837 19805 30849 19839
rect 30883 19836 30895 19839
rect 34698 19836 34704 19848
rect 30883 19808 34704 19836
rect 30883 19805 30895 19808
rect 30837 19799 30895 19805
rect 34698 19796 34704 19808
rect 34756 19796 34762 19848
rect 28626 19768 28632 19780
rect 28000 19740 28632 19768
rect 27893 19731 27951 19737
rect 28626 19728 28632 19740
rect 28684 19728 28690 19780
rect 19352 19672 22094 19700
rect 22465 19703 22523 19709
rect 22465 19669 22477 19703
rect 22511 19700 22523 19703
rect 23750 19700 23756 19712
rect 22511 19672 23756 19700
rect 22511 19669 22523 19672
rect 22465 19663 22523 19669
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 26142 19660 26148 19712
rect 26200 19700 26206 19712
rect 30929 19703 30987 19709
rect 30929 19700 30941 19703
rect 26200 19672 30941 19700
rect 26200 19660 26206 19672
rect 30929 19669 30941 19672
rect 30975 19669 30987 19703
rect 30929 19663 30987 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 5813 19499 5871 19505
rect 5813 19465 5825 19499
rect 5859 19496 5871 19499
rect 6822 19496 6828 19508
rect 5859 19468 6828 19496
rect 5859 19465 5871 19468
rect 5813 19459 5871 19465
rect 1596 19428 1624 19459
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 7374 19456 7380 19508
rect 7432 19496 7438 19508
rect 7745 19499 7803 19505
rect 7745 19496 7757 19499
rect 7432 19468 7757 19496
rect 7432 19456 7438 19468
rect 7745 19465 7757 19468
rect 7791 19465 7803 19499
rect 7745 19459 7803 19465
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8076 19468 8984 19496
rect 8076 19456 8082 19468
rect 8956 19428 8984 19468
rect 9030 19456 9036 19508
rect 9088 19496 9094 19508
rect 9125 19499 9183 19505
rect 9125 19496 9137 19499
rect 9088 19468 9137 19496
rect 9088 19456 9094 19468
rect 9125 19465 9137 19468
rect 9171 19465 9183 19499
rect 9125 19459 9183 19465
rect 9769 19499 9827 19505
rect 9769 19465 9781 19499
rect 9815 19496 9827 19499
rect 11606 19496 11612 19508
rect 9815 19468 11612 19496
rect 9815 19465 9827 19468
rect 9769 19459 9827 19465
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 12894 19496 12900 19508
rect 11756 19468 12900 19496
rect 11756 19456 11762 19468
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 23474 19496 23480 19508
rect 15028 19468 23480 19496
rect 10686 19428 10692 19440
rect 1596 19400 8800 19428
rect 8956 19400 9720 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 5994 19360 6000 19372
rect 4847 19332 5856 19360
rect 5955 19332 6000 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 5828 19292 5856 19332
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 6914 19360 6920 19372
rect 6104 19332 6920 19360
rect 6104 19292 6132 19332
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7101 19363 7159 19369
rect 7101 19329 7113 19363
rect 7147 19329 7159 19363
rect 7101 19323 7159 19329
rect 5828 19264 6132 19292
rect 7116 19292 7144 19323
rect 7190 19320 7196 19372
rect 7248 19360 7254 19372
rect 7926 19360 7932 19372
rect 7248 19332 7293 19360
rect 7887 19332 7932 19360
rect 7248 19320 7254 19332
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 8772 19364 8800 19400
rect 9692 19369 9720 19400
rect 10428 19400 10692 19428
rect 10428 19369 10456 19400
rect 10686 19388 10692 19400
rect 10744 19388 10750 19440
rect 10870 19388 10876 19440
rect 10928 19428 10934 19440
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 10928 19400 12173 19428
rect 10928 19388 10934 19400
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 13725 19431 13783 19437
rect 13725 19428 13737 19431
rect 12400 19400 13737 19428
rect 12400 19388 12406 19400
rect 13725 19397 13737 19400
rect 13771 19397 13783 19431
rect 14642 19428 14648 19440
rect 14555 19400 14648 19428
rect 13725 19391 13783 19397
rect 14642 19388 14648 19400
rect 14700 19428 14706 19440
rect 14918 19428 14924 19440
rect 14700 19400 14924 19428
rect 14700 19388 14706 19400
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 8772 19360 8892 19364
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8772 19336 9045 19360
rect 8864 19332 9045 19336
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19329 9735 19363
rect 9677 19323 9735 19329
rect 10413 19363 10471 19369
rect 10413 19329 10425 19363
rect 10459 19329 10471 19363
rect 10413 19323 10471 19329
rect 10502 19320 10508 19372
rect 10560 19360 10566 19372
rect 10560 19332 10605 19360
rect 10560 19320 10566 19332
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 10836 19332 11928 19360
rect 10836 19320 10842 19332
rect 8294 19292 8300 19304
rect 7116 19264 8300 19292
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 9214 19292 9220 19304
rect 8435 19264 9220 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 11606 19292 11612 19304
rect 9324 19264 11612 19292
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 9324 19224 9352 19264
rect 11606 19252 11612 19264
rect 11664 19252 11670 19304
rect 11900 19292 11928 19332
rect 13004 19332 13216 19360
rect 12069 19295 12127 19301
rect 12069 19292 12081 19295
rect 11900 19264 12081 19292
rect 12069 19261 12081 19264
rect 12115 19261 12127 19295
rect 12069 19255 12127 19261
rect 12342 19252 12348 19304
rect 12400 19292 12406 19304
rect 13004 19292 13032 19332
rect 12400 19264 13032 19292
rect 13081 19295 13139 19301
rect 12400 19252 12406 19264
rect 13081 19261 13093 19295
rect 13127 19261 13139 19295
rect 13188 19292 13216 19332
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 15028 19360 15056 19468
rect 15194 19428 15200 19440
rect 15155 19400 15200 19428
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 15289 19431 15347 19437
rect 15289 19397 15301 19431
rect 15335 19428 15347 19431
rect 15562 19428 15568 19440
rect 15335 19400 15568 19428
rect 15335 19397 15347 19400
rect 15289 19391 15347 19397
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 16224 19437 16252 19468
rect 23474 19456 23480 19468
rect 23532 19456 23538 19508
rect 16209 19431 16267 19437
rect 16209 19397 16221 19431
rect 16255 19397 16267 19431
rect 17586 19428 17592 19440
rect 16209 19391 16267 19397
rect 16316 19400 17592 19428
rect 16316 19360 16344 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 17954 19428 17960 19440
rect 17915 19400 17960 19428
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 18046 19388 18052 19440
rect 18104 19428 18110 19440
rect 19426 19428 19432 19440
rect 18104 19400 19432 19428
rect 18104 19388 18110 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 13320 19332 13492 19360
rect 13320 19320 13326 19332
rect 13464 19292 13492 19332
rect 14476 19332 15056 19360
rect 16040 19332 16344 19360
rect 16945 19363 17003 19369
rect 13633 19295 13691 19301
rect 13633 19292 13645 19295
rect 13188 19264 13400 19292
rect 13464 19264 13645 19292
rect 13081 19255 13139 19261
rect 8168 19196 9352 19224
rect 13096 19224 13124 19255
rect 13262 19224 13268 19236
rect 13096 19196 13268 19224
rect 8168 19184 8174 19196
rect 13262 19184 13268 19196
rect 13320 19184 13326 19236
rect 13372 19224 13400 19264
rect 13633 19261 13645 19264
rect 13679 19292 13691 19295
rect 14476 19292 14504 19332
rect 13679 19264 14504 19292
rect 16040 19280 16068 19332
rect 16945 19329 16957 19363
rect 16991 19360 17003 19363
rect 17678 19360 17684 19372
rect 16991 19332 17684 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 20916 19332 22017 19360
rect 17862 19292 17868 19304
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 15948 19252 16068 19280
rect 17823 19264 17868 19292
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 18230 19292 18236 19304
rect 18191 19264 18236 19292
rect 18230 19252 18236 19264
rect 18288 19252 18294 19304
rect 19429 19295 19487 19301
rect 19429 19261 19441 19295
rect 19475 19292 19487 19295
rect 19518 19292 19524 19304
rect 19475 19264 19524 19292
rect 19475 19261 19487 19264
rect 19429 19255 19487 19261
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 14550 19224 14556 19236
rect 13372 19196 14556 19224
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 4617 19159 4675 19165
rect 4617 19125 4629 19159
rect 4663 19156 4675 19159
rect 4706 19156 4712 19168
rect 4663 19128 4712 19156
rect 4663 19125 4675 19128
rect 4617 19119 4675 19125
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 9122 19156 9128 19168
rect 7984 19128 9128 19156
rect 7984 19116 7990 19128
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 13538 19156 13544 19168
rect 9640 19128 13544 19156
rect 9640 19116 9646 19128
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 15948 19156 15976 19252
rect 20916 19236 20944 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 28718 19360 28724 19372
rect 28679 19332 28724 19360
rect 22005 19323 22063 19329
rect 28718 19320 28724 19332
rect 28776 19320 28782 19372
rect 30098 19360 30104 19372
rect 30059 19332 30104 19360
rect 30098 19320 30104 19332
rect 30156 19320 30162 19372
rect 30190 19320 30196 19372
rect 30248 19360 30254 19372
rect 38102 19360 38108 19372
rect 30248 19332 30293 19360
rect 38063 19332 38108 19360
rect 30248 19320 30254 19332
rect 38102 19320 38108 19332
rect 38160 19320 38166 19372
rect 16666 19184 16672 19236
rect 16724 19224 16730 19236
rect 16724 19196 17080 19224
rect 16724 19184 16730 19196
rect 17052 19165 17080 19196
rect 17218 19184 17224 19236
rect 17276 19224 17282 19236
rect 20898 19224 20904 19236
rect 17276 19196 20904 19224
rect 17276 19184 17282 19196
rect 17880 19168 17908 19196
rect 20898 19184 20904 19196
rect 20956 19184 20962 19236
rect 14792 19128 15976 19156
rect 17037 19159 17095 19165
rect 14792 19116 14798 19128
rect 17037 19125 17049 19159
rect 17083 19125 17095 19159
rect 17037 19119 17095 19125
rect 17862 19116 17868 19168
rect 17920 19116 17926 19168
rect 22097 19159 22155 19165
rect 22097 19125 22109 19159
rect 22143 19156 22155 19159
rect 22554 19156 22560 19168
rect 22143 19128 22560 19156
rect 22143 19125 22155 19128
rect 22097 19119 22155 19125
rect 22554 19116 22560 19128
rect 22612 19116 22618 19168
rect 28534 19156 28540 19168
rect 28495 19128 28540 19156
rect 28534 19116 28540 19128
rect 28592 19116 28598 19168
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 6052 18924 6469 18952
rect 6052 18912 6058 18924
rect 6457 18921 6469 18924
rect 6503 18921 6515 18955
rect 6457 18915 6515 18921
rect 7837 18955 7895 18961
rect 7837 18921 7849 18955
rect 7883 18952 7895 18955
rect 8478 18952 8484 18964
rect 7883 18924 8484 18952
rect 7883 18921 7895 18924
rect 7837 18915 7895 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 10318 18912 10324 18964
rect 10376 18952 10382 18964
rect 16850 18952 16856 18964
rect 10376 18924 16856 18952
rect 10376 18912 10382 18924
rect 16850 18912 16856 18924
rect 16908 18912 16914 18964
rect 16942 18912 16948 18964
rect 17000 18952 17006 18964
rect 21082 18952 21088 18964
rect 17000 18924 21088 18952
rect 17000 18912 17006 18924
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 13722 18884 13728 18896
rect 7524 18856 9536 18884
rect 7524 18844 7530 18856
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 9214 18816 9220 18828
rect 7340 18788 9076 18816
rect 9175 18788 9220 18816
rect 7340 18776 7346 18788
rect 4706 18748 4712 18760
rect 4667 18720 4712 18748
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 5997 18751 6055 18757
rect 5997 18748 6009 18751
rect 5868 18720 6009 18748
rect 5868 18708 5874 18720
rect 5997 18717 6009 18720
rect 6043 18717 6055 18751
rect 5997 18711 6055 18717
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7374 18748 7380 18760
rect 7147 18720 7380 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 6656 18680 6684 18711
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 7742 18748 7748 18760
rect 7703 18720 7748 18748
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 8389 18751 8447 18757
rect 8389 18748 8401 18751
rect 8352 18720 8401 18748
rect 8352 18708 8358 18720
rect 8389 18717 8401 18720
rect 8435 18748 8447 18751
rect 8754 18748 8760 18760
rect 8435 18720 8760 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 7760 18680 7788 18708
rect 6656 18652 7788 18680
rect 9048 18680 9076 18788
rect 9214 18776 9220 18788
rect 9272 18776 9278 18828
rect 9508 18825 9536 18856
rect 10704 18856 13728 18884
rect 9493 18819 9551 18825
rect 9493 18785 9505 18819
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 10134 18776 10140 18828
rect 10192 18816 10198 18828
rect 10704 18825 10732 18856
rect 13722 18844 13728 18856
rect 13780 18844 13786 18896
rect 14550 18844 14556 18896
rect 14608 18884 14614 18896
rect 26510 18884 26516 18896
rect 14608 18856 19840 18884
rect 14608 18844 14614 18856
rect 10689 18819 10747 18825
rect 10689 18816 10701 18819
rect 10192 18788 10701 18816
rect 10192 18776 10198 18788
rect 10689 18785 10701 18788
rect 10735 18785 10747 18819
rect 11054 18816 11060 18828
rect 11015 18788 11060 18816
rect 10689 18779 10747 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 12342 18816 12348 18828
rect 11992 18788 12348 18816
rect 11992 18757 12020 18788
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 12713 18819 12771 18825
rect 12713 18785 12725 18819
rect 12759 18816 12771 18819
rect 12986 18816 12992 18828
rect 12759 18788 12992 18816
rect 12759 18785 12771 18788
rect 12713 18779 12771 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 14642 18816 14648 18828
rect 13679 18788 14648 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 15013 18819 15071 18825
rect 15013 18785 15025 18819
rect 15059 18816 15071 18819
rect 15838 18816 15844 18828
rect 15059 18788 15844 18816
rect 15059 18785 15071 18788
rect 15013 18779 15071 18785
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 17402 18816 17408 18828
rect 16684 18788 17408 18816
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18717 12035 18751
rect 11977 18711 12035 18717
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12216 18720 12572 18748
rect 12216 18708 12222 18720
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 9048 18652 9321 18680
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9309 18643 9367 18649
rect 10778 18640 10784 18692
rect 10836 18680 10842 18692
rect 12069 18683 12127 18689
rect 10836 18652 10881 18680
rect 10836 18640 10842 18652
rect 12069 18649 12081 18683
rect 12115 18649 12127 18683
rect 12544 18680 12572 18720
rect 14458 18708 14464 18760
rect 14516 18748 14522 18760
rect 14817 18751 14875 18757
rect 14817 18748 14829 18751
rect 14516 18720 14829 18748
rect 14516 18708 14522 18720
rect 14817 18717 14829 18720
rect 14863 18717 14875 18751
rect 16022 18748 16028 18760
rect 15983 18720 16028 18748
rect 14817 18711 14875 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 16684 18757 16712 18788
rect 17402 18776 17408 18788
rect 17460 18776 17466 18828
rect 19518 18816 19524 18828
rect 19479 18788 19524 18816
rect 19518 18776 19524 18788
rect 19576 18776 19582 18828
rect 19812 18825 19840 18856
rect 22066 18856 26516 18884
rect 19797 18819 19855 18825
rect 19797 18785 19809 18819
rect 19843 18816 19855 18819
rect 22066 18816 22094 18856
rect 26510 18844 26516 18856
rect 26568 18844 26574 18896
rect 22462 18816 22468 18828
rect 19843 18788 22094 18816
rect 22423 18788 22468 18816
rect 19843 18785 19855 18788
rect 19797 18779 19855 18785
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 24670 18776 24676 18828
rect 24728 18816 24734 18828
rect 24728 18788 26188 18816
rect 24728 18776 24734 18788
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16172 18720 16681 18748
rect 16172 18708 16178 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17497 18751 17555 18757
rect 17497 18748 17509 18751
rect 17276 18720 17509 18748
rect 17276 18708 17282 18720
rect 17497 18717 17509 18720
rect 17543 18717 17555 18751
rect 17497 18711 17555 18717
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 18693 18751 18751 18757
rect 18693 18748 18705 18751
rect 18564 18720 18705 18748
rect 18564 18708 18570 18720
rect 18693 18717 18705 18720
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21177 18751 21235 18757
rect 21177 18748 21189 18751
rect 20956 18720 21189 18748
rect 20956 18708 20962 18720
rect 21177 18717 21189 18720
rect 21223 18717 21235 18751
rect 23750 18748 23756 18760
rect 23711 18720 23756 18748
rect 21177 18711 21235 18717
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 26160 18757 26188 18788
rect 27522 18776 27528 18828
rect 27580 18816 27586 18828
rect 35986 18816 35992 18828
rect 27580 18788 35992 18816
rect 27580 18776 27586 18788
rect 35986 18776 35992 18788
rect 36044 18776 36050 18828
rect 25409 18751 25467 18757
rect 25409 18717 25421 18751
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 26145 18751 26203 18757
rect 26145 18717 26157 18751
rect 26191 18748 26203 18751
rect 27249 18751 27307 18757
rect 27249 18748 27261 18751
rect 26191 18720 27261 18748
rect 26191 18717 26203 18720
rect 26145 18711 26203 18717
rect 27249 18717 27261 18720
rect 27295 18717 27307 18751
rect 27249 18711 27307 18717
rect 12805 18683 12863 18689
rect 12805 18680 12817 18683
rect 12544 18652 12817 18680
rect 12069 18643 12127 18649
rect 12805 18649 12817 18652
rect 12851 18649 12863 18683
rect 16040 18680 16068 18708
rect 18785 18683 18843 18689
rect 16040 18652 17724 18680
rect 12805 18643 12863 18649
rect 4338 18572 4344 18624
rect 4396 18612 4402 18624
rect 4525 18615 4583 18621
rect 4525 18612 4537 18615
rect 4396 18584 4537 18612
rect 4396 18572 4402 18584
rect 4525 18581 4537 18584
rect 4571 18581 4583 18615
rect 4525 18575 4583 18581
rect 5813 18615 5871 18621
rect 5813 18581 5825 18615
rect 5859 18612 5871 18615
rect 6454 18612 6460 18624
rect 5859 18584 6460 18612
rect 5859 18581 5871 18584
rect 5813 18575 5871 18581
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 7156 18584 7205 18612
rect 7156 18572 7162 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7193 18575 7251 18581
rect 8481 18615 8539 18621
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 9122 18612 9128 18624
rect 8527 18584 9128 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 11330 18612 11336 18624
rect 9272 18584 11336 18612
rect 9272 18572 9278 18584
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 12084 18612 12112 18643
rect 12710 18612 12716 18624
rect 12084 18584 12716 18612
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 15473 18615 15531 18621
rect 15473 18612 15485 18615
rect 15344 18584 15485 18612
rect 15344 18572 15350 18584
rect 15473 18581 15485 18584
rect 15519 18581 15531 18615
rect 15473 18575 15531 18581
rect 15562 18572 15568 18624
rect 15620 18612 15626 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15620 18584 16129 18612
rect 15620 18572 15626 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16117 18575 16175 18581
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 16761 18615 16819 18621
rect 16761 18612 16773 18615
rect 16356 18584 16773 18612
rect 16356 18572 16362 18584
rect 16761 18581 16773 18584
rect 16807 18581 16819 18615
rect 16761 18575 16819 18581
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17589 18615 17647 18621
rect 17589 18612 17601 18615
rect 17092 18584 17601 18612
rect 17092 18572 17098 18584
rect 17589 18581 17601 18584
rect 17635 18581 17647 18615
rect 17696 18612 17724 18652
rect 18785 18649 18797 18683
rect 18831 18680 18843 18683
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 18831 18652 19625 18680
rect 18831 18649 18843 18652
rect 18785 18643 18843 18649
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 20990 18680 20996 18692
rect 19613 18643 19671 18649
rect 19720 18652 20996 18680
rect 19720 18612 19748 18652
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 22554 18680 22560 18692
rect 22515 18652 22560 18680
rect 22554 18640 22560 18652
rect 22612 18640 22618 18692
rect 23109 18683 23167 18689
rect 23109 18649 23121 18683
rect 23155 18680 23167 18683
rect 23198 18680 23204 18692
rect 23155 18652 23204 18680
rect 23155 18649 23167 18652
rect 23109 18643 23167 18649
rect 23198 18640 23204 18652
rect 23256 18640 23262 18692
rect 25424 18680 25452 18711
rect 26694 18680 26700 18692
rect 25424 18652 26700 18680
rect 26694 18640 26700 18652
rect 26752 18640 26758 18692
rect 17696 18584 19748 18612
rect 17589 18575 17647 18581
rect 20346 18572 20352 18624
rect 20404 18612 20410 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 20404 18584 21281 18612
rect 20404 18572 20410 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 23569 18615 23627 18621
rect 23569 18581 23581 18615
rect 23615 18612 23627 18615
rect 23750 18612 23756 18624
rect 23615 18584 23756 18612
rect 23615 18581 23627 18584
rect 23569 18575 23627 18581
rect 23750 18572 23756 18584
rect 23808 18572 23814 18624
rect 24854 18612 24860 18624
rect 24815 18584 24860 18612
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 25498 18612 25504 18624
rect 25459 18584 25504 18612
rect 25498 18572 25504 18584
rect 25556 18572 25562 18624
rect 26237 18615 26295 18621
rect 26237 18581 26249 18615
rect 26283 18612 26295 18615
rect 26326 18612 26332 18624
rect 26283 18584 26332 18612
rect 26283 18581 26295 18584
rect 26237 18575 26295 18581
rect 26326 18572 26332 18584
rect 26384 18572 26390 18624
rect 27065 18615 27123 18621
rect 27065 18581 27077 18615
rect 27111 18612 27123 18615
rect 27706 18612 27712 18624
rect 27111 18584 27712 18612
rect 27111 18581 27123 18584
rect 27065 18575 27123 18581
rect 27706 18572 27712 18584
rect 27764 18572 27770 18624
rect 28077 18615 28135 18621
rect 28077 18581 28089 18615
rect 28123 18612 28135 18615
rect 28350 18612 28356 18624
rect 28123 18584 28356 18612
rect 28123 18581 28135 18584
rect 28077 18575 28135 18581
rect 28350 18572 28356 18584
rect 28408 18572 28414 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 5810 18408 5816 18420
rect 5771 18380 5816 18408
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 8481 18411 8539 18417
rect 8481 18377 8493 18411
rect 8527 18408 8539 18411
rect 10778 18408 10784 18420
rect 8527 18380 10784 18408
rect 8527 18377 8539 18380
rect 8481 18371 8539 18377
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11054 18368 11060 18420
rect 11112 18408 11118 18420
rect 11698 18408 11704 18420
rect 11112 18380 11704 18408
rect 11112 18368 11118 18380
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 11793 18411 11851 18417
rect 11793 18377 11805 18411
rect 11839 18408 11851 18411
rect 12989 18411 13047 18417
rect 11839 18380 12756 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 4338 18340 4344 18352
rect 4299 18312 4344 18340
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 7650 18300 7656 18352
rect 7708 18340 7714 18352
rect 9125 18343 9183 18349
rect 7708 18312 9076 18340
rect 7708 18300 7714 18312
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 5997 18275 6055 18281
rect 5997 18272 6009 18275
rect 5776 18244 6009 18272
rect 5776 18232 5782 18244
rect 5997 18241 6009 18244
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 6972 18244 7113 18272
rect 6972 18232 6978 18244
rect 7101 18241 7113 18244
rect 7147 18272 7159 18275
rect 7282 18272 7288 18284
rect 7147 18244 7288 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 4249 18207 4307 18213
rect 4249 18173 4261 18207
rect 4295 18204 4307 18207
rect 4614 18204 4620 18216
rect 4295 18176 4620 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 4890 18204 4896 18216
rect 4851 18176 4896 18204
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 7760 18204 7788 18235
rect 7926 18232 7932 18284
rect 7984 18272 7990 18284
rect 9048 18281 9076 18312
rect 9125 18309 9137 18343
rect 9171 18340 9183 18343
rect 12728 18340 12756 18380
rect 12989 18377 13001 18411
rect 13035 18408 13047 18411
rect 15286 18408 15292 18420
rect 13035 18380 15292 18408
rect 13035 18377 13047 18380
rect 12989 18371 13047 18377
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 15764 18380 18521 18408
rect 13633 18343 13691 18349
rect 13633 18340 13645 18343
rect 9171 18312 11836 18340
rect 12728 18312 13645 18340
rect 9171 18309 9183 18312
rect 9125 18303 9183 18309
rect 8389 18275 8447 18281
rect 8389 18272 8401 18275
rect 7984 18244 8401 18272
rect 7984 18232 7990 18244
rect 8389 18241 8401 18244
rect 8435 18241 8447 18275
rect 8389 18235 8447 18241
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9214 18232 9220 18284
rect 9272 18272 9278 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9272 18244 9689 18272
rect 9272 18232 9278 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18272 10563 18275
rect 10870 18272 10876 18284
rect 10551 18244 10876 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11698 18272 11704 18284
rect 11020 18244 11065 18272
rect 11659 18244 11704 18272
rect 11020 18232 11026 18244
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 11808 18272 11836 18312
rect 13633 18309 13645 18312
rect 13679 18309 13691 18343
rect 14550 18340 14556 18352
rect 14511 18312 14556 18340
rect 13633 18303 13691 18309
rect 14550 18300 14556 18312
rect 14608 18300 14614 18352
rect 15764 18349 15792 18380
rect 18509 18377 18521 18380
rect 18555 18377 18567 18411
rect 18509 18371 18567 18377
rect 21269 18411 21327 18417
rect 21269 18377 21281 18411
rect 21315 18408 21327 18411
rect 21315 18380 27384 18408
rect 21315 18377 21327 18380
rect 21269 18371 21327 18377
rect 15742 18343 15800 18349
rect 15742 18309 15754 18343
rect 15788 18309 15800 18343
rect 15742 18303 15800 18309
rect 16942 18300 16948 18352
rect 17000 18340 17006 18352
rect 17037 18343 17095 18349
rect 17037 18340 17049 18343
rect 17000 18312 17049 18340
rect 17000 18300 17006 18312
rect 17037 18309 17049 18312
rect 17083 18309 17095 18343
rect 17037 18303 17095 18309
rect 17402 18300 17408 18352
rect 17460 18340 17466 18352
rect 22186 18340 22192 18352
rect 17460 18312 20484 18340
rect 22147 18312 22192 18340
rect 17460 18300 17466 18312
rect 12158 18272 12164 18284
rect 11808 18244 12164 18272
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12268 18244 12480 18272
rect 12268 18204 12296 18244
rect 7760 18176 12296 18204
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18173 12403 18207
rect 12452 18204 12480 18244
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 18414 18272 18420 18284
rect 12584 18244 12629 18272
rect 18375 18244 18420 18272
rect 12584 18232 12590 18244
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 19610 18272 19616 18284
rect 18748 18244 19616 18272
rect 18748 18232 18754 18244
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 20456 18281 20484 18312
rect 22186 18300 22192 18312
rect 22244 18300 22250 18352
rect 24854 18340 24860 18352
rect 24815 18312 24860 18340
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 26050 18340 26056 18352
rect 26011 18312 26056 18340
rect 26050 18300 26056 18312
rect 26108 18300 26114 18352
rect 27246 18340 27252 18352
rect 27207 18312 27252 18340
rect 27246 18300 27252 18312
rect 27304 18300 27310 18352
rect 27356 18349 27384 18380
rect 27341 18343 27399 18349
rect 27341 18309 27353 18343
rect 27387 18309 27399 18343
rect 27341 18303 27399 18309
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 21082 18232 21088 18284
rect 21140 18272 21146 18284
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 21140 18244 21189 18272
rect 21140 18232 21146 18244
rect 21177 18241 21189 18244
rect 21223 18272 21235 18275
rect 21450 18272 21456 18284
rect 21223 18244 21456 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 21450 18232 21456 18244
rect 21508 18232 21514 18284
rect 23750 18272 23756 18284
rect 23711 18244 23756 18272
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 28350 18272 28356 18284
rect 28311 18244 28356 18272
rect 28350 18232 28356 18244
rect 28408 18232 28414 18284
rect 28534 18272 28540 18284
rect 28495 18244 28540 18272
rect 28534 18232 28540 18244
rect 28592 18232 28598 18284
rect 13538 18204 13544 18216
rect 12452 18176 13216 18204
rect 13499 18176 13544 18204
rect 12345 18167 12403 18173
rect 7837 18139 7895 18145
rect 7837 18105 7849 18139
rect 7883 18136 7895 18139
rect 9858 18136 9864 18148
rect 7883 18108 9864 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 11057 18139 11115 18145
rect 10244 18108 11008 18136
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 6546 18068 6552 18080
rect 1627 18040 6552 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 7193 18071 7251 18077
rect 7193 18037 7205 18071
rect 7239 18068 7251 18071
rect 9674 18068 9680 18080
rect 7239 18040 9680 18068
rect 7239 18037 7251 18040
rect 7193 18031 7251 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 9769 18071 9827 18077
rect 9769 18037 9781 18071
rect 9815 18068 9827 18071
rect 10244 18068 10272 18108
rect 9815 18040 10272 18068
rect 9815 18037 9827 18040
rect 9769 18031 9827 18037
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 10980 18068 11008 18108
rect 11057 18105 11069 18139
rect 11103 18136 11115 18139
rect 12360 18136 12388 18167
rect 12894 18136 12900 18148
rect 11103 18108 11928 18136
rect 12360 18108 12900 18136
rect 11103 18105 11115 18108
rect 11057 18099 11115 18105
rect 11422 18068 11428 18080
rect 10376 18040 10421 18068
rect 10980 18040 11428 18068
rect 10376 18028 10382 18040
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 11900 18068 11928 18108
rect 12894 18096 12900 18108
rect 12952 18096 12958 18148
rect 13188 18136 13216 18176
rect 13538 18164 13544 18176
rect 13596 18164 13602 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16666 18204 16672 18216
rect 15703 18176 16672 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 16666 18164 16672 18176
rect 16724 18204 16730 18216
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16724 18176 16957 18204
rect 16724 18164 16730 18176
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18173 17279 18207
rect 17221 18167 17279 18173
rect 13188 18108 13492 18136
rect 13354 18068 13360 18080
rect 11900 18040 13360 18068
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 13464 18068 13492 18108
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 16206 18136 16212 18148
rect 14608 18108 16212 18136
rect 14608 18096 14614 18108
rect 16206 18096 16212 18108
rect 16264 18096 16270 18148
rect 16482 18096 16488 18148
rect 16540 18136 16546 18148
rect 17236 18136 17264 18167
rect 17310 18164 17316 18216
rect 17368 18204 17374 18216
rect 17368 18176 19472 18204
rect 17368 18164 17374 18176
rect 16540 18108 17264 18136
rect 19444 18136 19472 18176
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 23109 18207 23167 18213
rect 22152 18176 22197 18204
rect 22152 18164 22158 18176
rect 23109 18173 23121 18207
rect 23155 18204 23167 18207
rect 23290 18204 23296 18216
rect 23155 18176 23296 18204
rect 23155 18173 23167 18176
rect 23109 18167 23167 18173
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 23569 18207 23627 18213
rect 23569 18173 23581 18207
rect 23615 18173 23627 18207
rect 23569 18167 23627 18173
rect 24765 18207 24823 18213
rect 24765 18173 24777 18207
rect 24811 18204 24823 18207
rect 24854 18204 24860 18216
rect 24811 18176 24860 18204
rect 24811 18173 24823 18176
rect 24765 18167 24823 18173
rect 23584 18136 23612 18167
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 25041 18207 25099 18213
rect 25041 18173 25053 18207
rect 25087 18173 25099 18207
rect 25041 18167 25099 18173
rect 25961 18207 26019 18213
rect 25961 18173 25973 18207
rect 26007 18204 26019 18207
rect 26142 18204 26148 18216
rect 26007 18176 26148 18204
rect 26007 18173 26019 18176
rect 25961 18167 26019 18173
rect 25056 18136 25084 18167
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 26602 18204 26608 18216
rect 26563 18176 26608 18204
rect 26602 18164 26608 18176
rect 26660 18164 26666 18216
rect 27798 18136 27804 18148
rect 19444 18108 23612 18136
rect 23676 18108 25084 18136
rect 27759 18108 27804 18136
rect 16540 18096 16546 18108
rect 16758 18068 16764 18080
rect 13464 18040 16764 18068
rect 16758 18028 16764 18040
rect 16816 18028 16822 18080
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 19705 18071 19763 18077
rect 19705 18068 19717 18071
rect 18104 18040 19717 18068
rect 18104 18028 18110 18040
rect 19705 18037 19717 18040
rect 19751 18037 19763 18071
rect 19705 18031 19763 18037
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 20533 18071 20591 18077
rect 20533 18068 20545 18071
rect 20496 18040 20545 18068
rect 20496 18028 20502 18040
rect 20533 18037 20545 18040
rect 20579 18037 20591 18071
rect 20533 18031 20591 18037
rect 23198 18028 23204 18080
rect 23256 18068 23262 18080
rect 23676 18068 23704 18108
rect 27798 18096 27804 18108
rect 27856 18096 27862 18148
rect 23256 18040 23704 18068
rect 24213 18071 24271 18077
rect 23256 18028 23262 18040
rect 24213 18037 24225 18071
rect 24259 18068 24271 18071
rect 26234 18068 26240 18080
rect 24259 18040 26240 18068
rect 24259 18037 24271 18040
rect 24213 18031 24271 18037
rect 26234 18028 26240 18040
rect 26292 18028 26298 18080
rect 28994 18068 29000 18080
rect 28955 18040 29000 18068
rect 28994 18028 29000 18040
rect 29052 18028 29058 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 7561 17867 7619 17873
rect 7561 17864 7573 17867
rect 6788 17836 7573 17864
rect 6788 17824 6794 17836
rect 7561 17833 7573 17836
rect 7607 17864 7619 17867
rect 9398 17864 9404 17876
rect 7607 17836 9404 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 11701 17867 11759 17873
rect 11701 17864 11713 17867
rect 10928 17836 11713 17864
rect 10928 17824 10934 17836
rect 11701 17833 11713 17836
rect 11747 17833 11759 17867
rect 11701 17827 11759 17833
rect 11790 17824 11796 17876
rect 11848 17864 11854 17876
rect 14366 17864 14372 17876
rect 11848 17836 14372 17864
rect 11848 17824 11854 17836
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 14461 17867 14519 17873
rect 14461 17833 14473 17867
rect 14507 17864 14519 17867
rect 15102 17864 15108 17876
rect 14507 17836 15108 17864
rect 14507 17833 14519 17836
rect 14461 17827 14519 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 16206 17824 16212 17876
rect 16264 17864 16270 17876
rect 19426 17864 19432 17876
rect 16264 17836 19432 17864
rect 16264 17824 16270 17836
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22244 17836 22845 17864
rect 22244 17824 22250 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 22833 17827 22891 17833
rect 25593 17867 25651 17873
rect 25593 17833 25605 17867
rect 25639 17864 25651 17867
rect 26050 17864 26056 17876
rect 25639 17836 26056 17864
rect 25639 17833 25651 17836
rect 25593 17827 25651 17833
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 32122 17864 32128 17876
rect 32083 17836 32128 17864
rect 32122 17824 32128 17836
rect 32180 17824 32186 17876
rect 7466 17796 7472 17808
rect 5920 17768 7472 17796
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4614 17728 4620 17740
rect 4387 17700 4620 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5920 17669 5948 17768
rect 7466 17756 7472 17768
rect 7524 17756 7530 17808
rect 8570 17756 8576 17808
rect 8628 17796 8634 17808
rect 10410 17796 10416 17808
rect 8628 17768 10416 17796
rect 8628 17756 8634 17768
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 10686 17756 10692 17808
rect 10744 17796 10750 17808
rect 13262 17796 13268 17808
rect 10744 17768 13268 17796
rect 10744 17756 10750 17768
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 13633 17799 13691 17805
rect 13633 17765 13645 17799
rect 13679 17796 13691 17799
rect 15654 17796 15660 17808
rect 13679 17768 15660 17796
rect 13679 17765 13691 17768
rect 13633 17759 13691 17765
rect 15654 17756 15660 17768
rect 15712 17756 15718 17808
rect 20806 17796 20812 17808
rect 15764 17768 20812 17796
rect 6638 17728 6644 17740
rect 6012 17700 6644 17728
rect 5905 17663 5963 17669
rect 5905 17629 5917 17663
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 1854 17552 1860 17604
rect 1912 17592 1918 17604
rect 6012 17592 6040 17700
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 6880 17700 7389 17728
rect 6880 17688 6886 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 9950 17728 9956 17740
rect 7616 17700 9956 17728
rect 7616 17688 7622 17700
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10318 17728 10324 17740
rect 10231 17700 10324 17728
rect 10318 17688 10324 17700
rect 10376 17728 10382 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 10376 17700 13093 17728
rect 10376 17688 10382 17700
rect 13081 17697 13093 17700
rect 13127 17728 13139 17731
rect 15764 17728 15792 17768
rect 20806 17756 20812 17768
rect 20864 17756 20870 17808
rect 13127 17700 15792 17728
rect 17405 17731 17463 17737
rect 13127 17697 13139 17700
rect 13081 17691 13139 17697
rect 17405 17697 17417 17731
rect 17451 17728 17463 17731
rect 22094 17728 22100 17740
rect 17451 17700 22100 17728
rect 17451 17697 17463 17700
rect 17405 17691 17463 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 24854 17728 24860 17740
rect 24815 17700 24860 17728
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 26234 17728 26240 17740
rect 26195 17700 26240 17728
rect 26234 17688 26240 17700
rect 26292 17688 26298 17740
rect 26881 17731 26939 17737
rect 26881 17697 26893 17731
rect 26927 17728 26939 17731
rect 29086 17728 29092 17740
rect 26927 17700 29092 17728
rect 26927 17697 26939 17700
rect 26881 17691 26939 17697
rect 29086 17688 29092 17700
rect 29144 17688 29150 17740
rect 6546 17660 6552 17672
rect 6507 17632 6552 17660
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 6730 17620 6736 17672
rect 6788 17660 6794 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 6788 17632 7205 17660
rect 6788 17620 6794 17632
rect 7193 17629 7205 17632
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17660 8447 17663
rect 8662 17660 8668 17672
rect 8435 17632 8668 17660
rect 8435 17629 8447 17632
rect 8389 17623 8447 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 11606 17660 11612 17672
rect 10827 17632 11612 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 11606 17620 11612 17632
rect 11664 17620 11670 17672
rect 11885 17663 11943 17669
rect 11885 17629 11897 17663
rect 11931 17660 11943 17663
rect 11974 17660 11980 17672
rect 11931 17632 11980 17660
rect 11931 17629 11943 17632
rect 11885 17623 11943 17629
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12342 17660 12348 17672
rect 12303 17632 12348 17660
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14182 17660 14188 17672
rect 13872 17632 14188 17660
rect 13872 17620 13878 17632
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 14642 17660 14648 17672
rect 14415 17632 14648 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 14642 17620 14648 17632
rect 14700 17620 14706 17672
rect 16209 17663 16267 17669
rect 16209 17629 16221 17663
rect 16255 17660 16267 17663
rect 17126 17660 17132 17672
rect 16255 17632 17132 17660
rect 16255 17629 16267 17632
rect 16209 17623 16267 17629
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 18506 17660 18512 17672
rect 18467 17632 18512 17660
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 19518 17660 19524 17672
rect 19479 17632 19524 17660
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 19610 17620 19616 17672
rect 19668 17660 19674 17672
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 19668 17632 20545 17660
rect 19668 17620 19674 17632
rect 20533 17629 20545 17632
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17660 22799 17663
rect 25501 17663 25559 17669
rect 25501 17660 25513 17663
rect 22787 17632 25513 17660
rect 22787 17629 22799 17632
rect 22741 17623 22799 17629
rect 25501 17629 25513 17632
rect 25547 17660 25559 17663
rect 25774 17660 25780 17672
rect 25547 17632 25780 17660
rect 25547 17629 25559 17632
rect 25501 17623 25559 17629
rect 25774 17620 25780 17632
rect 25832 17620 25838 17672
rect 27706 17660 27712 17672
rect 27667 17632 27712 17660
rect 27706 17620 27712 17632
rect 27764 17620 27770 17672
rect 29178 17620 29184 17672
rect 29236 17660 29242 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29236 17632 29745 17660
rect 29236 17620 29242 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 32309 17663 32367 17669
rect 32309 17629 32321 17663
rect 32355 17660 32367 17663
rect 37274 17660 37280 17672
rect 32355 17632 37280 17660
rect 32355 17629 32367 17632
rect 32309 17623 32367 17629
rect 1912 17564 6040 17592
rect 1912 17552 1918 17564
rect 6086 17552 6092 17604
rect 6144 17592 6150 17604
rect 9677 17595 9735 17601
rect 9677 17592 9689 17595
rect 6144 17564 9689 17592
rect 6144 17552 6150 17564
rect 9677 17561 9689 17564
rect 9723 17561 9735 17595
rect 9677 17555 9735 17561
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 9824 17564 9869 17592
rect 9824 17552 9830 17564
rect 10962 17552 10968 17604
rect 11020 17592 11026 17604
rect 11057 17595 11115 17601
rect 11057 17592 11069 17595
rect 11020 17564 11069 17592
rect 11020 17552 11026 17564
rect 11057 17561 11069 17564
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 13173 17595 13231 17601
rect 13173 17561 13185 17595
rect 13219 17592 13231 17595
rect 13262 17592 13268 17604
rect 13219 17564 13268 17592
rect 13219 17561 13231 17564
rect 13173 17555 13231 17561
rect 13262 17552 13268 17564
rect 13320 17552 13326 17604
rect 15102 17592 15108 17604
rect 15063 17564 15108 17592
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 15197 17595 15255 17601
rect 15197 17561 15209 17595
rect 15243 17561 15255 17595
rect 17494 17592 17500 17604
rect 17455 17564 17500 17592
rect 15197 17555 15255 17561
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5960 17496 6009 17524
rect 5960 17484 5966 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 6641 17527 6699 17533
rect 6641 17493 6653 17527
rect 6687 17524 6699 17527
rect 8386 17524 8392 17536
rect 6687 17496 8392 17524
rect 6687 17493 6699 17496
rect 6641 17487 6699 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 8481 17527 8539 17533
rect 8481 17493 8493 17527
rect 8527 17524 8539 17527
rect 10686 17524 10692 17536
rect 8527 17496 10692 17524
rect 8527 17493 8539 17496
rect 8481 17487 8539 17493
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 12437 17527 12495 17533
rect 12437 17493 12449 17527
rect 12483 17524 12495 17527
rect 12526 17524 12532 17536
rect 12483 17496 12532 17524
rect 12483 17493 12495 17496
rect 12437 17487 12495 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 14826 17484 14832 17536
rect 14884 17524 14890 17536
rect 15212 17524 15240 17555
rect 17494 17552 17500 17564
rect 17552 17552 17558 17604
rect 17586 17552 17592 17604
rect 17644 17592 17650 17604
rect 18049 17595 18107 17601
rect 18049 17592 18061 17595
rect 17644 17564 18061 17592
rect 17644 17552 17650 17564
rect 18049 17561 18061 17564
rect 18095 17592 18107 17595
rect 18230 17592 18236 17604
rect 18095 17564 18236 17592
rect 18095 17561 18107 17564
rect 18049 17555 18107 17561
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 19150 17552 19156 17604
rect 19208 17592 19214 17604
rect 23198 17592 23204 17604
rect 19208 17564 23204 17592
rect 19208 17552 19214 17564
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 26326 17552 26332 17604
rect 26384 17592 26390 17604
rect 26384 17564 26429 17592
rect 26384 17552 26390 17564
rect 27154 17552 27160 17604
rect 27212 17592 27218 17604
rect 32324 17592 32352 17623
rect 37274 17620 37280 17632
rect 37332 17620 37338 17672
rect 27212 17564 32352 17592
rect 27212 17552 27218 17564
rect 14884 17496 15240 17524
rect 16301 17527 16359 17533
rect 14884 17484 14890 17496
rect 16301 17493 16313 17527
rect 16347 17524 16359 17527
rect 16390 17524 16396 17536
rect 16347 17496 16396 17524
rect 16347 17493 16359 17496
rect 16301 17487 16359 17493
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 17402 17484 17408 17536
rect 17460 17524 17466 17536
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 17460 17496 18613 17524
rect 17460 17484 17466 17496
rect 18601 17493 18613 17496
rect 18647 17493 18659 17527
rect 18601 17487 18659 17493
rect 19613 17527 19671 17533
rect 19613 17493 19625 17527
rect 19659 17524 19671 17527
rect 19978 17524 19984 17536
rect 19659 17496 19984 17524
rect 19659 17493 19671 17496
rect 19613 17487 19671 17493
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20622 17524 20628 17536
rect 20583 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 27525 17527 27583 17533
rect 27525 17493 27537 17527
rect 27571 17524 27583 17527
rect 27890 17524 27896 17536
rect 27571 17496 27896 17524
rect 27571 17493 27583 17496
rect 27525 17487 27583 17493
rect 27890 17484 27896 17496
rect 27948 17484 27954 17536
rect 29270 17484 29276 17536
rect 29328 17524 29334 17536
rect 29825 17527 29883 17533
rect 29825 17524 29837 17527
rect 29328 17496 29837 17524
rect 29328 17484 29334 17496
rect 29825 17493 29837 17496
rect 29871 17493 29883 17527
rect 29825 17487 29883 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 8570 17320 8576 17332
rect 6656 17292 8576 17320
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17184 3571 17187
rect 3694 17184 3700 17196
rect 3559 17156 3700 17184
rect 3559 17153 3571 17156
rect 3513 17147 3571 17153
rect 3694 17144 3700 17156
rect 3752 17144 3758 17196
rect 4154 17184 4160 17196
rect 4115 17156 4160 17184
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4982 17184 4988 17196
rect 4943 17156 4988 17184
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 5810 17184 5816 17196
rect 5771 17156 5816 17184
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 6656 17193 6684 17292
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 15102 17320 15108 17332
rect 8772 17292 8984 17320
rect 7190 17212 7196 17264
rect 7248 17252 7254 17264
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 7248 17224 7481 17252
rect 7248 17212 7254 17224
rect 7469 17221 7481 17224
rect 7515 17221 7527 17255
rect 7469 17215 7527 17221
rect 8018 17212 8024 17264
rect 8076 17252 8082 17264
rect 8772 17252 8800 17292
rect 8076 17224 8800 17252
rect 8956 17252 8984 17292
rect 11348 17292 15108 17320
rect 8956 17224 9352 17252
rect 8076 17212 8082 17224
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 8849 17187 8907 17193
rect 8536 17182 8800 17184
rect 8849 17182 8861 17187
rect 8536 17156 8861 17182
rect 8536 17144 8542 17156
rect 8772 17154 8861 17156
rect 8849 17153 8861 17154
rect 8895 17153 8907 17187
rect 9030 17184 9036 17196
rect 8991 17156 9036 17184
rect 8849 17147 8907 17153
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 9324 17184 9352 17224
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 9493 17255 9551 17261
rect 9493 17252 9505 17255
rect 9456 17224 9505 17252
rect 9456 17212 9462 17224
rect 9493 17221 9505 17224
rect 9539 17221 9551 17255
rect 9493 17215 9551 17221
rect 10502 17212 10508 17264
rect 10560 17252 10566 17264
rect 10597 17255 10655 17261
rect 10597 17252 10609 17255
rect 10560 17224 10609 17252
rect 10560 17212 10566 17224
rect 10597 17221 10609 17224
rect 10643 17221 10655 17255
rect 10597 17215 10655 17221
rect 10686 17212 10692 17264
rect 10744 17252 10750 17264
rect 11149 17255 11207 17261
rect 11149 17252 11161 17255
rect 10744 17224 11161 17252
rect 10744 17212 10750 17224
rect 11149 17221 11161 17224
rect 11195 17252 11207 17255
rect 11348 17252 11376 17292
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 19150 17320 19156 17332
rect 17788 17292 19156 17320
rect 11195 17224 11376 17252
rect 11195 17221 11207 17224
rect 11149 17215 11207 17221
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 14369 17255 14427 17261
rect 14369 17252 14381 17255
rect 11480 17224 14381 17252
rect 11480 17212 11486 17224
rect 14369 17221 14381 17224
rect 14415 17221 14427 17255
rect 14369 17215 14427 17221
rect 15749 17255 15807 17261
rect 15749 17221 15761 17255
rect 15795 17252 15807 17255
rect 16298 17252 16304 17264
rect 15795 17224 16304 17252
rect 15795 17221 15807 17224
rect 15749 17215 15807 17221
rect 16298 17212 16304 17224
rect 16356 17212 16362 17264
rect 11974 17184 11980 17196
rect 9324 17156 10364 17184
rect 11935 17156 11980 17184
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 6788 17088 7389 17116
rect 6788 17076 6794 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 10134 17116 10140 17128
rect 7616 17088 10140 17116
rect 7616 17076 7622 17088
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17048 5963 17051
rect 6822 17048 6828 17060
rect 5951 17020 6828 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 6822 17008 6828 17020
rect 6880 17008 6886 17060
rect 7929 17051 7987 17057
rect 7929 17017 7941 17051
rect 7975 17048 7987 17051
rect 10042 17048 10048 17060
rect 7975 17020 10048 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10336 17048 10364 17156
rect 11974 17144 11980 17156
rect 12032 17144 12038 17196
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 13262 17184 13268 17196
rect 13223 17156 13268 17184
rect 12621 17147 12679 17153
rect 10505 17119 10563 17125
rect 10505 17085 10517 17119
rect 10551 17116 10563 17119
rect 11238 17116 11244 17128
rect 10551 17088 11244 17116
rect 10551 17085 10563 17088
rect 10505 17079 10563 17085
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 12636 17116 12664 17147
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 17218 17184 17224 17196
rect 17179 17156 17224 17184
rect 17218 17144 17224 17156
rect 17276 17144 17282 17196
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 11992 17088 13461 17116
rect 11992 17048 12020 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13722 17076 13728 17128
rect 13780 17116 13786 17128
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 13780 17088 14289 17116
rect 13780 17076 13786 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14550 17116 14556 17128
rect 14511 17088 14556 17116
rect 14277 17079 14335 17085
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 15654 17116 15660 17128
rect 15615 17088 15660 17116
rect 15654 17076 15660 17088
rect 15712 17076 15718 17128
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17116 16359 17119
rect 17788 17116 17816 17292
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 22738 17320 22744 17332
rect 20312 17292 22744 17320
rect 20312 17280 20318 17292
rect 22738 17280 22744 17292
rect 22796 17280 22802 17332
rect 25038 17280 25044 17332
rect 25096 17320 25102 17332
rect 25225 17323 25283 17329
rect 25225 17320 25237 17323
rect 25096 17292 25237 17320
rect 25096 17280 25102 17292
rect 25225 17289 25237 17292
rect 25271 17289 25283 17323
rect 25225 17283 25283 17289
rect 18046 17252 18052 17264
rect 18007 17224 18052 17252
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 19242 17252 19248 17264
rect 19203 17224 19248 17252
rect 19242 17212 19248 17224
rect 19300 17212 19306 17264
rect 20438 17252 20444 17264
rect 20399 17224 20444 17252
rect 20438 17212 20444 17224
rect 20496 17212 20502 17264
rect 23382 17252 23388 17264
rect 23343 17224 23388 17252
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 23477 17255 23535 17261
rect 23477 17221 23489 17255
rect 23523 17252 23535 17255
rect 25498 17252 25504 17264
rect 23523 17224 25504 17252
rect 23523 17221 23535 17224
rect 23477 17215 23535 17221
rect 25498 17212 25504 17224
rect 25556 17212 25562 17264
rect 25958 17252 25964 17264
rect 25919 17224 25964 17252
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 26050 17212 26056 17264
rect 26108 17252 26114 17264
rect 27890 17252 27896 17264
rect 26108 17224 26153 17252
rect 27851 17224 27896 17252
rect 26108 17212 26114 17224
rect 27890 17212 27896 17224
rect 27948 17212 27954 17264
rect 28445 17255 28503 17261
rect 28445 17221 28457 17255
rect 28491 17252 28503 17255
rect 29086 17252 29092 17264
rect 28491 17224 29092 17252
rect 28491 17221 28503 17224
rect 28445 17215 28503 17221
rect 29086 17212 29092 17224
rect 29144 17212 29150 17264
rect 24489 17187 24547 17193
rect 24489 17153 24501 17187
rect 24535 17153 24547 17187
rect 24489 17147 24547 17153
rect 16347 17088 17816 17116
rect 17957 17119 18015 17125
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 17957 17085 17969 17119
rect 18003 17116 18015 17119
rect 18966 17116 18972 17128
rect 18003 17088 18972 17116
rect 18003 17085 18015 17088
rect 17957 17079 18015 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17116 19211 17119
rect 19794 17116 19800 17128
rect 19199 17088 19800 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 19794 17076 19800 17088
rect 19852 17116 19858 17128
rect 20349 17119 20407 17125
rect 20349 17116 20361 17119
rect 19852 17088 20361 17116
rect 19852 17076 19858 17088
rect 20349 17085 20361 17088
rect 20395 17085 20407 17119
rect 20349 17079 20407 17085
rect 20993 17119 21051 17125
rect 20993 17085 21005 17119
rect 21039 17116 21051 17119
rect 21266 17116 21272 17128
rect 21039 17088 21272 17116
rect 21039 17085 21051 17088
rect 20993 17079 21051 17085
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24210 17116 24216 17128
rect 24075 17088 24216 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 24210 17076 24216 17088
rect 24268 17076 24274 17128
rect 24504 17116 24532 17147
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 25133 17187 25191 17193
rect 25133 17184 25145 17187
rect 24636 17156 25145 17184
rect 24636 17144 24642 17156
rect 25133 17153 25145 17156
rect 25179 17153 25191 17187
rect 29270 17184 29276 17196
rect 29231 17156 29276 17184
rect 25133 17147 25191 17153
rect 29270 17144 29276 17156
rect 29328 17144 29334 17196
rect 38286 17184 38292 17196
rect 38247 17156 38292 17184
rect 38286 17144 38292 17156
rect 38344 17144 38350 17196
rect 24854 17116 24860 17128
rect 24504 17088 24860 17116
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 26602 17116 26608 17128
rect 26515 17088 26608 17116
rect 26602 17076 26608 17088
rect 26660 17116 26666 17128
rect 27062 17116 27068 17128
rect 26660 17088 27068 17116
rect 26660 17076 26666 17088
rect 27062 17076 27068 17088
rect 27120 17076 27126 17128
rect 27801 17119 27859 17125
rect 27801 17085 27813 17119
rect 27847 17116 27859 17119
rect 29089 17119 29147 17125
rect 27847 17088 28856 17116
rect 27847 17085 27859 17088
rect 27801 17079 27859 17085
rect 10336 17020 12020 17048
rect 12069 17051 12127 17057
rect 12069 17017 12081 17051
rect 12115 17048 12127 17051
rect 12115 17020 13860 17048
rect 12115 17017 12127 17020
rect 12069 17011 12127 17017
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 3605 16983 3663 16989
rect 3605 16980 3617 16983
rect 3384 16952 3617 16980
rect 3384 16940 3390 16952
rect 3605 16949 3617 16952
rect 3651 16949 3663 16983
rect 3605 16943 3663 16949
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 4706 16980 4712 16992
rect 4295 16952 4712 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 4801 16983 4859 16989
rect 4801 16949 4813 16983
rect 4847 16980 4859 16983
rect 5442 16980 5448 16992
rect 4847 16952 5448 16980
rect 4847 16949 4859 16952
rect 4801 16943 4859 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 6733 16983 6791 16989
rect 6733 16949 6745 16983
rect 6779 16980 6791 16983
rect 9950 16980 9956 16992
rect 6779 16952 9956 16980
rect 6779 16949 6791 16952
rect 6733 16943 6791 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 12713 16983 12771 16989
rect 12713 16949 12725 16983
rect 12759 16980 12771 16983
rect 13722 16980 13728 16992
rect 12759 16952 13728 16980
rect 12759 16949 12771 16952
rect 12713 16943 12771 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 13832 16980 13860 17020
rect 15102 17008 15108 17060
rect 15160 17048 15166 17060
rect 18509 17051 18567 17057
rect 18509 17048 18521 17051
rect 15160 17020 18521 17048
rect 15160 17008 15166 17020
rect 18509 17017 18521 17020
rect 18555 17017 18567 17051
rect 18509 17011 18567 17017
rect 19426 17008 19432 17060
rect 19484 17048 19490 17060
rect 19705 17051 19763 17057
rect 19705 17048 19717 17051
rect 19484 17020 19717 17048
rect 19484 17008 19490 17020
rect 19705 17017 19717 17020
rect 19751 17048 19763 17051
rect 20162 17048 20168 17060
rect 19751 17020 20168 17048
rect 19751 17017 19763 17020
rect 19705 17011 19763 17017
rect 20162 17008 20168 17020
rect 20220 17008 20226 17060
rect 28828 17048 28856 17088
rect 29089 17085 29101 17119
rect 29135 17116 29147 17119
rect 29822 17116 29828 17128
rect 29135 17088 29828 17116
rect 29135 17085 29147 17088
rect 29089 17079 29147 17085
rect 29822 17076 29828 17088
rect 29880 17116 29886 17128
rect 30190 17116 30196 17128
rect 29880 17088 30196 17116
rect 29880 17076 29886 17088
rect 30190 17076 30196 17088
rect 30248 17076 30254 17128
rect 28994 17048 29000 17060
rect 28828 17020 29000 17048
rect 28994 17008 29000 17020
rect 29052 17048 29058 17060
rect 29457 17051 29515 17057
rect 29457 17048 29469 17051
rect 29052 17020 29469 17048
rect 29052 17008 29058 17020
rect 29457 17017 29469 17020
rect 29503 17017 29515 17051
rect 29457 17011 29515 17017
rect 15194 16980 15200 16992
rect 13832 16952 15200 16980
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17313 16983 17371 16989
rect 17313 16980 17325 16983
rect 16632 16952 17325 16980
rect 16632 16940 16638 16952
rect 17313 16949 17325 16952
rect 17359 16949 17371 16983
rect 17313 16943 17371 16949
rect 17586 16940 17592 16992
rect 17644 16980 17650 16992
rect 19886 16980 19892 16992
rect 17644 16952 19892 16980
rect 17644 16940 17650 16952
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 22186 16940 22192 16992
rect 22244 16980 22250 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 22244 16952 24593 16980
rect 22244 16940 22250 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 38102 16980 38108 16992
rect 38063 16952 38108 16980
rect 24581 16943 24639 16949
rect 38102 16940 38108 16952
rect 38160 16940 38166 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 5810 16736 5816 16788
rect 5868 16776 5874 16788
rect 7926 16776 7932 16788
rect 5868 16748 7932 16776
rect 5868 16736 5874 16748
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 13262 16776 13268 16788
rect 8404 16748 13268 16776
rect 6362 16708 6368 16720
rect 5184 16680 6368 16708
rect 2682 16532 2688 16584
rect 2740 16572 2746 16584
rect 3237 16575 3295 16581
rect 3237 16572 3249 16575
rect 2740 16544 3249 16572
rect 2740 16532 2746 16544
rect 3237 16541 3249 16544
rect 3283 16541 3295 16575
rect 3237 16535 3295 16541
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16572 4583 16575
rect 4798 16572 4804 16584
rect 4571 16544 4804 16572
rect 4571 16541 4583 16544
rect 4525 16535 4583 16541
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 5184 16581 5212 16680
rect 6362 16668 6368 16680
rect 6420 16668 6426 16720
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 6546 16640 6552 16652
rect 5776 16612 5856 16640
rect 5776 16600 5782 16612
rect 5828 16581 5856 16612
rect 6472 16612 6552 16640
rect 6472 16581 6500 16612
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 7558 16640 7564 16652
rect 7116 16612 7564 16640
rect 7116 16581 7144 16612
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8110 16640 8116 16652
rect 7760 16612 8116 16640
rect 7760 16581 7788 16612
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 5813 16575 5871 16581
rect 5813 16541 5825 16575
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16541 6515 16575
rect 6457 16535 6515 16541
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7745 16575 7803 16581
rect 7745 16541 7757 16575
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16572 7895 16575
rect 8202 16572 8208 16584
rect 7883 16544 8208 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8404 16581 8432 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 13906 16776 13912 16788
rect 13464 16748 13912 16776
rect 8478 16668 8484 16720
rect 8536 16708 8542 16720
rect 10229 16711 10287 16717
rect 8536 16680 9720 16708
rect 8536 16668 8542 16680
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 9398 16640 9404 16652
rect 8628 16612 9404 16640
rect 8628 16600 8634 16612
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9692 16649 9720 16680
rect 10229 16677 10241 16711
rect 10275 16708 10287 16711
rect 10318 16708 10324 16720
rect 10275 16680 10324 16708
rect 10275 16677 10287 16680
rect 10229 16671 10287 16677
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 11330 16668 11336 16720
rect 11388 16708 11394 16720
rect 13464 16717 13492 16748
rect 13906 16736 13912 16748
rect 13964 16776 13970 16788
rect 17586 16776 17592 16788
rect 13964 16748 17592 16776
rect 13964 16736 13970 16748
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 18785 16779 18843 16785
rect 18785 16745 18797 16779
rect 18831 16776 18843 16779
rect 19242 16776 19248 16788
rect 18831 16748 19248 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19794 16776 19800 16788
rect 19755 16748 19800 16776
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 19886 16736 19892 16788
rect 19944 16776 19950 16788
rect 22278 16776 22284 16788
rect 19944 16748 22284 16776
rect 19944 16736 19950 16748
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 26050 16736 26056 16788
rect 26108 16776 26114 16788
rect 26145 16779 26203 16785
rect 26145 16776 26157 16779
rect 26108 16748 26157 16776
rect 26108 16736 26114 16748
rect 26145 16745 26157 16748
rect 26191 16745 26203 16779
rect 26145 16739 26203 16745
rect 13449 16711 13507 16717
rect 11388 16680 12940 16708
rect 11388 16668 11394 16680
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 9723 16612 11008 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16541 8447 16575
rect 8389 16535 8447 16541
rect 10594 16532 10600 16584
rect 10652 16572 10658 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10652 16544 10793 16572
rect 10652 16532 10658 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10980 16572 11008 16612
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11112 16612 11529 16640
rect 11112 16600 11118 16612
rect 11517 16609 11529 16612
rect 11563 16609 11575 16643
rect 11790 16640 11796 16652
rect 11751 16612 11796 16640
rect 11517 16603 11575 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 12912 16649 12940 16680
rect 13449 16677 13461 16711
rect 13495 16677 13507 16711
rect 13449 16671 13507 16677
rect 14366 16668 14372 16720
rect 14424 16708 14430 16720
rect 14424 16680 15148 16708
rect 14424 16668 14430 16680
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16609 12955 16643
rect 14458 16640 14464 16652
rect 12897 16603 12955 16609
rect 14384 16612 14464 16640
rect 11238 16572 11244 16584
rect 10980 16544 11244 16572
rect 10781 16535 10839 16541
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 14384 16581 14412 16612
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 15120 16649 15148 16680
rect 16022 16668 16028 16720
rect 16080 16708 16086 16720
rect 18506 16708 18512 16720
rect 16080 16680 18512 16708
rect 16080 16668 16086 16680
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 16666 16640 16672 16652
rect 15151 16612 16672 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16574 16819 16575
rect 16807 16572 16883 16574
rect 17126 16572 17132 16584
rect 16807 16546 17132 16572
rect 16807 16541 16819 16546
rect 16855 16544 17132 16546
rect 16761 16535 16819 16541
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 17420 16581 17448 16680
rect 18506 16668 18512 16680
rect 18564 16668 18570 16720
rect 18966 16668 18972 16720
rect 19024 16708 19030 16720
rect 21726 16708 21732 16720
rect 19024 16680 21732 16708
rect 19024 16668 19030 16680
rect 21726 16668 21732 16680
rect 21784 16708 21790 16720
rect 29825 16711 29883 16717
rect 29825 16708 29837 16711
rect 21784 16680 29837 16708
rect 21784 16668 21790 16680
rect 29825 16677 29837 16680
rect 29871 16677 29883 16711
rect 29825 16671 29883 16677
rect 20070 16640 20076 16652
rect 19352 16612 20076 16640
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 17586 16532 17592 16584
rect 17644 16572 17650 16584
rect 18233 16575 18291 16581
rect 17644 16544 18184 16572
rect 17644 16532 17650 16544
rect 7193 16507 7251 16513
rect 7193 16473 7205 16507
rect 7239 16504 7251 16507
rect 9398 16504 9404 16516
rect 7239 16476 9404 16504
rect 7239 16473 7251 16476
rect 7193 16467 7251 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 9769 16507 9827 16513
rect 9769 16473 9781 16507
rect 9815 16473 9827 16507
rect 9769 16467 9827 16473
rect 2409 16439 2467 16445
rect 2409 16405 2421 16439
rect 2455 16436 2467 16439
rect 2774 16436 2780 16448
rect 2455 16408 2780 16436
rect 2455 16405 2467 16408
rect 2409 16399 2467 16405
rect 2774 16396 2780 16408
rect 2832 16396 2838 16448
rect 2866 16396 2872 16448
rect 2924 16436 2930 16448
rect 3053 16439 3111 16445
rect 3053 16436 3065 16439
rect 2924 16408 3065 16436
rect 2924 16396 2930 16408
rect 3053 16405 3065 16408
rect 3099 16405 3111 16439
rect 3053 16399 3111 16405
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 3476 16408 4629 16436
rect 3476 16396 3482 16408
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 5132 16408 5273 16436
rect 5132 16396 5138 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16436 5963 16439
rect 6270 16436 6276 16448
rect 5951 16408 6276 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 6549 16439 6607 16445
rect 6549 16405 6561 16439
rect 6595 16436 6607 16439
rect 8294 16436 8300 16448
rect 6595 16408 8300 16436
rect 6595 16405 6607 16408
rect 6549 16399 6607 16405
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8478 16436 8484 16448
rect 8439 16408 8484 16436
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 9122 16396 9128 16448
rect 9180 16436 9186 16448
rect 9784 16436 9812 16467
rect 9858 16464 9864 16516
rect 9916 16504 9922 16516
rect 11609 16507 11667 16513
rect 11609 16504 11621 16507
rect 9916 16476 11621 16504
rect 9916 16464 9922 16476
rect 11609 16473 11621 16476
rect 11655 16473 11667 16507
rect 11609 16467 11667 16473
rect 12710 16464 12716 16516
rect 12768 16504 12774 16516
rect 12989 16507 13047 16513
rect 12989 16504 13001 16507
rect 12768 16476 13001 16504
rect 12768 16464 12774 16476
rect 12989 16473 13001 16476
rect 13035 16473 13047 16507
rect 12989 16467 13047 16473
rect 15197 16507 15255 16513
rect 15197 16473 15209 16507
rect 15243 16504 15255 16507
rect 15562 16504 15568 16516
rect 15243 16476 15568 16504
rect 15243 16473 15255 16476
rect 15197 16467 15255 16473
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 16117 16507 16175 16513
rect 16117 16473 16129 16507
rect 16163 16504 16175 16507
rect 16482 16504 16488 16516
rect 16163 16476 16488 16504
rect 16163 16473 16175 16476
rect 16117 16467 16175 16473
rect 16482 16464 16488 16476
rect 16540 16464 16546 16516
rect 16853 16507 16911 16513
rect 16853 16473 16865 16507
rect 16899 16504 16911 16507
rect 17954 16504 17960 16516
rect 16899 16476 17960 16504
rect 16899 16473 16911 16476
rect 16853 16467 16911 16473
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 10870 16436 10876 16448
rect 9180 16408 9812 16436
rect 10831 16408 10876 16436
rect 9180 16396 9186 16408
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 13262 16436 13268 16448
rect 11756 16408 13268 16436
rect 11756 16396 11762 16408
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 14461 16439 14519 16445
rect 14461 16405 14473 16439
rect 14507 16436 14519 16439
rect 14826 16436 14832 16448
rect 14507 16408 14832 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17497 16439 17555 16445
rect 17497 16436 17509 16439
rect 17092 16408 17509 16436
rect 17092 16396 17098 16408
rect 17497 16405 17509 16408
rect 17543 16405 17555 16439
rect 18046 16436 18052 16448
rect 18007 16408 18052 16436
rect 17497 16399 17555 16405
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 18156 16436 18184 16544
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18690 16572 18696 16584
rect 18651 16544 18696 16572
rect 18233 16535 18291 16541
rect 18248 16504 18276 16535
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19352 16572 19380 16612
rect 19720 16581 19748 16612
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 20530 16640 20536 16652
rect 20491 16612 20536 16640
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 20806 16640 20812 16652
rect 20767 16612 20812 16640
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 38102 16640 38108 16652
rect 20956 16612 26096 16640
rect 20956 16600 20962 16612
rect 18800 16544 19380 16572
rect 19705 16575 19763 16581
rect 18800 16504 18828 16544
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 24596 16581 24624 16612
rect 26068 16581 26096 16612
rect 29748 16612 38108 16640
rect 23477 16575 23535 16581
rect 23477 16572 23489 16575
rect 22704 16544 23489 16572
rect 22704 16532 22710 16544
rect 23477 16541 23489 16544
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 26053 16575 26111 16581
rect 26053 16541 26065 16575
rect 26099 16541 26111 16575
rect 27154 16572 27160 16584
rect 27115 16544 27160 16572
rect 26053 16535 26111 16541
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 29748 16581 29776 16612
rect 38102 16600 38108 16612
rect 38160 16600 38166 16652
rect 29733 16575 29791 16581
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 18248 16476 18828 16504
rect 20622 16464 20628 16516
rect 20680 16504 20686 16516
rect 21726 16504 21732 16516
rect 20680 16476 20725 16504
rect 21687 16476 21732 16504
rect 20680 16464 20686 16476
rect 21726 16464 21732 16476
rect 21784 16464 21790 16516
rect 21821 16507 21879 16513
rect 21821 16473 21833 16507
rect 21867 16504 21879 16507
rect 22186 16504 22192 16516
rect 21867 16476 22192 16504
rect 21867 16473 21879 16476
rect 21821 16467 21879 16473
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 22370 16504 22376 16516
rect 22331 16476 22376 16504
rect 22370 16464 22376 16476
rect 22428 16464 22434 16516
rect 22462 16464 22468 16516
rect 22520 16504 22526 16516
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 22520 16476 24685 16504
rect 22520 16464 22526 16476
rect 24673 16473 24685 16476
rect 24719 16473 24731 16507
rect 24673 16467 24731 16473
rect 22094 16436 22100 16448
rect 18156 16408 22100 16436
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 22830 16436 22836 16448
rect 22791 16408 22836 16436
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 23569 16439 23627 16445
rect 23569 16405 23581 16439
rect 23615 16436 23627 16439
rect 24486 16436 24492 16448
rect 23615 16408 24492 16436
rect 23615 16405 23627 16408
rect 23569 16399 23627 16405
rect 24486 16396 24492 16408
rect 24544 16396 24550 16448
rect 27246 16436 27252 16448
rect 27207 16408 27252 16436
rect 27246 16396 27252 16408
rect 27304 16396 27310 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2682 16232 2688 16244
rect 2643 16204 2688 16232
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 7374 16232 7380 16244
rect 3528 16204 7380 16232
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 3528 16105 3556 16204
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8386 16232 8392 16244
rect 8343 16204 8392 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 8536 16204 13308 16232
rect 8536 16192 8542 16204
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 4709 16167 4767 16173
rect 4709 16164 4721 16167
rect 4120 16136 4721 16164
rect 4120 16124 4126 16136
rect 4709 16133 4721 16136
rect 4755 16133 4767 16167
rect 5442 16164 5448 16176
rect 5403 16136 5448 16164
rect 4709 16127 4767 16133
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 6270 16124 6276 16176
rect 6328 16164 6334 16176
rect 9030 16164 9036 16176
rect 6328 16136 9036 16164
rect 6328 16124 6334 16136
rect 9030 16124 9036 16136
rect 9088 16124 9094 16176
rect 9122 16124 9128 16176
rect 9180 16164 9186 16176
rect 9585 16167 9643 16173
rect 9585 16164 9597 16167
rect 9180 16136 9597 16164
rect 9180 16124 9186 16136
rect 9585 16133 9597 16136
rect 9631 16133 9643 16167
rect 9585 16127 9643 16133
rect 9677 16167 9735 16173
rect 9677 16133 9689 16167
rect 9723 16164 9735 16167
rect 10042 16164 10048 16176
rect 9723 16136 10048 16164
rect 9723 16133 9735 16136
rect 9677 16127 9735 16133
rect 10042 16124 10048 16136
rect 10100 16124 10106 16176
rect 12066 16124 12072 16176
rect 12124 16164 12130 16176
rect 13280 16173 13308 16204
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15746 16232 15752 16244
rect 15344 16204 15752 16232
rect 15344 16192 15350 16204
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 16209 16235 16267 16241
rect 16209 16201 16221 16235
rect 16255 16232 16267 16235
rect 17494 16232 17500 16244
rect 16255 16204 17500 16232
rect 16255 16201 16267 16204
rect 16209 16195 16267 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 23290 16232 23296 16244
rect 22152 16204 23296 16232
rect 22152 16192 22158 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23382 16192 23388 16244
rect 23440 16232 23446 16244
rect 27246 16232 27252 16244
rect 23440 16204 27252 16232
rect 23440 16192 23446 16204
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 13173 16167 13231 16173
rect 13173 16164 13185 16167
rect 12124 16136 13185 16164
rect 12124 16124 12130 16136
rect 13173 16133 13185 16136
rect 13219 16133 13231 16167
rect 13173 16127 13231 16133
rect 13265 16167 13323 16173
rect 13265 16133 13277 16167
rect 13311 16133 13323 16167
rect 13265 16127 13323 16133
rect 15930 16124 15936 16176
rect 15988 16164 15994 16176
rect 17129 16167 17187 16173
rect 17129 16164 17141 16167
rect 15988 16136 17141 16164
rect 15988 16124 15994 16136
rect 17129 16133 17141 16136
rect 17175 16164 17187 16167
rect 19242 16164 19248 16176
rect 17175 16136 19248 16164
rect 17175 16133 17187 16136
rect 17129 16127 17187 16133
rect 19242 16124 19248 16136
rect 19300 16124 19306 16176
rect 20346 16164 20352 16176
rect 20307 16136 20352 16164
rect 20346 16124 20352 16136
rect 20404 16124 20410 16176
rect 20438 16124 20444 16176
rect 20496 16164 20502 16176
rect 20622 16164 20628 16176
rect 20496 16136 20628 16164
rect 20496 16124 20502 16136
rect 20622 16124 20628 16136
rect 20680 16124 20686 16176
rect 22830 16164 22836 16176
rect 22791 16136 22836 16164
rect 22830 16124 22836 16136
rect 22888 16124 22894 16176
rect 22922 16124 22928 16176
rect 22980 16164 22986 16176
rect 24486 16164 24492 16176
rect 22980 16136 23025 16164
rect 24447 16136 24492 16164
rect 22980 16124 22986 16136
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 26050 16164 26056 16176
rect 26011 16136 26056 16164
rect 26050 16124 26056 16136
rect 26108 16124 26114 16176
rect 26605 16167 26663 16173
rect 26605 16133 26617 16167
rect 26651 16164 26663 16167
rect 27798 16164 27804 16176
rect 26651 16136 27804 16164
rect 26651 16133 26663 16136
rect 26605 16127 26663 16133
rect 27798 16124 27804 16136
rect 27856 16124 27862 16176
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 3513 16099 3571 16105
rect 3513 16065 3525 16099
rect 3559 16065 3571 16099
rect 3970 16096 3976 16108
rect 3931 16068 3976 16096
rect 3513 16059 3571 16065
rect 2884 16028 2912 16059
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4614 16096 4620 16108
rect 4575 16068 4620 16096
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 6914 16096 6920 16108
rect 6875 16068 6920 16096
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8202 16096 8208 16108
rect 8163 16068 8208 16096
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 8895 16068 9444 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 3694 16028 3700 16040
rect 2884 16000 3700 16028
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 5350 16028 5356 16040
rect 5311 16000 5356 16028
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5997 16031 6055 16037
rect 5997 15997 6009 16031
rect 6043 16028 6055 16031
rect 6086 16028 6092 16040
rect 6043 16000 6092 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 6086 15988 6092 16000
rect 6144 15988 6150 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 9122 16028 9128 16040
rect 7156 16000 9128 16028
rect 7156 15988 7162 16000
rect 9122 15988 9128 16000
rect 9180 15988 9186 16040
rect 9416 16028 9444 16068
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 12161 16099 12219 16105
rect 10744 16068 11192 16096
rect 10744 16056 10750 16068
rect 9674 16028 9680 16040
rect 9416 16000 9680 16028
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10597 16031 10655 16037
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 11054 16028 11060 16040
rect 10643 16000 11060 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11164 16028 11192 16068
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12434 16096 12440 16108
rect 12207 16068 12440 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12434 16056 12440 16068
rect 12492 16096 12498 16108
rect 15194 16096 15200 16108
rect 12492 16068 13032 16096
rect 15155 16068 15200 16096
rect 12492 16056 12498 16068
rect 12345 16031 12403 16037
rect 12345 16028 12357 16031
rect 11164 16000 12357 16028
rect 12345 15997 12357 16000
rect 12391 15997 12403 16031
rect 13004 16028 13032 16068
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16206 16096 16212 16108
rect 16163 16068 16212 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 17310 16096 17316 16108
rect 16899 16068 17316 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17954 16096 17960 16108
rect 17915 16068 17960 16096
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18288 16068 19073 16096
rect 18288 16056 18294 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 19061 16059 19119 16065
rect 22002 16056 22008 16068
rect 22060 16096 22066 16108
rect 22646 16096 22652 16108
rect 22060 16068 22652 16096
rect 22060 16056 22066 16068
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 38286 16096 38292 16108
rect 25332 16068 25820 16096
rect 38247 16068 38292 16096
rect 13170 16028 13176 16040
rect 13004 16000 13176 16028
rect 12345 15991 12403 15997
rect 13170 15988 13176 16000
rect 13228 15988 13234 16040
rect 14182 16028 14188 16040
rect 14143 16000 14188 16028
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 16028 15071 16031
rect 15059 16000 16988 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 2222 15920 2228 15972
rect 2280 15960 2286 15972
rect 4065 15963 4123 15969
rect 4065 15960 4077 15963
rect 2280 15932 4077 15960
rect 2280 15920 2286 15932
rect 4065 15929 4077 15932
rect 4111 15929 4123 15963
rect 7653 15963 7711 15969
rect 4065 15923 4123 15929
rect 6840 15932 7604 15960
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 3329 15895 3387 15901
rect 3329 15892 3341 15895
rect 3108 15864 3341 15892
rect 3108 15852 3114 15864
rect 3329 15861 3341 15864
rect 3375 15861 3387 15895
rect 3329 15855 3387 15861
rect 4890 15852 4896 15904
rect 4948 15892 4954 15904
rect 6840 15892 6868 15932
rect 7006 15892 7012 15904
rect 4948 15864 6868 15892
rect 6967 15864 7012 15892
rect 4948 15852 4954 15864
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 7576 15892 7604 15932
rect 7653 15929 7665 15963
rect 7699 15960 7711 15963
rect 7699 15932 9674 15960
rect 7699 15929 7711 15932
rect 7653 15923 7711 15929
rect 8570 15892 8576 15904
rect 7576 15864 8576 15892
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 8938 15892 8944 15904
rect 8899 15864 8944 15892
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 9646 15892 9674 15932
rect 9766 15920 9772 15972
rect 9824 15960 9830 15972
rect 15381 15963 15439 15969
rect 15381 15960 15393 15963
rect 9824 15932 15393 15960
rect 9824 15920 9830 15932
rect 15381 15929 15393 15932
rect 15427 15960 15439 15963
rect 16758 15960 16764 15972
rect 15427 15932 16764 15960
rect 15427 15929 15439 15932
rect 15381 15923 15439 15929
rect 16758 15920 16764 15932
rect 16816 15920 16822 15972
rect 16960 15960 16988 16000
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18046 16028 18052 16040
rect 17920 16000 18052 16028
rect 17920 15988 17926 16000
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 18156 16000 20269 16028
rect 17770 15960 17776 15972
rect 16960 15932 17776 15960
rect 17770 15920 17776 15932
rect 17828 15960 17834 15972
rect 18156 15960 18184 16000
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 16028 20959 16031
rect 21266 16028 21272 16040
rect 20947 16000 21272 16028
rect 20947 15997 20959 16000
rect 20901 15991 20959 15997
rect 21266 15988 21272 16000
rect 21324 15988 21330 16040
rect 21358 15988 21364 16040
rect 21416 16028 21422 16040
rect 23106 16028 23112 16040
rect 21416 16000 23112 16028
rect 21416 15988 21422 16000
rect 23106 15988 23112 16000
rect 23164 15988 23170 16040
rect 24394 16028 24400 16040
rect 24355 16000 24400 16028
rect 24394 15988 24400 16000
rect 24452 15988 24458 16040
rect 17828 15932 18184 15960
rect 17828 15920 17834 15932
rect 18966 15920 18972 15972
rect 19024 15960 19030 15972
rect 22097 15963 22155 15969
rect 22097 15960 22109 15963
rect 19024 15932 22109 15960
rect 19024 15920 19030 15932
rect 22097 15929 22109 15932
rect 22143 15929 22155 15963
rect 22097 15923 22155 15929
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 25332 15960 25360 16068
rect 25409 16031 25467 16037
rect 25409 15997 25421 16031
rect 25455 15997 25467 16031
rect 25409 15991 25467 15997
rect 23440 15932 25360 15960
rect 23440 15920 23446 15932
rect 12158 15892 12164 15904
rect 9646 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13630 15892 13636 15904
rect 12860 15864 13636 15892
rect 12860 15852 12866 15864
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 17586 15892 17592 15904
rect 14240 15864 17592 15892
rect 14240 15852 14246 15864
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 17920 15864 18061 15892
rect 17920 15852 17926 15864
rect 18049 15861 18061 15864
rect 18095 15861 18107 15895
rect 18049 15855 18107 15861
rect 19153 15895 19211 15901
rect 19153 15861 19165 15895
rect 19199 15892 19211 15895
rect 19426 15892 19432 15904
rect 19199 15864 19432 15892
rect 19199 15861 19211 15864
rect 19153 15855 19211 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 22370 15852 22376 15904
rect 22428 15892 22434 15904
rect 24118 15892 24124 15904
rect 22428 15864 24124 15892
rect 22428 15852 22434 15864
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 25424 15892 25452 15991
rect 25792 15960 25820 16068
rect 38286 16056 38292 16068
rect 38344 16056 38350 16108
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 16028 26019 16031
rect 26142 16028 26148 16040
rect 26007 16000 26148 16028
rect 26007 15997 26019 16000
rect 25961 15991 26019 15997
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 29638 15960 29644 15972
rect 25792 15932 29644 15960
rect 29638 15920 29644 15932
rect 29696 15920 29702 15972
rect 25958 15892 25964 15904
rect 25424 15864 25964 15892
rect 25958 15852 25964 15864
rect 26016 15852 26022 15904
rect 28994 15852 29000 15904
rect 29052 15892 29058 15904
rect 38105 15895 38163 15901
rect 38105 15892 38117 15895
rect 29052 15864 38117 15892
rect 29052 15852 29058 15864
rect 38105 15861 38117 15864
rect 38151 15861 38163 15895
rect 38105 15855 38163 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 4982 15688 4988 15700
rect 1995 15660 4988 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 4982 15648 4988 15660
rect 5040 15648 5046 15700
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 9858 15688 9864 15700
rect 7064 15660 9864 15688
rect 7064 15648 7070 15660
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 15654 15688 15660 15700
rect 11112 15660 12388 15688
rect 11112 15648 11118 15660
rect 12360 15632 12388 15660
rect 13188 15660 15660 15688
rect 3970 15580 3976 15632
rect 4028 15620 4034 15632
rect 7282 15620 7288 15632
rect 4028 15592 7288 15620
rect 4028 15580 4034 15592
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 7558 15580 7564 15632
rect 7616 15620 7622 15632
rect 9122 15620 9128 15632
rect 7616 15592 9128 15620
rect 7616 15580 7622 15592
rect 9122 15580 9128 15592
rect 9180 15580 9186 15632
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 10686 15620 10692 15632
rect 9548 15592 10692 15620
rect 9548 15580 9554 15592
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 10870 15580 10876 15632
rect 10928 15620 10934 15632
rect 10928 15592 12296 15620
rect 10928 15580 10934 15592
rect 2130 15484 2136 15496
rect 2091 15456 2136 15484
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 2682 15444 2688 15496
rect 2740 15484 2746 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 2740 15456 3249 15484
rect 2740 15444 2746 15456
rect 3237 15453 3249 15456
rect 3283 15484 3295 15487
rect 3988 15484 4016 15580
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 6454 15552 6460 15564
rect 4672 15524 5672 15552
rect 6415 15524 6460 15552
rect 4672 15512 4678 15524
rect 4246 15484 4252 15496
rect 3283 15456 4016 15484
rect 4159 15456 4252 15484
rect 3283 15453 3295 15456
rect 3237 15447 3295 15453
rect 4246 15444 4252 15456
rect 4304 15484 4310 15496
rect 4798 15484 4804 15496
rect 4304 15456 4804 15484
rect 4304 15444 4310 15456
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 2593 15419 2651 15425
rect 2593 15385 2605 15419
rect 2639 15416 2651 15419
rect 4985 15419 5043 15425
rect 4985 15416 4997 15419
rect 2639 15388 4997 15416
rect 2639 15385 2651 15388
rect 2593 15379 2651 15385
rect 4985 15385 4997 15388
rect 5031 15385 5043 15419
rect 4985 15379 5043 15385
rect 5074 15376 5080 15428
rect 5132 15416 5138 15428
rect 5644 15425 5672 15524
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 7760 15524 11008 15552
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15484 6331 15487
rect 7098 15484 7104 15496
rect 6319 15456 7104 15484
rect 6319 15453 6331 15456
rect 6273 15447 6331 15453
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 7760 15493 7788 15524
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8570 15484 8576 15496
rect 8435 15456 8576 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 5629 15419 5687 15425
rect 5132 15388 5177 15416
rect 5132 15376 5138 15388
rect 5629 15385 5641 15419
rect 5675 15416 5687 15419
rect 7374 15416 7380 15428
rect 5675 15388 7380 15416
rect 5675 15385 5687 15388
rect 5629 15379 5687 15385
rect 7374 15376 7380 15388
rect 7432 15376 7438 15428
rect 7834 15416 7840 15428
rect 7795 15388 7840 15416
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 9766 15416 9772 15428
rect 8404 15388 9628 15416
rect 9727 15388 9772 15416
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 3329 15351 3387 15357
rect 3329 15348 3341 15351
rect 3292 15320 3341 15348
rect 3292 15308 3298 15320
rect 3329 15317 3341 15320
rect 3375 15317 3387 15351
rect 4338 15348 4344 15360
rect 4299 15320 4344 15348
rect 3329 15311 3387 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 7006 15348 7012 15360
rect 6963 15320 7012 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 7006 15308 7012 15320
rect 7064 15348 7070 15360
rect 8404 15348 8432 15388
rect 7064 15320 8432 15348
rect 7064 15308 7070 15320
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 9600 15348 9628 15388
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 9861 15419 9919 15425
rect 9861 15385 9873 15419
rect 9907 15416 9919 15419
rect 9950 15416 9956 15428
rect 9907 15388 9956 15416
rect 9907 15385 9919 15388
rect 9861 15379 9919 15385
rect 9950 15376 9956 15388
rect 10008 15376 10014 15428
rect 10413 15419 10471 15425
rect 10413 15416 10425 15419
rect 10336 15388 10425 15416
rect 10336 15360 10364 15388
rect 10413 15385 10425 15388
rect 10459 15385 10471 15419
rect 10980 15416 11008 15524
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 12069 15555 12127 15561
rect 12069 15552 12081 15555
rect 11940 15524 12081 15552
rect 11940 15512 11946 15524
rect 12069 15521 12081 15524
rect 12115 15521 12127 15555
rect 12268 15552 12296 15592
rect 12342 15580 12348 15632
rect 12400 15620 12406 15632
rect 13188 15620 13216 15660
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 16758 15688 16764 15700
rect 16719 15660 16764 15688
rect 16758 15648 16764 15660
rect 16816 15648 16822 15700
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 20809 15691 20867 15697
rect 20809 15688 20821 15691
rect 18840 15660 20821 15688
rect 18840 15648 18846 15660
rect 20809 15657 20821 15660
rect 20855 15657 20867 15691
rect 20809 15651 20867 15657
rect 21637 15691 21695 15697
rect 21637 15657 21649 15691
rect 21683 15688 21695 15691
rect 22922 15688 22928 15700
rect 21683 15660 22928 15688
rect 21683 15657 21695 15660
rect 21637 15651 21695 15657
rect 22922 15648 22928 15660
rect 22980 15648 22986 15700
rect 23014 15648 23020 15700
rect 23072 15688 23078 15700
rect 24394 15688 24400 15700
rect 23072 15660 24400 15688
rect 23072 15648 23078 15660
rect 24394 15648 24400 15660
rect 24452 15688 24458 15700
rect 29089 15691 29147 15697
rect 29089 15688 29101 15691
rect 24452 15660 29101 15688
rect 24452 15648 24458 15660
rect 29089 15657 29101 15660
rect 29135 15657 29147 15691
rect 29089 15651 29147 15657
rect 12400 15592 13216 15620
rect 12400 15580 12406 15592
rect 13081 15555 13139 15561
rect 12268 15524 13032 15552
rect 12069 15515 12127 15521
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15484 11115 15487
rect 11606 15484 11612 15496
rect 11103 15456 11612 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 11333 15419 11391 15425
rect 11333 15416 11345 15419
rect 10980 15388 11345 15416
rect 10413 15379 10471 15385
rect 11333 15385 11345 15388
rect 11379 15416 11391 15419
rect 11422 15416 11428 15428
rect 11379 15388 11428 15416
rect 11379 15385 11391 15388
rect 11333 15379 11391 15385
rect 11422 15376 11428 15388
rect 11480 15376 11486 15428
rect 12158 15376 12164 15428
rect 12216 15416 12222 15428
rect 13004 15416 13032 15524
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13188 15552 13216 15592
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 15562 15620 15568 15632
rect 13780 15592 15568 15620
rect 13780 15580 13786 15592
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 18325 15623 18383 15629
rect 18325 15589 18337 15623
rect 18371 15620 18383 15623
rect 22370 15620 22376 15632
rect 18371 15592 22376 15620
rect 18371 15589 18383 15592
rect 18325 15583 18383 15589
rect 22370 15580 22376 15592
rect 22428 15580 22434 15632
rect 23106 15580 23112 15632
rect 23164 15620 23170 15632
rect 23164 15592 30144 15620
rect 23164 15580 23170 15592
rect 13127 15524 13216 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 13320 15524 14933 15552
rect 13320 15512 13326 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 15378 15552 15384 15564
rect 15339 15524 15384 15552
rect 14921 15515 14979 15521
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 16390 15552 16396 15564
rect 16351 15524 16396 15552
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 16850 15552 16856 15564
rect 16623 15524 16856 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 16850 15512 16856 15524
rect 16908 15512 16914 15564
rect 17773 15555 17831 15561
rect 17773 15521 17785 15555
rect 17819 15552 17831 15555
rect 18138 15552 18144 15564
rect 17819 15524 18144 15552
rect 17819 15521 17831 15524
rect 17773 15515 17831 15521
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 19613 15555 19671 15561
rect 19613 15521 19625 15555
rect 19659 15552 19671 15555
rect 20898 15552 20904 15564
rect 19659 15524 20904 15552
rect 19659 15521 19671 15524
rect 19613 15515 19671 15521
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 22738 15552 22744 15564
rect 22699 15524 22744 15552
rect 22738 15512 22744 15524
rect 22796 15512 22802 15564
rect 23658 15512 23664 15564
rect 23716 15552 23722 15564
rect 29822 15552 29828 15564
rect 23716 15524 24624 15552
rect 29783 15524 29828 15552
rect 23716 15512 23722 15524
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14274 15484 14280 15496
rect 13587 15456 14280 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15484 20315 15487
rect 20438 15484 20444 15496
rect 20303 15456 20444 15484
rect 20303 15453 20315 15456
rect 20257 15447 20315 15453
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 20714 15484 20720 15496
rect 20675 15456 20720 15484
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 15013 15419 15071 15425
rect 15013 15416 15025 15419
rect 12216 15388 12261 15416
rect 13004 15388 15025 15416
rect 12216 15376 12222 15388
rect 15013 15385 15025 15388
rect 15059 15385 15071 15419
rect 15013 15379 15071 15385
rect 17862 15376 17868 15428
rect 17920 15416 17926 15428
rect 19705 15419 19763 15425
rect 17920 15388 17965 15416
rect 17920 15376 17926 15388
rect 19705 15385 19717 15419
rect 19751 15416 19763 15419
rect 19978 15416 19984 15428
rect 19751 15388 19984 15416
rect 19751 15385 19763 15388
rect 19705 15379 19763 15385
rect 19978 15376 19984 15388
rect 20036 15376 20042 15428
rect 21560 15416 21588 15447
rect 23382 15444 23388 15496
rect 23440 15484 23446 15496
rect 23842 15484 23848 15496
rect 23440 15456 23485 15484
rect 23803 15456 23848 15484
rect 23440 15444 23446 15456
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 24596 15493 24624 15524
rect 29822 15512 29828 15524
rect 29880 15512 29886 15564
rect 30116 15561 30144 15592
rect 30101 15555 30159 15561
rect 30101 15521 30113 15555
rect 30147 15552 30159 15555
rect 36354 15552 36360 15564
rect 30147 15524 36360 15552
rect 30147 15521 30159 15524
rect 30101 15515 30159 15521
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 37734 15552 37740 15564
rect 37695 15524 37740 15552
rect 37734 15512 37740 15524
rect 37792 15512 37798 15564
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 24762 15484 24768 15496
rect 24627 15456 24768 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 24854 15444 24860 15496
rect 24912 15484 24918 15496
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 24912 15456 25237 15484
rect 24912 15444 24918 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 28994 15484 29000 15496
rect 28955 15456 29000 15484
rect 25225 15447 25283 15453
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 37182 15444 37188 15496
rect 37240 15484 37246 15496
rect 37461 15487 37519 15493
rect 37461 15484 37473 15487
rect 37240 15456 37473 15484
rect 37240 15444 37246 15456
rect 37461 15453 37473 15456
rect 37507 15453 37519 15487
rect 37461 15447 37519 15453
rect 20364 15388 21588 15416
rect 22833 15419 22891 15425
rect 10042 15348 10048 15360
rect 8536 15320 8581 15348
rect 9600 15320 10048 15348
rect 8536 15308 8542 15320
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 10318 15308 10324 15360
rect 10376 15308 10382 15360
rect 13630 15348 13636 15360
rect 13591 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 20364 15348 20392 15388
rect 22833 15385 22845 15419
rect 22879 15385 22891 15419
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 22833 15379 22891 15385
rect 23492 15388 24685 15416
rect 20128 15320 20392 15348
rect 22848 15348 22876 15379
rect 23492 15348 23520 15388
rect 24673 15385 24685 15388
rect 24719 15385 24731 15419
rect 29914 15416 29920 15428
rect 29875 15388 29920 15416
rect 24673 15379 24731 15385
rect 29914 15376 29920 15388
rect 29972 15376 29978 15428
rect 23934 15348 23940 15360
rect 22848 15320 23520 15348
rect 23895 15320 23940 15348
rect 20128 15308 20134 15320
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24026 15308 24032 15360
rect 24084 15348 24090 15360
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 24084 15320 25329 15348
rect 24084 15308 24090 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 25317 15311 25375 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2041 15147 2099 15153
rect 2041 15113 2053 15147
rect 2087 15144 2099 15147
rect 9490 15144 9496 15156
rect 2087 15116 6868 15144
rect 2087 15113 2099 15116
rect 2041 15107 2099 15113
rect 4246 15076 4252 15088
rect 2608 15048 4252 15076
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2406 15008 2412 15020
rect 1995 14980 2412 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2406 14968 2412 14980
rect 2464 14968 2470 15020
rect 2608 15017 2636 15048
rect 4246 15036 4252 15048
rect 4304 15036 4310 15088
rect 6270 15076 6276 15088
rect 4540 15048 6276 15076
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 15008 3295 15011
rect 3786 15008 3792 15020
rect 3283 14980 3792 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 3786 14968 3792 14980
rect 3844 15008 3850 15020
rect 4540 15017 4568 15048
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 3844 14980 3893 15008
rect 3844 14968 3850 14980
rect 3881 14977 3893 14980
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 14977 5227 15011
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 5169 14971 5227 14977
rect 3602 14900 3608 14952
rect 3660 14940 3666 14952
rect 5184 14940 5212 14971
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 3660 14912 5212 14940
rect 3660 14900 3666 14912
rect 3973 14875 4031 14881
rect 3973 14841 3985 14875
rect 4019 14872 4031 14875
rect 4982 14872 4988 14884
rect 4019 14844 4988 14872
rect 4019 14841 4031 14844
rect 3973 14835 4031 14841
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 6840 14872 6868 15116
rect 8220 15116 9496 15144
rect 7282 15036 7288 15088
rect 7340 15076 7346 15088
rect 8018 15076 8024 15088
rect 7340 15048 8024 15076
rect 7340 15036 7346 15048
rect 8018 15036 8024 15048
rect 8076 15036 8082 15088
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 6963 14980 7573 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7561 14977 7573 14980
rect 7607 15008 7619 15011
rect 7834 15008 7840 15020
rect 7607 14980 7840 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 7834 14968 7840 14980
rect 7892 15008 7898 15020
rect 8220 15017 8248 15116
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 9631 15116 15332 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 8294 15036 8300 15088
rect 8352 15076 8358 15088
rect 10321 15079 10379 15085
rect 10321 15076 10333 15079
rect 8352 15048 10333 15076
rect 8352 15036 8358 15048
rect 10321 15045 10333 15048
rect 10367 15045 10379 15079
rect 12434 15076 12440 15088
rect 10321 15039 10379 15045
rect 12268 15048 12440 15076
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7892 14980 8217 15008
rect 7892 14968 7898 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 8938 15008 8944 15020
rect 8895 14980 8944 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 9490 15008 9496 15020
rect 9451 14980 9496 15008
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 12268 15017 12296 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 12529 15079 12587 15085
rect 12529 15045 12541 15079
rect 12575 15076 12587 15079
rect 12986 15076 12992 15088
rect 12575 15048 12992 15076
rect 12575 15045 12587 15048
rect 12529 15039 12587 15045
rect 12986 15036 12992 15048
rect 13044 15036 13050 15088
rect 13354 15076 13360 15088
rect 13315 15048 13360 15076
rect 13354 15036 13360 15048
rect 13412 15036 13418 15088
rect 13906 15076 13912 15088
rect 13867 15048 13912 15076
rect 13906 15036 13912 15048
rect 13964 15036 13970 15088
rect 15304 15085 15332 15116
rect 15654 15104 15660 15156
rect 15712 15144 15718 15156
rect 15712 15116 19334 15144
rect 15712 15104 15718 15116
rect 15289 15079 15347 15085
rect 15289 15045 15301 15079
rect 15335 15045 15347 15079
rect 17402 15076 17408 15088
rect 17363 15048 17408 15076
rect 15289 15039 15347 15045
rect 17402 15036 17408 15048
rect 17460 15036 17466 15088
rect 18598 15076 18604 15088
rect 18559 15048 18604 15076
rect 18598 15036 18604 15048
rect 18656 15036 18662 15088
rect 19306 15076 19334 15116
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 20162 15144 20168 15156
rect 19576 15116 20168 15144
rect 19576 15104 19582 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20254 15104 20260 15156
rect 20312 15104 20318 15156
rect 23566 15144 23572 15156
rect 20916 15116 23572 15144
rect 20272 15076 20300 15104
rect 19306 15048 20300 15076
rect 12253 15011 12311 15017
rect 11296 14980 12204 15008
rect 11296 14968 11302 14980
rect 7374 14900 7380 14952
rect 7432 14940 7438 14952
rect 10229 14943 10287 14949
rect 7432 14928 9168 14940
rect 9324 14928 9628 14940
rect 7432 14912 9628 14928
rect 7432 14900 7438 14912
rect 9140 14900 9352 14912
rect 8386 14872 8392 14884
rect 6840 14844 8392 14872
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 8941 14875 8999 14881
rect 8941 14841 8953 14875
rect 8987 14872 8999 14875
rect 9600 14872 9628 14912
rect 10229 14909 10241 14943
rect 10275 14940 10287 14943
rect 11790 14940 11796 14952
rect 10275 14912 11796 14940
rect 10275 14909 10287 14912
rect 10229 14903 10287 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 12176 14940 12204 14980
rect 12253 14977 12265 15011
rect 12299 14977 12311 15011
rect 14369 15011 14427 15017
rect 12253 14971 12311 14977
rect 12406 14980 12848 15008
rect 12406 14940 12434 14980
rect 12176 14912 12434 14940
rect 12820 14940 12848 14980
rect 14369 14977 14381 15011
rect 14415 14977 14427 15011
rect 16390 15008 16396 15020
rect 14369 14971 14427 14977
rect 16040 14980 16396 15008
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 12820 14912 13277 14940
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 13354 14900 13360 14952
rect 13412 14940 13418 14952
rect 14384 14940 14412 14971
rect 13412 14912 14412 14940
rect 15197 14943 15255 14949
rect 13412 14900 13418 14912
rect 15197 14909 15209 14943
rect 15243 14940 15255 14943
rect 16040 14940 16068 14980
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19300 14980 19625 15008
rect 19300 14968 19306 14980
rect 19613 14977 19625 14980
rect 19659 15008 19671 15011
rect 19794 15008 19800 15020
rect 19659 14980 19800 15008
rect 19659 14977 19671 14980
rect 19613 14971 19671 14977
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20438 15008 20444 15020
rect 20303 14980 20444 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 20916 15017 20944 15116
rect 23566 15104 23572 15116
rect 23624 15104 23630 15156
rect 26234 15144 26240 15156
rect 23676 15116 26240 15144
rect 20993 15079 21051 15085
rect 20993 15045 21005 15079
rect 21039 15076 21051 15079
rect 21174 15076 21180 15088
rect 21039 15048 21180 15076
rect 21039 15045 21051 15048
rect 20993 15039 21051 15045
rect 21174 15036 21180 15048
rect 21232 15036 21238 15088
rect 22189 15079 22247 15085
rect 22189 15045 22201 15079
rect 22235 15076 22247 15079
rect 22462 15076 22468 15088
rect 22235 15048 22468 15076
rect 22235 15045 22247 15048
rect 22189 15039 22247 15045
rect 22462 15036 22468 15048
rect 22520 15036 22526 15088
rect 23676 15085 23704 15116
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 27525 15147 27583 15153
rect 27525 15113 27537 15147
rect 27571 15144 27583 15147
rect 27614 15144 27620 15156
rect 27571 15116 27620 15144
rect 27571 15113 27583 15116
rect 27525 15107 27583 15113
rect 27614 15104 27620 15116
rect 27672 15104 27678 15156
rect 28077 15147 28135 15153
rect 28077 15113 28089 15147
rect 28123 15113 28135 15147
rect 28077 15107 28135 15113
rect 23661 15079 23719 15085
rect 23661 15045 23673 15079
rect 23707 15045 23719 15079
rect 23661 15039 23719 15045
rect 23753 15079 23811 15085
rect 23753 15045 23765 15079
rect 23799 15076 23811 15079
rect 24026 15076 24032 15088
rect 23799 15048 24032 15076
rect 23799 15045 23811 15048
rect 23753 15039 23811 15045
rect 24026 15036 24032 15048
rect 24084 15036 24090 15088
rect 24762 15036 24768 15088
rect 24820 15036 24826 15088
rect 28092 15076 28120 15107
rect 28092 15048 28948 15076
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 14977 20959 15011
rect 24780 15008 24808 15036
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 24780 14980 26249 15008
rect 20901 14971 20959 14977
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 27433 15011 27491 15017
rect 27433 14977 27445 15011
rect 27479 14977 27491 15011
rect 28258 15008 28264 15020
rect 28219 14980 28264 15008
rect 27433 14971 27491 14977
rect 15243 14912 16068 14940
rect 16209 14943 16267 14949
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16482 14940 16488 14952
rect 16255 14912 16488 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16666 14900 16672 14952
rect 16724 14940 16730 14952
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 16724 14912 17325 14940
rect 16724 14900 16730 14912
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17586 14940 17592 14952
rect 17547 14912 17592 14940
rect 17313 14903 17371 14909
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 17736 14912 18521 14940
rect 17736 14900 17742 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 19150 14940 19156 14952
rect 19063 14912 19156 14940
rect 18509 14903 18567 14909
rect 19150 14900 19156 14912
rect 19208 14940 19214 14952
rect 21910 14940 21916 14952
rect 19208 14912 21916 14940
rect 19208 14900 19214 14912
rect 21910 14900 21916 14912
rect 21968 14900 21974 14952
rect 22097 14943 22155 14949
rect 22097 14909 22109 14943
rect 22143 14940 22155 14943
rect 23014 14940 23020 14952
rect 22143 14912 23020 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 23014 14900 23020 14912
rect 23072 14900 23078 14952
rect 23109 14943 23167 14949
rect 23109 14909 23121 14943
rect 23155 14940 23167 14943
rect 23290 14940 23296 14952
rect 23155 14912 23296 14940
rect 23155 14909 23167 14912
rect 23109 14903 23167 14909
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23937 14943 23995 14949
rect 23937 14909 23949 14943
rect 23983 14909 23995 14943
rect 23937 14903 23995 14909
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 8987 14844 9536 14872
rect 9600 14844 10793 14872
rect 8987 14841 8999 14844
rect 8941 14835 8999 14841
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2648 14776 2697 14804
rect 2648 14764 2654 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 2685 14767 2743 14773
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3329 14807 3387 14813
rect 3329 14804 3341 14807
rect 3016 14776 3341 14804
rect 3016 14764 3022 14776
rect 3329 14773 3341 14776
rect 3375 14773 3387 14807
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 3329 14767 3387 14773
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 5261 14807 5319 14813
rect 5261 14773 5273 14807
rect 5307 14804 5319 14807
rect 5626 14804 5632 14816
rect 5307 14776 5632 14804
rect 5307 14773 5319 14776
rect 5261 14767 5319 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 5905 14807 5963 14813
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 6914 14804 6920 14816
rect 5951 14776 6920 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7009 14807 7067 14813
rect 7009 14773 7021 14807
rect 7055 14804 7067 14807
rect 7098 14804 7104 14816
rect 7055 14776 7104 14804
rect 7055 14773 7067 14776
rect 7009 14767 7067 14773
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 8202 14804 8208 14816
rect 7699 14776 8208 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8297 14807 8355 14813
rect 8297 14773 8309 14807
rect 8343 14804 8355 14807
rect 9398 14804 9404 14816
rect 8343 14776 9404 14804
rect 8343 14773 8355 14776
rect 8297 14767 8355 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 9508 14804 9536 14844
rect 10781 14841 10793 14844
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 12986 14832 12992 14884
rect 13044 14872 13050 14884
rect 20162 14872 20168 14884
rect 13044 14844 20168 14872
rect 13044 14832 13050 14844
rect 20162 14832 20168 14844
rect 20220 14832 20226 14884
rect 20349 14875 20407 14881
rect 20349 14841 20361 14875
rect 20395 14872 20407 14875
rect 20395 14844 21220 14872
rect 20395 14841 20407 14844
rect 20349 14835 20407 14841
rect 12710 14804 12716 14816
rect 9508 14776 12716 14804
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13998 14804 14004 14816
rect 12860 14776 14004 14804
rect 12860 14764 12866 14776
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 14550 14764 14556 14776
rect 14608 14804 14614 14816
rect 16850 14804 16856 14816
rect 14608 14776 16856 14804
rect 14608 14764 14614 14776
rect 16850 14764 16856 14776
rect 16908 14804 16914 14816
rect 17310 14804 17316 14816
rect 16908 14776 17316 14804
rect 16908 14764 16914 14776
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 19705 14807 19763 14813
rect 19705 14804 19717 14807
rect 17736 14776 19717 14804
rect 17736 14764 17742 14776
rect 19705 14773 19717 14776
rect 19751 14773 19763 14807
rect 19705 14767 19763 14773
rect 19794 14764 19800 14816
rect 19852 14804 19858 14816
rect 21082 14804 21088 14816
rect 19852 14776 21088 14804
rect 19852 14764 19858 14776
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 21192 14804 21220 14844
rect 21266 14832 21272 14884
rect 21324 14872 21330 14884
rect 22370 14872 22376 14884
rect 21324 14844 22376 14872
rect 21324 14832 21330 14844
rect 22370 14832 22376 14844
rect 22428 14872 22434 14884
rect 23952 14872 23980 14903
rect 24670 14900 24676 14952
rect 24728 14940 24734 14952
rect 27448 14940 27476 14971
rect 28258 14968 28264 14980
rect 28316 14968 28322 15020
rect 28920 15017 28948 15048
rect 28905 15011 28963 15017
rect 28905 14977 28917 15011
rect 28951 14977 28963 15011
rect 38010 15008 38016 15020
rect 37971 14980 38016 15008
rect 28905 14971 28963 14977
rect 38010 14968 38016 14980
rect 38068 14968 38074 15020
rect 28350 14940 28356 14952
rect 24728 14912 28356 14940
rect 24728 14900 24734 14912
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 30006 14900 30012 14952
rect 30064 14940 30070 14952
rect 30101 14943 30159 14949
rect 30101 14940 30113 14943
rect 30064 14912 30113 14940
rect 30064 14900 30070 14912
rect 30101 14909 30113 14912
rect 30147 14909 30159 14943
rect 30101 14903 30159 14909
rect 22428 14844 23980 14872
rect 22428 14832 22434 14844
rect 22738 14804 22744 14816
rect 21192 14776 22744 14804
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 26053 14807 26111 14813
rect 26053 14773 26065 14807
rect 26099 14804 26111 14807
rect 27246 14804 27252 14816
rect 26099 14776 27252 14804
rect 26099 14773 26111 14776
rect 26053 14767 26111 14773
rect 27246 14764 27252 14776
rect 27304 14764 27310 14816
rect 28721 14807 28779 14813
rect 28721 14773 28733 14807
rect 28767 14804 28779 14807
rect 30190 14804 30196 14816
rect 28767 14776 30196 14804
rect 28767 14773 28779 14776
rect 28721 14767 28779 14773
rect 30190 14764 30196 14776
rect 30248 14764 30254 14816
rect 37829 14807 37887 14813
rect 37829 14773 37841 14807
rect 37875 14804 37887 14807
rect 37918 14804 37924 14816
rect 37875 14776 37924 14804
rect 37875 14773 37887 14776
rect 37829 14767 37887 14773
rect 37918 14764 37924 14776
rect 37976 14764 37982 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 8478 14600 8484 14612
rect 4580 14572 8484 14600
rect 4580 14560 4586 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14569 9551 14603
rect 9493 14563 9551 14569
rect 6914 14492 6920 14544
rect 6972 14532 6978 14544
rect 8386 14532 8392 14544
rect 6972 14504 8392 14532
rect 6972 14492 6978 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 4433 14467 4491 14473
rect 2832 14436 2877 14464
rect 2832 14424 2838 14436
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4614 14464 4620 14476
rect 4479 14436 4620 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 7193 14467 7251 14473
rect 7193 14433 7205 14467
rect 7239 14464 7251 14467
rect 9214 14464 9220 14476
rect 7239 14436 9220 14464
rect 7239 14433 7251 14436
rect 7193 14427 7251 14433
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9508 14464 9536 14563
rect 12710 14560 12716 14612
rect 12768 14600 12774 14612
rect 14182 14600 14188 14612
rect 12768 14572 14188 14600
rect 12768 14560 12774 14572
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 17402 14600 17408 14612
rect 16224 14572 17408 14600
rect 11606 14532 11612 14544
rect 9324 14436 9536 14464
rect 9600 14504 11612 14532
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 2498 14396 2504 14408
rect 1627 14368 2504 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6328 14368 6469 14396
rect 6328 14356 6334 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14396 7159 14399
rect 7282 14396 7288 14408
rect 7147 14368 7288 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14398 7803 14399
rect 7791 14370 7880 14398
rect 8386 14396 8392 14408
rect 7791 14365 7803 14370
rect 7745 14359 7803 14365
rect 2866 14288 2872 14340
rect 2924 14328 2930 14340
rect 3421 14331 3479 14337
rect 2924 14300 2969 14328
rect 2924 14288 2930 14300
rect 3421 14297 3433 14331
rect 3467 14328 3479 14331
rect 3510 14328 3516 14340
rect 3467 14300 3516 14328
rect 3467 14297 3479 14300
rect 3421 14291 3479 14297
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 4525 14331 4583 14337
rect 4525 14297 4537 14331
rect 4571 14328 4583 14331
rect 4706 14328 4712 14340
rect 4571 14300 4712 14328
rect 4571 14297 4583 14300
rect 4525 14291 4583 14297
rect 4706 14288 4712 14300
rect 4764 14288 4770 14340
rect 5442 14328 5448 14340
rect 5403 14300 5448 14328
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 6549 14331 6607 14337
rect 6549 14297 6561 14331
rect 6595 14328 6607 14331
rect 7650 14328 7656 14340
rect 6595 14300 7656 14328
rect 6595 14297 6607 14300
rect 6549 14291 6607 14297
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 7852 14328 7880 14370
rect 8347 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9324 14396 9352 14436
rect 8904 14368 9352 14396
rect 9401 14399 9459 14405
rect 8904 14356 8910 14368
rect 9401 14365 9413 14399
rect 9447 14390 9459 14399
rect 9600 14390 9628 14504
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 13722 14492 13728 14544
rect 13780 14532 13786 14544
rect 16224 14532 16252 14572
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 20714 14600 20720 14612
rect 17828 14572 20720 14600
rect 17828 14560 17834 14572
rect 20714 14560 20720 14572
rect 20772 14560 20778 14612
rect 21637 14603 21695 14609
rect 21637 14569 21649 14603
rect 21683 14600 21695 14603
rect 26050 14600 26056 14612
rect 21683 14572 26056 14600
rect 21683 14569 21695 14572
rect 21637 14563 21695 14569
rect 26050 14560 26056 14572
rect 26108 14560 26114 14612
rect 26234 14600 26240 14612
rect 26195 14572 26240 14600
rect 26234 14560 26240 14572
rect 26292 14600 26298 14612
rect 26602 14600 26608 14612
rect 26292 14572 26608 14600
rect 26292 14560 26298 14572
rect 26602 14560 26608 14572
rect 26660 14560 26666 14612
rect 27706 14560 27712 14612
rect 27764 14600 27770 14612
rect 38010 14600 38016 14612
rect 27764 14572 38016 14600
rect 27764 14560 27770 14572
rect 38010 14560 38016 14572
rect 38068 14560 38074 14612
rect 13780 14504 16252 14532
rect 13780 14492 13786 14504
rect 16298 14492 16304 14544
rect 16356 14532 16362 14544
rect 22094 14532 22100 14544
rect 16356 14504 22100 14532
rect 16356 14492 16362 14504
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 22186 14492 22192 14544
rect 22244 14532 22250 14544
rect 22244 14504 24624 14532
rect 22244 14492 22250 14504
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10781 14467 10839 14473
rect 10781 14464 10793 14467
rect 10284 14436 10793 14464
rect 10284 14424 10290 14436
rect 10781 14433 10793 14436
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12124 14436 12725 14464
rect 12124 14424 12130 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 12713 14427 12771 14433
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 14550 14464 14556 14476
rect 13228 14436 14556 14464
rect 13228 14424 13234 14436
rect 14292 14405 14320 14436
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 16758 14464 16764 14476
rect 16540 14436 16764 14464
rect 16540 14424 16546 14436
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 17770 14464 17776 14476
rect 17731 14436 17776 14464
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 18693 14467 18751 14473
rect 18693 14433 18705 14467
rect 18739 14464 18751 14467
rect 20346 14464 20352 14476
rect 18739 14436 20352 14464
rect 18739 14433 18751 14436
rect 18693 14427 18751 14433
rect 20346 14424 20352 14436
rect 20404 14424 20410 14476
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14464 20591 14467
rect 21910 14464 21916 14476
rect 20579 14436 21916 14464
rect 20579 14433 20591 14436
rect 20533 14427 20591 14433
rect 21910 14424 21916 14436
rect 21968 14424 21974 14476
rect 23474 14464 23480 14476
rect 23435 14436 23480 14464
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 9447 14365 9628 14390
rect 9401 14362 9628 14365
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14365 10103 14399
rect 9401 14359 9459 14362
rect 10045 14359 10103 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 8570 14328 8576 14340
rect 7852 14300 8576 14328
rect 8570 14288 8576 14300
rect 8628 14328 8634 14340
rect 10060 14328 10088 14359
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17368 14368 17509 14396
rect 17368 14356 17374 14368
rect 17497 14365 17509 14368
rect 17543 14396 17555 14399
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 17543 14368 18429 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 18417 14365 18429 14368
rect 18463 14365 18475 14399
rect 21542 14396 21548 14408
rect 21503 14368 21548 14396
rect 18417 14359 18475 14365
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 24596 14405 24624 14504
rect 29362 14492 29368 14544
rect 29420 14532 29426 14544
rect 30377 14535 30435 14541
rect 30377 14532 30389 14535
rect 29420 14504 30389 14532
rect 29420 14492 29426 14504
rect 30377 14501 30389 14504
rect 30423 14501 30435 14535
rect 30377 14495 30435 14501
rect 30006 14464 30012 14476
rect 26160 14436 28994 14464
rect 29967 14436 30012 14464
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 25222 14396 25228 14408
rect 25183 14368 25228 14396
rect 24581 14359 24639 14365
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 25590 14356 25596 14408
rect 25648 14396 25654 14408
rect 26160 14405 26188 14436
rect 26145 14399 26203 14405
rect 26145 14396 26157 14399
rect 25648 14368 26157 14396
rect 25648 14356 25654 14368
rect 26145 14365 26157 14368
rect 26191 14365 26203 14399
rect 27246 14396 27252 14408
rect 27207 14368 27252 14396
rect 26145 14359 26203 14365
rect 27246 14356 27252 14368
rect 27304 14356 27310 14408
rect 27706 14396 27712 14408
rect 27667 14368 27712 14396
rect 27706 14356 27712 14368
rect 27764 14356 27770 14408
rect 28350 14396 28356 14408
rect 28311 14368 28356 14396
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 8628 14300 9260 14328
rect 8628 14288 8634 14300
rect 1762 14260 1768 14272
rect 1723 14232 1768 14260
rect 1762 14220 1768 14232
rect 1820 14220 1826 14272
rect 7837 14263 7895 14269
rect 7837 14229 7849 14263
rect 7883 14260 7895 14263
rect 8018 14260 8024 14272
rect 7883 14232 8024 14260
rect 7883 14229 7895 14232
rect 7837 14223 7895 14229
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8478 14260 8484 14272
rect 8439 14232 8484 14260
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 9232 14260 9260 14300
rect 9416 14300 10824 14328
rect 9416 14260 9444 14300
rect 9232 14232 9444 14260
rect 10137 14263 10195 14269
rect 10137 14229 10149 14263
rect 10183 14260 10195 14263
rect 10686 14260 10692 14272
rect 10183 14232 10692 14260
rect 10183 14229 10195 14232
rect 10137 14223 10195 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 10796 14260 10824 14300
rect 10870 14288 10876 14340
rect 10928 14328 10934 14340
rect 11238 14328 11244 14340
rect 10928 14300 10973 14328
rect 11072 14300 11244 14328
rect 10928 14288 10934 14300
rect 11072 14260 11100 14300
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 11793 14331 11851 14337
rect 11793 14297 11805 14331
rect 11839 14328 11851 14331
rect 12342 14328 12348 14340
rect 11839 14300 12348 14328
rect 11839 14297 11851 14300
rect 11793 14291 11851 14297
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 12805 14331 12863 14337
rect 12805 14297 12817 14331
rect 12851 14297 12863 14331
rect 13722 14328 13728 14340
rect 13683 14300 13728 14328
rect 12805 14291 12863 14297
rect 10796 14232 11100 14260
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 12820 14260 12848 14291
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 14826 14288 14832 14340
rect 14884 14328 14890 14340
rect 15013 14331 15071 14337
rect 15013 14328 15025 14331
rect 14884 14300 15025 14328
rect 14884 14288 14890 14300
rect 15013 14297 15025 14300
rect 15059 14297 15071 14331
rect 15654 14328 15660 14340
rect 15615 14300 15660 14328
rect 15013 14291 15071 14297
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 16390 14328 16396 14340
rect 16351 14300 16396 14328
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 16482 14288 16488 14340
rect 16540 14328 16546 14340
rect 19242 14328 19248 14340
rect 16540 14300 19248 14328
rect 16540 14288 16546 14300
rect 19242 14288 19248 14300
rect 19300 14288 19306 14340
rect 19518 14328 19524 14340
rect 19479 14300 19524 14328
rect 19518 14288 19524 14300
rect 19576 14288 19582 14340
rect 19613 14331 19671 14337
rect 19613 14297 19625 14331
rect 19659 14297 19671 14331
rect 22830 14328 22836 14340
rect 22791 14300 22836 14328
rect 19613 14291 19671 14297
rect 11204 14232 12848 14260
rect 11204 14220 11210 14232
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 13446 14260 13452 14272
rect 13136 14232 13452 14260
rect 13136 14220 13142 14232
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 18966 14260 18972 14272
rect 15804 14232 18972 14260
rect 15804 14220 15810 14232
rect 18966 14220 18972 14232
rect 19024 14220 19030 14272
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 19628 14260 19656 14291
rect 22830 14288 22836 14300
rect 22888 14288 22894 14340
rect 22925 14331 22983 14337
rect 22925 14297 22937 14331
rect 22971 14297 22983 14331
rect 22925 14291 22983 14297
rect 19484 14232 19656 14260
rect 19484 14220 19490 14232
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 22002 14260 22008 14272
rect 20036 14232 22008 14260
rect 20036 14220 20042 14232
rect 22002 14220 22008 14232
rect 22060 14220 22066 14272
rect 22940 14260 22968 14291
rect 27338 14288 27344 14340
rect 27396 14328 27402 14340
rect 27801 14331 27859 14337
rect 27801 14328 27813 14331
rect 27396 14300 27813 14328
rect 27396 14288 27402 14300
rect 27801 14297 27813 14300
rect 27847 14297 27859 14331
rect 28966 14328 28994 14436
rect 30006 14424 30012 14436
rect 30064 14424 30070 14476
rect 30190 14464 30196 14476
rect 30151 14436 30196 14464
rect 30190 14424 30196 14436
rect 30248 14424 30254 14476
rect 38194 14328 38200 14340
rect 28966 14300 38200 14328
rect 27801 14291 27859 14297
rect 38194 14288 38200 14300
rect 38252 14288 38258 14340
rect 24673 14263 24731 14269
rect 24673 14260 24685 14263
rect 22940 14232 24685 14260
rect 24673 14229 24685 14232
rect 24719 14229 24731 14263
rect 25314 14260 25320 14272
rect 25275 14232 25320 14260
rect 24673 14223 24731 14229
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 27065 14263 27123 14269
rect 27065 14229 27077 14263
rect 27111 14260 27123 14263
rect 27706 14260 27712 14272
rect 27111 14232 27712 14260
rect 27111 14229 27123 14232
rect 27065 14223 27123 14229
rect 27706 14220 27712 14232
rect 27764 14220 27770 14272
rect 28166 14220 28172 14272
rect 28224 14260 28230 14272
rect 28445 14263 28503 14269
rect 28445 14260 28457 14263
rect 28224 14232 28457 14260
rect 28224 14220 28230 14232
rect 28445 14229 28457 14232
rect 28491 14229 28503 14263
rect 28445 14223 28503 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 4856 14028 5917 14056
rect 4856 14016 4862 14028
rect 5905 14025 5917 14028
rect 5951 14025 5963 14059
rect 5905 14019 5963 14025
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 8294 14056 8300 14068
rect 6687 14028 8300 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 12066 14056 12072 14068
rect 9048 14028 12072 14056
rect 3050 13988 3056 14000
rect 1596 13960 3056 13988
rect 1596 13929 1624 13960
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 3326 13988 3332 14000
rect 3287 13960 3332 13988
rect 3326 13948 3332 13960
rect 3384 13948 3390 14000
rect 4617 13991 4675 13997
rect 4617 13957 4629 13991
rect 4663 13988 4675 13991
rect 5258 13988 5264 14000
rect 4663 13960 5264 13988
rect 4663 13957 4675 13960
rect 4617 13951 4675 13957
rect 5258 13948 5264 13960
rect 5316 13948 5322 14000
rect 7282 13988 7288 14000
rect 7243 13960 7288 13988
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 7650 13948 7656 14000
rect 7708 13988 7714 14000
rect 9048 13988 9076 14028
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 15102 14056 15108 14068
rect 12406 14028 15108 14056
rect 10134 13988 10140 14000
rect 7708 13960 9076 13988
rect 9324 13960 10140 13988
rect 7708 13948 7714 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2682 13920 2688 13932
rect 2547 13892 2688 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 4522 13920 4528 13932
rect 4483 13892 4528 13920
rect 4522 13880 4528 13892
rect 4580 13920 4586 13932
rect 4706 13920 4712 13932
rect 4580 13892 4712 13920
rect 4580 13880 4586 13892
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 4890 13880 4896 13932
rect 4948 13920 4954 13932
rect 5169 13923 5227 13929
rect 5169 13920 5181 13923
rect 4948 13892 5181 13920
rect 4948 13880 4954 13892
rect 5169 13889 5181 13892
rect 5215 13920 5227 13923
rect 5442 13920 5448 13932
rect 5215 13892 5448 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5592 13892 5825 13920
rect 5592 13880 5598 13892
rect 5813 13889 5825 13892
rect 5859 13920 5871 13923
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 5859 13892 6561 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6549 13889 6561 13892
rect 6595 13920 6607 13923
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6595 13892 7205 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 7193 13889 7205 13892
rect 7239 13920 7251 13923
rect 7834 13920 7840 13932
rect 7239 13892 7840 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8352 13892 8493 13920
rect 8352 13880 8358 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 9324 13918 9352 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 10229 13991 10287 13997
rect 10229 13957 10241 13991
rect 10275 13988 10287 13991
rect 12406 13988 12434 14028
rect 15102 14016 15108 14028
rect 15160 14056 15166 14068
rect 15654 14056 15660 14068
rect 15160 14028 15660 14056
rect 15160 14016 15166 14028
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 19150 14056 19156 14068
rect 17604 14028 19156 14056
rect 12526 13988 12532 14000
rect 10275 13960 12434 13988
rect 12487 13960 12532 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 12621 13991 12679 13997
rect 12621 13957 12633 13991
rect 12667 13988 12679 13991
rect 13446 13988 13452 14000
rect 12667 13960 13452 13988
rect 12667 13957 12679 13960
rect 12621 13951 12679 13957
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 14182 13988 14188 14000
rect 14143 13960 14188 13988
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 15746 13988 15752 14000
rect 14700 13960 15332 13988
rect 15707 13960 15752 13988
rect 14700 13948 14706 13960
rect 8481 13883 8539 13889
rect 9140 13890 9352 13918
rect 9769 13923 9827 13929
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3510 13852 3516 13864
rect 3283 13824 3372 13852
rect 3471 13824 3516 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3344 13784 3372 13824
rect 3510 13812 3516 13824
rect 3568 13852 3574 13864
rect 3878 13852 3884 13864
rect 3568 13824 3884 13852
rect 3568 13812 3574 13824
rect 3878 13812 3884 13824
rect 3936 13812 3942 13864
rect 3988 13824 5028 13852
rect 3988 13784 4016 13824
rect 3344 13756 4016 13784
rect 5000 13784 5028 13824
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5132 13824 5273 13852
rect 5132 13812 5138 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 7006 13852 7012 13864
rect 5261 13815 5319 13821
rect 5368 13824 7012 13852
rect 5368 13784 5396 13824
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13852 8631 13855
rect 8846 13852 8852 13864
rect 8619 13824 8852 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9140 13861 9168 13890
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 9950 13920 9956 13932
rect 9815 13892 9956 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12158 13920 12164 13932
rect 11931 13892 12164 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 9309 13855 9367 13861
rect 9309 13821 9321 13855
rect 9355 13821 9367 13855
rect 11054 13852 11060 13864
rect 11015 13824 11060 13852
rect 9309 13815 9367 13821
rect 6454 13784 6460 13796
rect 5000 13756 5396 13784
rect 5920 13756 6460 13784
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 3970 13716 3976 13728
rect 2639 13688 3976 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 5166 13716 5172 13728
rect 4948 13688 5172 13716
rect 4948 13676 4954 13688
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5920 13716 5948 13756
rect 6454 13744 6460 13756
rect 6512 13744 6518 13796
rect 5408 13688 5948 13716
rect 5408 13676 5414 13688
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 7006 13716 7012 13728
rect 6052 13688 7012 13716
rect 6052 13676 6058 13688
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 7929 13719 7987 13725
rect 7929 13685 7941 13719
rect 7975 13716 7987 13719
rect 8570 13716 8576 13728
rect 7975 13688 8576 13716
rect 7975 13685 7987 13688
rect 7929 13679 7987 13685
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 9030 13676 9036 13728
rect 9088 13716 9094 13728
rect 9324 13716 9352 13815
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11808 13852 11836 13883
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13906 13920 13912 13932
rect 13372 13892 13912 13920
rect 13372 13852 13400 13892
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 15194 13920 15200 13932
rect 15028 13892 15200 13920
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 11808 13824 13400 13852
rect 13464 13824 13553 13852
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 13464 13784 13492 13824
rect 13541 13821 13553 13824
rect 13587 13852 13599 13855
rect 14090 13852 14096 13864
rect 13587 13824 13952 13852
rect 14051 13824 14096 13852
rect 13587 13821 13599 13824
rect 13541 13815 13599 13821
rect 13044 13756 13492 13784
rect 13924 13784 13952 13824
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 15028 13852 15056 13892
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15304 13920 15332 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 16298 13988 16304 14000
rect 16259 13960 16304 13988
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 17034 13988 17040 14000
rect 16995 13960 17040 13988
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 17604 13997 17632 14028
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 20254 14016 20260 14068
rect 20312 14056 20318 14068
rect 24857 14059 24915 14065
rect 24857 14056 24869 14059
rect 20312 14028 24869 14056
rect 20312 14016 20318 14028
rect 24857 14025 24869 14028
rect 24903 14025 24915 14059
rect 24857 14019 24915 14025
rect 25501 14059 25559 14065
rect 25501 14025 25513 14059
rect 25547 14056 25559 14059
rect 29914 14056 29920 14068
rect 25547 14028 29920 14056
rect 25547 14025 25559 14028
rect 25501 14019 25559 14025
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 17589 13991 17647 13997
rect 17589 13957 17601 13991
rect 17635 13957 17647 13991
rect 17589 13951 17647 13957
rect 17770 13948 17776 14000
rect 17828 13988 17834 14000
rect 18969 13991 19027 13997
rect 18969 13988 18981 13991
rect 17828 13960 18981 13988
rect 17828 13948 17834 13960
rect 18969 13957 18981 13960
rect 19015 13957 19027 13991
rect 18969 13951 19027 13957
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19889 13991 19947 13997
rect 19889 13988 19901 13991
rect 19300 13960 19901 13988
rect 19300 13948 19306 13960
rect 19889 13957 19901 13960
rect 19935 13957 19947 13991
rect 19889 13951 19947 13957
rect 20533 13991 20591 13997
rect 20533 13957 20545 13991
rect 20579 13988 20591 13991
rect 21082 13988 21088 14000
rect 20579 13960 21088 13988
rect 20579 13957 20591 13960
rect 20533 13951 20591 13957
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 23106 13988 23112 14000
rect 22152 13960 23112 13988
rect 22152 13948 22158 13960
rect 23106 13948 23112 13960
rect 23164 13948 23170 14000
rect 23385 13991 23443 13997
rect 23385 13957 23397 13991
rect 23431 13988 23443 13991
rect 25314 13988 25320 14000
rect 23431 13960 25320 13988
rect 23431 13957 23443 13960
rect 23385 13951 23443 13957
rect 25314 13948 25320 13960
rect 25372 13948 25378 14000
rect 27338 13988 27344 14000
rect 27299 13960 27344 13988
rect 27338 13948 27344 13960
rect 27396 13948 27402 14000
rect 27706 13948 27712 14000
rect 27764 13988 27770 14000
rect 29457 13991 29515 13997
rect 29457 13988 29469 13991
rect 27764 13960 29469 13988
rect 27764 13948 27770 13960
rect 29457 13957 29469 13960
rect 29503 13957 29515 13991
rect 29457 13951 29515 13957
rect 18138 13920 18144 13932
rect 15304 13892 15516 13920
rect 18099 13892 18144 13920
rect 14200 13824 15056 13852
rect 15105 13855 15163 13861
rect 14200 13784 14228 13824
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15378 13852 15384 13864
rect 15151 13824 15384 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15488 13852 15516 13892
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21284 13892 22017 13920
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 15488 13824 15669 13852
rect 15657 13821 15669 13824
rect 15703 13821 15715 13855
rect 15657 13815 15715 13821
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 15896 13824 16957 13852
rect 15896 13812 15902 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 16945 13815 17003 13821
rect 18233 13855 18291 13861
rect 18233 13821 18245 13855
rect 18279 13852 18291 13855
rect 18877 13855 18935 13861
rect 18279 13824 18828 13852
rect 18279 13821 18291 13824
rect 18233 13815 18291 13821
rect 13924 13756 14228 13784
rect 15396 13784 15424 13812
rect 16666 13784 16672 13796
rect 15396 13756 16672 13784
rect 13044 13744 13050 13756
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 18800 13784 18828 13824
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 19242 13852 19248 13864
rect 18923 13824 19248 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 19334 13812 19340 13864
rect 19392 13812 19398 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 20364 13824 20453 13852
rect 19352 13784 19380 13812
rect 20364 13796 20392 13824
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 21284 13852 21312 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 22005 13883 22063 13889
rect 24136 13892 24777 13920
rect 20680 13824 21312 13852
rect 20680 13812 20686 13824
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 21416 13824 21509 13852
rect 21416 13812 21422 13824
rect 22830 13812 22836 13864
rect 22888 13852 22894 13864
rect 23293 13855 23351 13861
rect 23293 13852 23305 13855
rect 22888 13824 23305 13852
rect 22888 13812 22894 13824
rect 23293 13821 23305 13824
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 18800 13756 19380 13784
rect 20346 13744 20352 13796
rect 20404 13744 20410 13796
rect 20714 13744 20720 13796
rect 20772 13784 20778 13796
rect 21376 13784 21404 13812
rect 20772 13756 21404 13784
rect 23308 13784 23336 13815
rect 23382 13812 23388 13864
rect 23440 13852 23446 13864
rect 24136 13852 24164 13892
rect 24765 13889 24777 13892
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 24302 13852 24308 13864
rect 23440 13824 24164 13852
rect 24263 13824 24308 13852
rect 23440 13812 23446 13824
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 24394 13812 24400 13864
rect 24452 13852 24458 13864
rect 25424 13852 25452 13883
rect 27890 13880 27896 13932
rect 27948 13920 27954 13932
rect 27948 13892 27993 13920
rect 27948 13880 27954 13892
rect 37274 13880 37280 13932
rect 37332 13920 37338 13932
rect 37737 13923 37795 13929
rect 37737 13920 37749 13923
rect 37332 13892 37749 13920
rect 37332 13880 37338 13892
rect 37737 13889 37749 13892
rect 37783 13889 37795 13923
rect 37737 13883 37795 13889
rect 27246 13852 27252 13864
rect 24452 13824 25452 13852
rect 25516 13824 27108 13852
rect 27207 13824 27252 13852
rect 24452 13812 24458 13824
rect 24578 13784 24584 13796
rect 23308 13756 24584 13784
rect 20772 13744 20778 13756
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 9088 13688 9352 13716
rect 9088 13676 9094 13688
rect 10134 13676 10140 13728
rect 10192 13716 10198 13728
rect 11330 13716 11336 13728
rect 10192 13688 11336 13716
rect 10192 13676 10198 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 18690 13716 18696 13728
rect 13780 13688 18696 13716
rect 13780 13676 13786 13688
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 21910 13716 21916 13728
rect 20220 13688 21916 13716
rect 20220 13676 20226 13688
rect 21910 13676 21916 13688
rect 21968 13676 21974 13728
rect 22094 13716 22100 13728
rect 22055 13688 22100 13716
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 23106 13676 23112 13728
rect 23164 13716 23170 13728
rect 24302 13716 24308 13728
rect 23164 13688 24308 13716
rect 23164 13676 23170 13688
rect 24302 13676 24308 13688
rect 24360 13716 24366 13728
rect 25516 13716 25544 13824
rect 27080 13784 27108 13824
rect 27246 13812 27252 13824
rect 27304 13812 27310 13864
rect 27908 13852 27936 13880
rect 29362 13852 29368 13864
rect 27356 13824 27936 13852
rect 29323 13824 29368 13852
rect 27356 13784 27384 13824
rect 29362 13812 29368 13824
rect 29420 13812 29426 13864
rect 29638 13852 29644 13864
rect 29599 13824 29644 13852
rect 29638 13812 29644 13824
rect 29696 13812 29702 13864
rect 37182 13812 37188 13864
rect 37240 13852 37246 13864
rect 37461 13855 37519 13861
rect 37461 13852 37473 13855
rect 37240 13824 37473 13852
rect 37240 13812 37246 13824
rect 37461 13821 37473 13824
rect 37507 13821 37519 13855
rect 37461 13815 37519 13821
rect 27080 13756 27384 13784
rect 24360 13688 25544 13716
rect 24360 13676 24366 13688
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 3786 13472 3792 13524
rect 3844 13512 3850 13524
rect 5994 13512 6000 13524
rect 3844 13484 6000 13512
rect 3844 13472 3850 13484
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 7282 13512 7288 13524
rect 6236 13484 7288 13512
rect 6236 13472 6242 13484
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9122 13512 9128 13524
rect 8812 13484 9128 13512
rect 8812 13472 8818 13484
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 12710 13512 12716 13524
rect 9646 13484 12716 13512
rect 9646 13444 9674 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12860 13484 13001 13512
rect 12860 13472 12866 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 15378 13512 15384 13524
rect 14424 13484 15384 13512
rect 14424 13472 14430 13484
rect 15378 13472 15384 13484
rect 15436 13472 15442 13524
rect 16114 13472 16120 13524
rect 16172 13512 16178 13524
rect 16298 13512 16304 13524
rect 16172 13484 16304 13512
rect 16172 13472 16178 13484
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 16724 13484 21404 13512
rect 16724 13472 16730 13484
rect 2884 13416 9674 13444
rect 2884 13385 2912 13416
rect 11238 13404 11244 13456
rect 11296 13444 11302 13456
rect 15930 13444 15936 13456
rect 11296 13416 11376 13444
rect 11296 13404 11302 13416
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 6914 13376 6920 13388
rect 4663 13348 6920 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7282 13376 7288 13388
rect 7243 13348 7288 13376
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 9766 13376 9772 13388
rect 9727 13348 9772 13376
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 11348 13376 11376 13416
rect 13556 13416 15936 13444
rect 13556 13376 13584 13416
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 11348 13348 13584 13376
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5534 13308 5540 13320
rect 5399 13280 5540 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 1946 13200 1952 13252
rect 2004 13240 2010 13252
rect 4540 13240 4568 13271
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5684 13280 6009 13308
rect 5684 13268 5690 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 6178 13308 6184 13320
rect 6135 13280 6184 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 2004 13212 2049 13240
rect 4540 13212 5580 13240
rect 2004 13200 2010 13212
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5445 13175 5503 13181
rect 5445 13172 5457 13175
rect 5224 13144 5457 13172
rect 5224 13132 5230 13144
rect 5445 13141 5457 13144
rect 5491 13141 5503 13175
rect 5552 13172 5580 13212
rect 5810 13200 5816 13252
rect 5868 13240 5874 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 5868 13212 6745 13240
rect 5868 13200 5874 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6733 13203 6791 13209
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 6880 13212 6925 13240
rect 6880 13200 6886 13212
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 8294 13240 8300 13252
rect 7064 13212 8300 13240
rect 7064 13200 7070 13212
rect 8294 13200 8300 13212
rect 8352 13240 8358 13252
rect 8404 13240 8432 13271
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 13556 13317 13584 13348
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 17310 13376 17316 13388
rect 13679 13348 17316 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 18800 13385 18828 13484
rect 19150 13404 19156 13456
rect 19208 13444 19214 13456
rect 21376 13444 21404 13484
rect 21450 13472 21456 13524
rect 21508 13512 21514 13524
rect 25038 13512 25044 13524
rect 21508 13484 25044 13512
rect 21508 13472 21514 13484
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 27982 13444 27988 13456
rect 19208 13416 21312 13444
rect 21376 13416 27988 13444
rect 19208 13404 19214 13416
rect 18785 13379 18843 13385
rect 17604 13348 18736 13376
rect 11241 13311 11299 13317
rect 11241 13310 11253 13311
rect 11164 13308 11253 13310
rect 11112 13282 11253 13308
rect 11112 13280 11192 13282
rect 11112 13268 11118 13280
rect 11241 13277 11253 13282
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 9582 13240 9588 13252
rect 8352 13212 9588 13240
rect 8352 13200 8358 13212
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 9861 13243 9919 13249
rect 9861 13240 9873 13243
rect 9824 13212 9873 13240
rect 9824 13200 9830 13212
rect 9861 13209 9873 13212
rect 9907 13209 9919 13243
rect 9861 13203 9919 13209
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 11514 13240 11520 13252
rect 11204 13212 11520 13240
rect 11204 13200 11210 13212
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 12526 13200 12532 13252
rect 12584 13200 12590 13252
rect 14366 13240 14372 13252
rect 14327 13212 14372 13240
rect 14366 13200 14372 13212
rect 14424 13200 14430 13252
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 14516 13212 14561 13240
rect 14516 13200 14522 13212
rect 15194 13200 15200 13252
rect 15252 13240 15258 13252
rect 15381 13243 15439 13249
rect 15381 13240 15393 13243
rect 15252 13212 15393 13240
rect 15252 13200 15258 13212
rect 15381 13209 15393 13212
rect 15427 13209 15439 13243
rect 15381 13203 15439 13209
rect 8110 13172 8116 13184
rect 5552 13144 8116 13172
rect 5445 13135 5503 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8386 13132 8392 13184
rect 8444 13172 8450 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8444 13144 8493 13172
rect 8444 13132 8450 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 12342 13172 12348 13184
rect 9272 13144 12348 13172
rect 9272 13132 9278 13144
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 12802 13132 12808 13184
rect 12860 13172 12866 13184
rect 13998 13172 14004 13184
rect 12860 13144 14004 13172
rect 12860 13132 12866 13144
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 15396 13172 15424 13203
rect 15838 13200 15844 13252
rect 15896 13240 15902 13252
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15896 13212 16221 13240
rect 15896 13200 15902 13212
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 16301 13243 16359 13249
rect 16301 13209 16313 13243
rect 16347 13240 16359 13243
rect 16574 13240 16580 13252
rect 16347 13212 16580 13240
rect 16347 13209 16359 13212
rect 16301 13203 16359 13209
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 17221 13243 17279 13249
rect 17221 13209 17233 13243
rect 17267 13240 17279 13243
rect 17402 13240 17408 13252
rect 17267 13212 17408 13240
rect 17267 13209 17279 13212
rect 17221 13203 17279 13209
rect 17402 13200 17408 13212
rect 17460 13200 17466 13252
rect 17604 13240 17632 13348
rect 18708 13308 18736 13348
rect 18785 13345 18797 13379
rect 18831 13345 18843 13379
rect 20806 13376 20812 13388
rect 18785 13339 18843 13345
rect 19306 13348 20812 13376
rect 19306 13308 19334 13348
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 21177 13311 21235 13317
rect 21177 13308 21189 13311
rect 18708 13280 19334 13308
rect 20548 13280 21189 13308
rect 17773 13243 17831 13249
rect 17773 13240 17785 13243
rect 17604 13212 17785 13240
rect 17773 13209 17785 13212
rect 17819 13209 17831 13243
rect 17773 13203 17831 13209
rect 16482 13172 16488 13184
rect 15396 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 17034 13132 17040 13184
rect 17092 13172 17098 13184
rect 17788 13172 17816 13203
rect 17862 13200 17868 13252
rect 17920 13240 17926 13252
rect 17920 13212 17965 13240
rect 17920 13200 17926 13212
rect 18322 13200 18328 13252
rect 18380 13240 18386 13252
rect 19426 13240 19432 13252
rect 18380 13212 19432 13240
rect 18380 13200 18386 13212
rect 19426 13200 19432 13212
rect 19484 13240 19490 13252
rect 19705 13243 19763 13249
rect 19705 13240 19717 13243
rect 19484 13212 19717 13240
rect 19484 13200 19490 13212
rect 19705 13209 19717 13212
rect 19751 13209 19763 13243
rect 19705 13203 19763 13209
rect 19794 13200 19800 13252
rect 19852 13240 19858 13252
rect 19852 13212 19897 13240
rect 19852 13200 19858 13212
rect 20162 13200 20168 13252
rect 20220 13240 20226 13252
rect 20548 13240 20576 13280
rect 21177 13277 21189 13280
rect 21223 13277 21235 13311
rect 21177 13271 21235 13277
rect 20220 13212 20576 13240
rect 20220 13200 20226 13212
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 21284 13240 21312 13416
rect 27982 13404 27988 13416
rect 28040 13404 28046 13456
rect 25866 13376 25872 13388
rect 22480 13348 25872 13376
rect 21358 13268 21364 13320
rect 21416 13308 21422 13320
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 21416 13280 21833 13308
rect 21416 13268 21422 13280
rect 21821 13277 21833 13280
rect 21867 13277 21879 13311
rect 21821 13271 21879 13277
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22480 13317 22508 13348
rect 25866 13336 25872 13348
rect 25924 13336 25930 13388
rect 25958 13336 25964 13388
rect 26016 13376 26022 13388
rect 28353 13379 28411 13385
rect 28353 13376 28365 13379
rect 26016 13348 28365 13376
rect 26016 13336 26022 13348
rect 28353 13345 28365 13348
rect 28399 13345 28411 13379
rect 28353 13339 28411 13345
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 21968 13280 22477 13308
rect 21968 13268 21974 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 22646 13268 22652 13320
rect 22704 13308 22710 13320
rect 22830 13308 22836 13320
rect 22704 13280 22836 13308
rect 22704 13268 22710 13280
rect 22830 13268 22836 13280
rect 22888 13308 22894 13320
rect 23109 13311 23167 13317
rect 23109 13308 23121 13311
rect 22888 13280 23121 13308
rect 22888 13268 22894 13280
rect 23109 13277 23121 13280
rect 23155 13308 23167 13311
rect 23382 13308 23388 13320
rect 23155 13280 23388 13308
rect 23155 13277 23167 13280
rect 23109 13271 23167 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23750 13308 23756 13320
rect 23711 13280 23756 13308
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 23201 13243 23259 13249
rect 23201 13240 23213 13243
rect 20772 13212 20817 13240
rect 21284 13212 23213 13240
rect 20772 13200 20778 13212
rect 23201 13209 23213 13212
rect 23247 13209 23259 13243
rect 23201 13203 23259 13209
rect 24302 13200 24308 13252
rect 24360 13240 24366 13252
rect 24673 13243 24731 13249
rect 24673 13240 24685 13243
rect 24360 13212 24685 13240
rect 24360 13200 24366 13212
rect 24673 13209 24685 13212
rect 24719 13209 24731 13243
rect 24673 13203 24731 13209
rect 24765 13243 24823 13249
rect 24765 13209 24777 13243
rect 24811 13209 24823 13243
rect 25682 13240 25688 13252
rect 25643 13212 25688 13240
rect 24765 13203 24823 13209
rect 17092 13144 17816 13172
rect 17092 13132 17098 13144
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 18966 13172 18972 13184
rect 18564 13144 18972 13172
rect 18564 13132 18570 13144
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 21266 13132 21272 13184
rect 21324 13172 21330 13184
rect 21913 13175 21971 13181
rect 21324 13144 21369 13172
rect 21324 13132 21330 13144
rect 21913 13141 21925 13175
rect 21959 13172 21971 13175
rect 22002 13172 22008 13184
rect 21959 13144 22008 13172
rect 21959 13141 21971 13144
rect 21913 13135 21971 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22557 13175 22615 13181
rect 22557 13172 22569 13175
rect 22152 13144 22569 13172
rect 22152 13132 22158 13144
rect 22557 13141 22569 13144
rect 22603 13141 22615 13175
rect 22557 13135 22615 13141
rect 23845 13175 23903 13181
rect 23845 13141 23857 13175
rect 23891 13172 23903 13175
rect 24780 13172 24808 13203
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 26237 13243 26295 13249
rect 26237 13209 26249 13243
rect 26283 13209 26295 13243
rect 26237 13203 26295 13209
rect 23891 13144 24808 13172
rect 26252 13172 26280 13203
rect 26326 13200 26332 13252
rect 26384 13240 26390 13252
rect 26384 13212 26429 13240
rect 26384 13200 26390 13212
rect 27154 13200 27160 13252
rect 27212 13240 27218 13252
rect 27249 13243 27307 13249
rect 27249 13240 27261 13243
rect 27212 13212 27261 13240
rect 27212 13200 27218 13212
rect 27249 13209 27261 13212
rect 27295 13209 27307 13243
rect 28074 13240 28080 13252
rect 28035 13212 28080 13240
rect 27249 13203 27307 13209
rect 28074 13200 28080 13212
rect 28132 13200 28138 13252
rect 28166 13200 28172 13252
rect 28224 13240 28230 13252
rect 28224 13212 28269 13240
rect 28224 13200 28230 13212
rect 29454 13172 29460 13184
rect 26252 13144 29460 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 29454 13132 29460 13144
rect 29512 13132 29518 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 3970 12928 3976 12980
rect 4028 12968 4034 12980
rect 4028 12940 8156 12968
rect 4028 12928 4034 12940
rect 5626 12900 5632 12912
rect 3436 12872 5632 12900
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 2774 12792 2780 12844
rect 2832 12832 2838 12844
rect 3436 12841 3464 12872
rect 5626 12860 5632 12872
rect 5684 12900 5690 12912
rect 6270 12900 6276 12912
rect 5684 12872 6276 12900
rect 5684 12860 5690 12872
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 6822 12900 6828 12912
rect 6783 12872 6828 12900
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 7374 12900 7380 12912
rect 7335 12872 7380 12900
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 7466 12860 7472 12912
rect 7524 12900 7530 12912
rect 8021 12903 8079 12909
rect 8021 12900 8033 12903
rect 7524 12872 8033 12900
rect 7524 12860 7530 12872
rect 8021 12869 8033 12872
rect 8067 12869 8079 12903
rect 8128 12900 8156 12940
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9398 12968 9404 12980
rect 9272 12940 9404 12968
rect 9272 12928 9278 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9640 12940 11008 12968
rect 9640 12928 9646 12940
rect 8128 12872 10166 12900
rect 8021 12863 8079 12869
rect 3421 12835 3479 12841
rect 2832 12804 2877 12832
rect 2832 12792 2838 12804
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3786 12792 3792 12844
rect 3844 12832 3850 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3844 12804 4077 12832
rect 3844 12792 3850 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4706 12832 4712 12844
rect 4667 12804 4712 12832
rect 4065 12795 4123 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5534 12832 5540 12844
rect 5399 12804 5540 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 10980 12832 11008 12940
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11882 12968 11888 12980
rect 11756 12940 11888 12968
rect 11756 12928 11762 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 15654 12968 15660 12980
rect 12492 12940 14044 12968
rect 12492 12928 12498 12940
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 11112 12872 11836 12900
rect 11112 12860 11118 12872
rect 11238 12832 11244 12844
rect 10980 12804 11244 12832
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11572 12804 11713 12832
rect 11572 12792 11578 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11808 12832 11836 12872
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12124 12872 13110 12900
rect 12124 12860 12130 12872
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 11808 12804 12357 12832
rect 11701 12795 11759 12801
rect 12345 12801 12357 12804
rect 12391 12801 12403 12835
rect 12345 12795 12403 12801
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4203 12668 4936 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 4908 12640 4936 12668
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 2866 12628 2872 12640
rect 2827 12600 2872 12628
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3510 12628 3516 12640
rect 3471 12600 3516 12628
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 4706 12588 4712 12640
rect 4764 12628 4770 12640
rect 4801 12631 4859 12637
rect 4801 12628 4813 12631
rect 4764 12600 4813 12628
rect 4764 12588 4770 12600
rect 4801 12597 4813 12600
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 4890 12588 4896 12640
rect 4948 12588 4954 12640
rect 5000 12628 5028 12792
rect 6564 12764 6592 12792
rect 6733 12767 6791 12773
rect 6733 12764 6745 12767
rect 6564 12736 6745 12764
rect 6733 12733 6745 12736
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12764 8999 12767
rect 9214 12764 9220 12776
rect 8987 12736 9220 12764
rect 8987 12733 8999 12736
rect 8941 12727 8999 12733
rect 5445 12699 5503 12705
rect 5445 12665 5457 12699
rect 5491 12696 5503 12699
rect 6086 12696 6092 12708
rect 5491 12668 6092 12696
rect 5491 12665 5503 12668
rect 5445 12659 5503 12665
rect 6086 12656 6092 12668
rect 6144 12656 6150 12708
rect 6454 12656 6460 12708
rect 6512 12696 6518 12708
rect 7944 12696 7972 12727
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9398 12764 9404 12776
rect 9359 12736 9404 12764
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 10042 12764 10048 12776
rect 9723 12736 10048 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 10042 12724 10048 12736
rect 10100 12764 10106 12776
rect 10410 12764 10416 12776
rect 10100 12736 10416 12764
rect 10100 12724 10106 12736
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 12618 12764 12624 12776
rect 12579 12736 12624 12764
rect 12618 12724 12624 12736
rect 12676 12724 12682 12776
rect 14016 12764 14044 12940
rect 14568 12940 15660 12968
rect 14568 12844 14596 12940
rect 15654 12928 15660 12940
rect 15712 12968 15718 12980
rect 16390 12968 16396 12980
rect 15712 12940 16396 12968
rect 15712 12928 15718 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 23569 12971 23627 12977
rect 23569 12968 23581 12971
rect 18616 12940 23581 12968
rect 14734 12860 14740 12912
rect 14792 12900 14798 12912
rect 14829 12903 14887 12909
rect 14829 12900 14841 12903
rect 14792 12872 14841 12900
rect 14792 12860 14798 12872
rect 14829 12869 14841 12872
rect 14875 12869 14887 12903
rect 18616 12900 18644 12940
rect 23569 12937 23581 12940
rect 23615 12937 23627 12971
rect 23569 12931 23627 12937
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 24762 12968 24768 12980
rect 24268 12940 24768 12968
rect 24268 12928 24274 12940
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25314 12928 25320 12980
rect 25372 12968 25378 12980
rect 25682 12968 25688 12980
rect 25372 12940 25688 12968
rect 25372 12928 25378 12940
rect 25682 12928 25688 12940
rect 25740 12968 25746 12980
rect 25740 12940 28396 12968
rect 25740 12928 25746 12940
rect 21177 12903 21235 12909
rect 21177 12900 21189 12903
rect 16054 12872 18644 12900
rect 19458 12872 21189 12900
rect 14829 12863 14887 12869
rect 21177 12869 21189 12872
rect 21223 12869 21235 12903
rect 22370 12900 22376 12912
rect 22331 12872 22376 12900
rect 21177 12863 21235 12869
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 22465 12903 22523 12909
rect 22465 12869 22477 12903
rect 22511 12900 22523 12903
rect 24857 12903 24915 12909
rect 24857 12900 24869 12903
rect 22511 12872 24869 12900
rect 22511 12869 22523 12872
rect 22465 12863 22523 12869
rect 24857 12869 24869 12872
rect 24903 12869 24915 12903
rect 24857 12863 24915 12869
rect 26786 12860 26792 12912
rect 26844 12900 26850 12912
rect 28368 12909 28396 12940
rect 29362 12928 29368 12980
rect 29420 12968 29426 12980
rect 29457 12971 29515 12977
rect 29457 12968 29469 12971
rect 29420 12940 29469 12968
rect 29420 12928 29426 12940
rect 29457 12937 29469 12940
rect 29503 12937 29515 12971
rect 29457 12931 29515 12937
rect 27433 12903 27491 12909
rect 27433 12900 27445 12903
rect 26844 12872 27445 12900
rect 26844 12860 26850 12872
rect 27433 12869 27445 12872
rect 27479 12869 27491 12903
rect 27433 12863 27491 12869
rect 28353 12903 28411 12909
rect 28353 12869 28365 12903
rect 28399 12900 28411 12903
rect 36722 12900 36728 12912
rect 28399 12872 36728 12900
rect 28399 12869 28411 12872
rect 28353 12863 28411 12869
rect 36722 12860 36728 12872
rect 36780 12860 36786 12912
rect 14550 12832 14556 12844
rect 14463 12804 14556 12832
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 16850 12832 16856 12844
rect 16811 12804 16856 12832
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 20438 12832 20444 12844
rect 19628 12804 20444 12832
rect 16114 12764 16120 12776
rect 14016 12736 16120 12764
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16298 12764 16304 12776
rect 16259 12736 16304 12764
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 17034 12764 17040 12776
rect 16995 12736 17040 12764
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17954 12764 17960 12776
rect 17915 12736 17960 12764
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18230 12764 18236 12776
rect 18191 12736 18236 12764
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 18690 12724 18696 12776
rect 18748 12764 18754 12776
rect 19628 12764 19656 12804
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21085 12835 21143 12841
rect 21085 12832 21097 12835
rect 20772 12804 21097 12832
rect 20772 12792 20778 12804
rect 21085 12801 21097 12804
rect 21131 12832 21143 12835
rect 21450 12832 21456 12844
rect 21131 12804 21456 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 23477 12835 23535 12841
rect 23477 12832 23489 12835
rect 23440 12804 23489 12832
rect 23440 12792 23446 12804
rect 23477 12801 23489 12804
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12832 24179 12835
rect 24302 12832 24308 12844
rect 24167 12804 24308 12832
rect 24167 12801 24179 12804
rect 24121 12795 24179 12801
rect 18748 12736 19656 12764
rect 19705 12767 19763 12773
rect 18748 12724 18754 12736
rect 19705 12733 19717 12767
rect 19751 12764 19763 12767
rect 20346 12764 20352 12776
rect 19751 12736 20352 12764
rect 19751 12733 19763 12736
rect 19705 12727 19763 12733
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 20456 12764 20484 12792
rect 22646 12764 22652 12776
rect 20456 12736 22652 12764
rect 22646 12724 22652 12736
rect 22704 12724 22710 12776
rect 24136 12764 24164 12795
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 24765 12835 24823 12841
rect 24765 12801 24777 12835
rect 24811 12801 24823 12835
rect 24765 12795 24823 12801
rect 22756 12736 24164 12764
rect 6512 12668 7972 12696
rect 11149 12699 11207 12705
rect 6512 12656 6518 12668
rect 11149 12665 11161 12699
rect 11195 12696 11207 12699
rect 11698 12696 11704 12708
rect 11195 12668 11704 12696
rect 11195 12665 11207 12668
rect 11149 12659 11207 12665
rect 11698 12656 11704 12668
rect 11756 12656 11762 12708
rect 10226 12628 10232 12640
rect 5000 12600 10232 12628
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11238 12628 11244 12640
rect 11112 12600 11244 12628
rect 11112 12588 11118 12600
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 12066 12628 12072 12640
rect 11839 12600 12072 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 14093 12631 14151 12637
rect 14093 12628 14105 12631
rect 13780 12600 14105 12628
rect 13780 12588 13786 12600
rect 14093 12597 14105 12600
rect 14139 12597 14151 12631
rect 17052 12628 17080 12724
rect 22756 12696 22784 12736
rect 22922 12696 22928 12708
rect 19306 12668 22784 12696
rect 22883 12668 22928 12696
rect 19306 12628 19334 12668
rect 22922 12656 22928 12668
rect 22980 12656 22986 12708
rect 24780 12696 24808 12795
rect 36906 12792 36912 12844
rect 36964 12832 36970 12844
rect 38013 12835 38071 12841
rect 38013 12832 38025 12835
rect 36964 12804 38025 12832
rect 36964 12792 36970 12804
rect 38013 12801 38025 12804
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 27341 12767 27399 12773
rect 27341 12733 27353 12767
rect 27387 12764 27399 12767
rect 27614 12764 27620 12776
rect 27387 12736 27620 12764
rect 27387 12733 27399 12736
rect 27341 12727 27399 12733
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 28810 12764 28816 12776
rect 28771 12736 28816 12764
rect 28810 12724 28816 12736
rect 28868 12724 28874 12776
rect 28994 12764 29000 12776
rect 28955 12736 29000 12764
rect 28994 12724 29000 12736
rect 29052 12724 29058 12776
rect 23032 12668 24808 12696
rect 17052 12600 19334 12628
rect 14093 12591 14151 12597
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 20438 12628 20444 12640
rect 19484 12600 20444 12628
rect 19484 12588 19490 12600
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 20533 12631 20591 12637
rect 20533 12597 20545 12631
rect 20579 12628 20591 12631
rect 20806 12628 20812 12640
rect 20579 12600 20812 12628
rect 20579 12597 20591 12600
rect 20533 12591 20591 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 21726 12588 21732 12640
rect 21784 12628 21790 12640
rect 23032 12628 23060 12668
rect 24210 12628 24216 12640
rect 21784 12600 23060 12628
rect 24171 12600 24216 12628
rect 21784 12588 21790 12600
rect 24210 12588 24216 12600
rect 24268 12588 24274 12640
rect 24302 12588 24308 12640
rect 24360 12628 24366 12640
rect 27522 12628 27528 12640
rect 24360 12600 27528 12628
rect 24360 12588 24366 12600
rect 27522 12588 27528 12600
rect 27580 12588 27586 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2004 12396 2421 12424
rect 2004 12384 2010 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 2409 12387 2467 12393
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6546 12424 6552 12436
rect 6144 12396 6552 12424
rect 6144 12384 6150 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 8478 12424 8484 12436
rect 7432 12396 8484 12424
rect 7432 12384 7438 12396
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 10410 12424 10416 12436
rect 8904 12396 10416 12424
rect 8904 12384 8910 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11388 12396 14044 12424
rect 11388 12384 11394 12396
rect 7668 12328 9628 12356
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 4617 12291 4675 12297
rect 4617 12288 4629 12291
rect 2924 12260 4629 12288
rect 2924 12248 2930 12260
rect 4617 12257 4629 12260
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5040 12260 5457 12288
rect 5040 12248 5046 12260
rect 5445 12257 5457 12260
rect 5491 12288 5503 12291
rect 7668 12288 7696 12328
rect 5491 12260 7696 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 9398 12288 9404 12300
rect 8536 12260 9404 12288
rect 8536 12248 8542 12260
rect 9398 12248 9404 12260
rect 9456 12288 9462 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9456 12260 9505 12288
rect 9456 12248 9462 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9600 12288 9628 12328
rect 9766 12288 9772 12300
rect 9600 12260 9772 12288
rect 9493 12251 9551 12257
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10318 12288 10324 12300
rect 9916 12260 10324 12288
rect 9916 12248 9922 12260
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 11606 12248 11612 12300
rect 11664 12288 11670 12300
rect 13722 12288 13728 12300
rect 11664 12260 13728 12288
rect 11664 12248 11670 12260
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 2130 12180 2136 12232
rect 2188 12220 2194 12232
rect 2317 12223 2375 12229
rect 2317 12220 2329 12223
rect 2188 12192 2329 12220
rect 2188 12180 2194 12192
rect 2317 12189 2329 12192
rect 2363 12189 2375 12223
rect 5902 12220 5908 12232
rect 2317 12183 2375 12189
rect 5552 12192 5908 12220
rect 4709 12155 4767 12161
rect 4709 12121 4721 12155
rect 4755 12152 4767 12155
rect 5552 12152 5580 12192
rect 5902 12180 5908 12192
rect 5960 12180 5966 12232
rect 6086 12220 6092 12232
rect 6047 12192 6092 12220
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8386 12220 8392 12232
rect 8168 12192 8392 12220
rect 8168 12180 8174 12192
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11940 12192 11989 12220
rect 11940 12180 11946 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 4755 12124 5580 12152
rect 6365 12155 6423 12161
rect 4755 12121 4767 12124
rect 4709 12115 4767 12121
rect 6365 12121 6377 12155
rect 6411 12121 6423 12155
rect 6365 12115 6423 12121
rect 6380 12084 6408 12115
rect 6914 12112 6920 12164
rect 6972 12112 6978 12164
rect 9769 12155 9827 12161
rect 7760 12124 9720 12152
rect 7760 12084 7788 12124
rect 6380 12056 7788 12084
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8478 12084 8484 12096
rect 7892 12056 7937 12084
rect 8439 12056 8484 12084
rect 7892 12044 7898 12056
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9692 12084 9720 12124
rect 9769 12121 9781 12155
rect 9815 12152 9827 12155
rect 9858 12152 9864 12164
rect 9815 12124 9864 12152
rect 9815 12121 9827 12124
rect 9769 12115 9827 12121
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10226 12112 10232 12164
rect 10284 12112 10290 12164
rect 11790 12112 11796 12164
rect 11848 12152 11854 12164
rect 12253 12155 12311 12161
rect 12253 12152 12265 12155
rect 11848 12124 12265 12152
rect 11848 12112 11854 12124
rect 12253 12121 12265 12124
rect 12299 12121 12311 12155
rect 12253 12115 12311 12121
rect 12342 12112 12348 12164
rect 12400 12152 12406 12164
rect 13906 12152 13912 12164
rect 12400 12124 12742 12152
rect 13648 12124 13912 12152
rect 12400 12112 12406 12124
rect 11054 12084 11060 12096
rect 9692 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11241 12087 11299 12093
rect 11241 12053 11253 12087
rect 11287 12084 11299 12087
rect 11330 12084 11336 12096
rect 11287 12056 11336 12084
rect 11287 12053 11299 12056
rect 11241 12047 11299 12053
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 11974 12044 11980 12096
rect 12032 12084 12038 12096
rect 13648 12084 13676 12124
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 14016 12152 14044 12396
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 15914 12427 15972 12433
rect 15914 12424 15926 12427
rect 14240 12396 15926 12424
rect 14240 12384 14246 12396
rect 15914 12393 15926 12396
rect 15960 12424 15972 12427
rect 16298 12424 16304 12436
rect 15960 12396 16304 12424
rect 15960 12393 15972 12396
rect 15914 12387 15972 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 23750 12424 23756 12436
rect 17236 12396 21128 12424
rect 14090 12316 14096 12368
rect 14148 12356 14154 12368
rect 14734 12356 14740 12368
rect 14148 12328 14740 12356
rect 14148 12316 14154 12328
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 15488 12328 15792 12356
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 15488 12220 15516 12328
rect 15654 12288 15660 12300
rect 15615 12260 15660 12288
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15764 12288 15792 12328
rect 16666 12288 16672 12300
rect 15764 12260 16672 12288
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 14783 12192 15516 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 15013 12155 15071 12161
rect 15013 12152 15025 12155
rect 14016 12124 15025 12152
rect 15013 12121 15025 12124
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 12032 12056 13676 12084
rect 15028 12084 15056 12115
rect 16390 12112 16396 12164
rect 16448 12112 16454 12164
rect 15194 12084 15200 12096
rect 15028 12056 15200 12084
rect 12032 12044 12038 12056
rect 15194 12044 15200 12056
rect 15252 12084 15258 12096
rect 17236 12084 17264 12396
rect 21100 12368 21128 12396
rect 21284 12396 23756 12424
rect 21284 12368 21312 12396
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 27065 12427 27123 12433
rect 27065 12393 27077 12427
rect 27111 12424 27123 12427
rect 27338 12424 27344 12436
rect 27111 12396 27344 12424
rect 27111 12393 27123 12396
rect 27065 12387 27123 12393
rect 27338 12384 27344 12396
rect 27396 12384 27402 12436
rect 28353 12427 28411 12433
rect 28353 12393 28365 12427
rect 28399 12424 28411 12427
rect 28994 12424 29000 12436
rect 28399 12396 29000 12424
rect 28399 12393 28411 12396
rect 28353 12387 28411 12393
rect 28994 12384 29000 12396
rect 29052 12384 29058 12436
rect 17405 12359 17463 12365
rect 17405 12325 17417 12359
rect 17451 12356 17463 12359
rect 19426 12356 19432 12368
rect 17451 12328 19432 12356
rect 17451 12325 17463 12328
rect 17405 12319 17463 12325
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 21082 12316 21088 12368
rect 21140 12316 21146 12368
rect 21266 12316 21272 12368
rect 21324 12316 21330 12368
rect 22002 12316 22008 12368
rect 22060 12356 22066 12368
rect 22060 12328 24624 12356
rect 22060 12316 22066 12328
rect 22281 12291 22339 12297
rect 18432 12260 21128 12288
rect 18432 12229 18460 12260
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 18509 12155 18567 12161
rect 18509 12121 18521 12155
rect 18555 12152 18567 12155
rect 18598 12152 18604 12164
rect 18555 12124 18604 12152
rect 18555 12121 18567 12124
rect 18509 12115 18567 12121
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 15252 12056 17264 12084
rect 15252 12044 15258 12056
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 18874 12084 18880 12096
rect 18380 12056 18880 12084
rect 18380 12044 18386 12056
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19536 12084 19564 12183
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 19797 12155 19855 12161
rect 19797 12152 19809 12155
rect 19760 12124 19809 12152
rect 19760 12112 19766 12124
rect 19797 12121 19809 12124
rect 19843 12121 19855 12155
rect 19797 12115 19855 12121
rect 19300 12056 19564 12084
rect 19812 12084 19840 12115
rect 20806 12112 20812 12164
rect 20864 12112 20870 12164
rect 20530 12084 20536 12096
rect 19812 12056 20536 12084
rect 19300 12044 19306 12056
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 20714 12044 20720 12096
rect 20772 12084 20778 12096
rect 21100 12084 21128 12260
rect 22281 12257 22293 12291
rect 22327 12288 22339 12291
rect 22370 12288 22376 12300
rect 22327 12260 22376 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 23014 12248 23020 12300
rect 23072 12288 23078 12300
rect 23072 12260 23244 12288
rect 23072 12248 23078 12260
rect 23216 12232 23244 12260
rect 22922 12180 22928 12232
rect 22980 12220 22986 12232
rect 22980 12192 23025 12220
rect 22980 12180 22986 12192
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 23290 12180 23296 12232
rect 23348 12220 23354 12232
rect 24596 12229 24624 12328
rect 27614 12288 27620 12300
rect 27575 12260 27620 12288
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 30834 12288 30840 12300
rect 30795 12260 30840 12288
rect 30834 12248 30840 12260
rect 30892 12248 30898 12300
rect 23385 12223 23443 12229
rect 23385 12220 23397 12223
rect 23348 12192 23397 12220
rect 23348 12180 23354 12192
rect 23385 12189 23397 12192
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24946 12180 24952 12232
rect 25004 12220 25010 12232
rect 26145 12223 26203 12229
rect 26145 12220 26157 12223
rect 25004 12192 26157 12220
rect 25004 12180 25010 12192
rect 26145 12189 26157 12192
rect 26191 12189 26203 12223
rect 26145 12183 26203 12189
rect 26878 12180 26884 12232
rect 26936 12220 26942 12232
rect 26973 12223 27031 12229
rect 26973 12220 26985 12223
rect 26936 12192 26985 12220
rect 26936 12180 26942 12192
rect 26973 12189 26985 12192
rect 27019 12189 27031 12223
rect 28258 12220 28264 12232
rect 28219 12192 28264 12220
rect 26973 12183 27031 12189
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 22373 12155 22431 12161
rect 22373 12121 22385 12155
rect 22419 12152 22431 12155
rect 24673 12155 24731 12161
rect 24673 12152 24685 12155
rect 22419 12124 24685 12152
rect 22419 12121 22431 12124
rect 22373 12115 22431 12121
rect 24673 12121 24685 12124
rect 24719 12121 24731 12155
rect 29822 12152 29828 12164
rect 29783 12124 29828 12152
rect 24673 12115 24731 12121
rect 29822 12112 29828 12124
rect 29880 12112 29886 12164
rect 29917 12155 29975 12161
rect 29917 12121 29929 12155
rect 29963 12121 29975 12155
rect 29917 12115 29975 12121
rect 21266 12084 21272 12096
rect 20772 12056 21128 12084
rect 21227 12056 21272 12084
rect 20772 12044 20778 12056
rect 21266 12044 21272 12056
rect 21324 12084 21330 12096
rect 21634 12084 21640 12096
rect 21324 12056 21640 12084
rect 21324 12044 21330 12056
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 23014 12044 23020 12096
rect 23072 12084 23078 12096
rect 23477 12087 23535 12093
rect 23477 12084 23489 12087
rect 23072 12056 23489 12084
rect 23072 12044 23078 12056
rect 23477 12053 23489 12056
rect 23523 12053 23535 12087
rect 23477 12047 23535 12053
rect 26237 12087 26295 12093
rect 26237 12053 26249 12087
rect 26283 12084 26295 12087
rect 29932 12084 29960 12115
rect 26283 12056 29960 12084
rect 26283 12053 26295 12056
rect 26237 12047 26295 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2774 11880 2780 11892
rect 1627 11852 2780 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11849 3295 11883
rect 3237 11843 3295 11849
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 11330 11880 11336 11892
rect 4663 11852 11336 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 2498 11772 2504 11824
rect 2556 11812 2562 11824
rect 3252 11812 3280 11843
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 16298 11880 16304 11892
rect 12084 11852 14320 11880
rect 16259 11852 16304 11880
rect 2556 11784 3280 11812
rect 5261 11815 5319 11821
rect 2556 11772 2562 11784
rect 5261 11781 5273 11815
rect 5307 11812 5319 11815
rect 6822 11812 6828 11824
rect 5307 11784 6828 11812
rect 5307 11781 5319 11784
rect 5261 11775 5319 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 8110 11772 8116 11824
rect 8168 11772 8174 11824
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 10229 11815 10287 11821
rect 10229 11812 10241 11815
rect 9088 11784 10241 11812
rect 9088 11772 9094 11784
rect 10229 11781 10241 11784
rect 10275 11781 10287 11815
rect 10229 11775 10287 11781
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 11882 11812 11888 11824
rect 11296 11784 11888 11812
rect 11296 11772 11302 11784
rect 11882 11772 11888 11784
rect 11940 11772 11946 11824
rect 1762 11744 1768 11756
rect 1723 11716 1768 11744
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 3418 11744 3424 11756
rect 3379 11716 3424 11744
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 4062 11744 4068 11756
rect 4023 11716 4068 11744
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 1578 11568 1584 11620
rect 1636 11608 1642 11620
rect 3881 11611 3939 11617
rect 3881 11608 3893 11611
rect 1636 11580 3893 11608
rect 1636 11568 1642 11580
rect 3881 11577 3893 11580
rect 3927 11577 3939 11611
rect 4540 11608 4568 11707
rect 5184 11676 5212 11707
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5684 11716 5825 11744
rect 5684 11704 5690 11716
rect 5813 11713 5825 11716
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 7006 11744 7012 11756
rect 6779 11716 7012 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7374 11744 7380 11756
rect 7335 11716 7380 11744
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 12084 11753 12112 11852
rect 14292 11824 14320 11852
rect 16298 11840 16304 11852
rect 16356 11840 16362 11892
rect 21266 11880 21272 11892
rect 18524 11852 21272 11880
rect 12342 11772 12348 11824
rect 12400 11812 12406 11824
rect 12618 11812 12624 11824
rect 12400 11784 12624 11812
rect 12400 11772 12406 11784
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 12802 11772 12808 11824
rect 12860 11772 12866 11824
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 13872 11784 13952 11812
rect 13872 11772 13878 11784
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11713 12127 11747
rect 13924 11744 13952 11784
rect 14274 11772 14280 11824
rect 14332 11812 14338 11824
rect 18524 11821 18552 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 22094 11880 22100 11892
rect 21508 11852 22100 11880
rect 21508 11840 21514 11852
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 22572 11852 23152 11880
rect 18509 11815 18567 11821
rect 14332 11784 14596 11812
rect 14332 11772 14338 11784
rect 14568 11756 14596 11784
rect 18509 11781 18521 11815
rect 18555 11781 18567 11815
rect 18509 11775 18567 11781
rect 19518 11772 19524 11824
rect 19576 11772 19582 11824
rect 20901 11815 20959 11821
rect 20901 11781 20913 11815
rect 20947 11812 20959 11815
rect 22281 11815 22339 11821
rect 22281 11812 22293 11815
rect 20947 11784 22293 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 22281 11781 22293 11784
rect 22327 11781 22339 11815
rect 22281 11775 22339 11781
rect 14366 11744 14372 11756
rect 13924 11716 14372 11744
rect 12069 11707 12127 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14550 11744 14556 11756
rect 14511 11716 14556 11744
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 5994 11676 6000 11688
rect 5184 11648 6000 11676
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 7190 11676 7196 11688
rect 6656 11648 7196 11676
rect 5626 11608 5632 11620
rect 4540 11580 5632 11608
rect 3881 11571 3939 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 5905 11611 5963 11617
rect 5905 11577 5917 11611
rect 5951 11608 5963 11611
rect 6656 11608 6684 11648
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8294 11676 8300 11688
rect 7699 11648 8300 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 11054 11676 11060 11688
rect 10183 11648 11060 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11645 11207 11679
rect 11149 11639 11207 11645
rect 5951 11580 6684 11608
rect 5951 11577 5963 11580
rect 5905 11571 5963 11577
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 11164 11608 11192 11639
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 12345 11679 12403 11685
rect 11756 11648 12112 11676
rect 11756 11636 11762 11648
rect 12084 11620 12112 11648
rect 12345 11645 12357 11679
rect 12391 11676 12403 11679
rect 13078 11676 13084 11688
rect 12391 11648 13084 11676
rect 12391 11645 12403 11648
rect 12345 11639 12403 11645
rect 13078 11636 13084 11648
rect 13136 11676 13142 11688
rect 13814 11676 13820 11688
rect 13136 11648 13820 11676
rect 13136 11636 13142 11648
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 11882 11608 11888 11620
rect 9272 11580 11888 11608
rect 9272 11568 9278 11580
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 12066 11568 12072 11620
rect 12124 11568 12130 11620
rect 14108 11608 14136 11639
rect 14182 11636 14188 11688
rect 14240 11676 14246 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 14240 11648 14841 11676
rect 14240 11636 14246 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 14550 11608 14556 11620
rect 14108 11580 14556 11608
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7650 11540 7656 11552
rect 6871 11512 7656 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 9088 11512 9137 11540
rect 9088 11500 9094 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9125 11503 9183 11509
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 15948 11540 15976 11730
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16724 11716 16865 11744
rect 16724 11704 16730 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 18046 11704 18052 11756
rect 18104 11744 18110 11756
rect 18233 11747 18291 11753
rect 18233 11744 18245 11747
rect 18104 11716 18245 11744
rect 18104 11704 18110 11716
rect 18233 11713 18245 11716
rect 18279 11713 18291 11747
rect 22186 11744 22192 11756
rect 22147 11716 22192 11744
rect 18233 11707 18291 11713
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 17034 11676 17040 11688
rect 16995 11648 17040 11676
rect 17034 11636 17040 11648
rect 17092 11676 17098 11688
rect 18506 11676 18512 11688
rect 17092 11648 18512 11676
rect 17092 11636 17098 11648
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 20257 11679 20315 11685
rect 20257 11676 20269 11679
rect 19116 11648 20269 11676
rect 19116 11636 19122 11648
rect 20257 11645 20269 11648
rect 20303 11645 20315 11679
rect 20257 11639 20315 11645
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11676 20867 11679
rect 20898 11676 20904 11688
rect 20855 11648 20904 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 20272 11608 20300 11639
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 21082 11676 21088 11688
rect 21043 11648 21088 11676
rect 21082 11636 21088 11648
rect 21140 11636 21146 11688
rect 22278 11676 22284 11688
rect 21192 11648 22284 11676
rect 21192 11608 21220 11648
rect 22278 11636 22284 11648
rect 22336 11676 22342 11688
rect 22572 11676 22600 11852
rect 23014 11812 23020 11824
rect 22975 11784 23020 11812
rect 23014 11772 23020 11784
rect 23072 11772 23078 11824
rect 23124 11812 23152 11852
rect 23382 11840 23388 11892
rect 23440 11880 23446 11892
rect 25406 11880 25412 11892
rect 23440 11852 25412 11880
rect 23440 11840 23446 11852
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 25777 11883 25835 11889
rect 25777 11849 25789 11883
rect 25823 11880 25835 11883
rect 26786 11880 26792 11892
rect 25823 11852 26792 11880
rect 25823 11849 25835 11852
rect 25777 11843 25835 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 28258 11880 28264 11892
rect 26896 11852 28264 11880
rect 26896 11812 26924 11852
rect 28258 11840 28264 11852
rect 28316 11840 28322 11892
rect 35713 11883 35771 11889
rect 35713 11849 35725 11883
rect 35759 11880 35771 11883
rect 36906 11880 36912 11892
rect 35759 11852 36912 11880
rect 35759 11849 35771 11852
rect 35713 11843 35771 11849
rect 36906 11840 36912 11852
rect 36964 11840 36970 11892
rect 27246 11812 27252 11824
rect 23124 11784 26924 11812
rect 27207 11784 27252 11812
rect 27246 11772 27252 11784
rect 27304 11772 27310 11824
rect 27338 11772 27344 11824
rect 27396 11812 27402 11824
rect 27396 11784 27441 11812
rect 27396 11772 27402 11784
rect 24394 11744 24400 11756
rect 24355 11716 24400 11744
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11744 25099 11747
rect 25130 11744 25136 11756
rect 25087 11716 25136 11744
rect 25087 11713 25099 11716
rect 25041 11707 25099 11713
rect 25130 11704 25136 11716
rect 25188 11704 25194 11756
rect 25682 11744 25688 11756
rect 25643 11716 25688 11744
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 33226 11704 33232 11756
rect 33284 11744 33290 11756
rect 35897 11747 35955 11753
rect 35897 11744 35909 11747
rect 33284 11716 35909 11744
rect 33284 11704 33290 11716
rect 35897 11713 35909 11716
rect 35943 11713 35955 11747
rect 35897 11707 35955 11713
rect 22336 11648 22600 11676
rect 22925 11679 22983 11685
rect 22336 11636 22342 11648
rect 22925 11645 22937 11679
rect 22971 11676 22983 11679
rect 23106 11676 23112 11688
rect 22971 11648 23112 11676
rect 22971 11645 22983 11648
rect 22925 11639 22983 11645
rect 23106 11636 23112 11648
rect 23164 11636 23170 11688
rect 23937 11679 23995 11685
rect 23937 11645 23949 11679
rect 23983 11676 23995 11679
rect 26142 11676 26148 11688
rect 23983 11648 26148 11676
rect 23983 11645 23995 11648
rect 23937 11639 23995 11645
rect 26142 11636 26148 11648
rect 26200 11636 26206 11688
rect 27430 11636 27436 11688
rect 27488 11676 27494 11688
rect 27525 11679 27583 11685
rect 27525 11676 27537 11679
rect 27488 11648 27537 11676
rect 27488 11636 27494 11648
rect 27525 11645 27537 11648
rect 27571 11676 27583 11679
rect 27614 11676 27620 11688
rect 27571 11648 27620 11676
rect 27571 11645 27583 11648
rect 27525 11639 27583 11645
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 24670 11608 24676 11620
rect 20272 11580 21220 11608
rect 23400 11580 24676 11608
rect 9548 11512 15976 11540
rect 9548 11500 9554 11512
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 21266 11540 21272 11552
rect 16172 11512 21272 11540
rect 16172 11500 16178 11512
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 22370 11500 22376 11552
rect 22428 11540 22434 11552
rect 23400 11540 23428 11580
rect 24670 11568 24676 11580
rect 24728 11568 24734 11620
rect 25133 11611 25191 11617
rect 25133 11577 25145 11611
rect 25179 11608 25191 11611
rect 26326 11608 26332 11620
rect 25179 11580 26332 11608
rect 25179 11577 25191 11580
rect 25133 11571 25191 11577
rect 26326 11568 26332 11580
rect 26384 11568 26390 11620
rect 22428 11512 23428 11540
rect 22428 11500 22434 11512
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 24489 11543 24547 11549
rect 24489 11540 24501 11543
rect 23532 11512 24501 11540
rect 23532 11500 23538 11512
rect 24489 11509 24501 11512
rect 24535 11509 24547 11543
rect 24489 11503 24547 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 3476 11308 4261 11336
rect 3476 11296 3482 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 6822 11336 6828 11348
rect 5132 11308 6828 11336
rect 5132 11296 5138 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7558 11336 7564 11348
rect 6972 11308 7564 11336
rect 6972 11296 6978 11308
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8352 11308 8585 11336
rect 8352 11296 8358 11308
rect 8573 11305 8585 11308
rect 8619 11336 8631 11339
rect 9306 11336 9312 11348
rect 8619 11308 9312 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 12434 11336 12440 11348
rect 9447 11308 12440 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 13446 11336 13452 11348
rect 13407 11308 13452 11336
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 16850 11345 16856 11348
rect 16840 11339 16856 11345
rect 16840 11336 16852 11339
rect 16763 11308 16852 11336
rect 16840 11305 16852 11308
rect 16908 11336 16914 11348
rect 17494 11336 17500 11348
rect 16908 11308 17500 11336
rect 16840 11299 16856 11305
rect 16850 11296 16856 11299
rect 16908 11296 16914 11308
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18322 11336 18328 11348
rect 18283 11308 18328 11336
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 19968 11339 20026 11345
rect 19968 11305 19980 11339
rect 20014 11336 20026 11339
rect 21266 11336 21272 11348
rect 20014 11308 21272 11336
rect 20014 11305 20026 11308
rect 19968 11299 20026 11305
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 21358 11296 21364 11348
rect 21416 11336 21422 11348
rect 21453 11339 21511 11345
rect 21453 11336 21465 11339
rect 21416 11308 21465 11336
rect 21416 11296 21422 11308
rect 21453 11305 21465 11308
rect 21499 11305 21511 11339
rect 21453 11299 21511 11305
rect 21542 11296 21548 11348
rect 21600 11336 21606 11348
rect 22002 11336 22008 11348
rect 21600 11308 22008 11336
rect 21600 11296 21606 11308
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22152 11308 24532 11336
rect 22152 11296 22158 11308
rect 8754 11228 8760 11280
rect 8812 11268 8818 11280
rect 10045 11271 10103 11277
rect 10045 11268 10057 11271
rect 8812 11240 10057 11268
rect 8812 11228 8818 11240
rect 10045 11237 10057 11240
rect 10091 11237 10103 11271
rect 10045 11231 10103 11237
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 12986 11268 12992 11280
rect 11940 11240 12992 11268
rect 11940 11228 11946 11240
rect 12986 11228 12992 11240
rect 13044 11228 13050 11280
rect 18046 11228 18052 11280
rect 18104 11268 18110 11280
rect 19242 11268 19248 11280
rect 18104 11240 19248 11268
rect 18104 11228 18110 11240
rect 19242 11228 19248 11240
rect 19300 11268 19306 11280
rect 19300 11240 19748 11268
rect 19300 11228 19306 11240
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11200 1915 11203
rect 2682 11200 2688 11212
rect 1903 11172 2688 11200
rect 1903 11169 1915 11172
rect 1857 11163 1915 11169
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 9214 11200 9220 11212
rect 4172 11172 9220 11200
rect 1578 11132 1584 11144
rect 1539 11104 1584 11132
rect 1578 11092 1584 11104
rect 1636 11092 1642 11144
rect 4172 11141 4200 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9398 11160 9404 11212
rect 9456 11200 9462 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 9456 11172 10609 11200
rect 9456 11160 9462 11172
rect 10597 11169 10609 11172
rect 10643 11200 10655 11203
rect 11238 11200 11244 11212
rect 10643 11172 11244 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12621 11203 12679 11209
rect 12621 11200 12633 11203
rect 11664 11172 12633 11200
rect 11664 11160 11670 11172
rect 12621 11169 12633 11172
rect 12667 11200 12679 11203
rect 13170 11200 13176 11212
rect 12667 11172 13176 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 14274 11200 14280 11212
rect 14235 11172 14280 11200
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 14550 11200 14556 11212
rect 14511 11172 14556 11200
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 15930 11160 15936 11212
rect 15988 11200 15994 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15988 11172 16037 11200
rect 15988 11160 15994 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 18064 11200 18092 11228
rect 19720 11209 19748 11240
rect 16623 11172 18092 11200
rect 19705 11203 19763 11209
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19751 11172 21956 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 4982 11132 4988 11144
rect 4847 11104 4988 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 6144 11104 6193 11132
rect 6144 11092 6150 11104
rect 6181 11101 6193 11104
rect 6227 11132 6239 11135
rect 6822 11132 6828 11144
rect 6227 11104 6828 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 9309 11135 9367 11141
rect 8588 11104 9168 11132
rect 4893 11067 4951 11073
rect 4893 11033 4905 11067
rect 4939 11064 4951 11067
rect 5445 11067 5503 11073
rect 4939 11036 5304 11064
rect 4939 11033 4951 11036
rect 4893 11027 4951 11033
rect 5276 11008 5304 11036
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 5534 11064 5540 11076
rect 5491 11036 5540 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 7064 11036 7113 11064
rect 7064 11024 7070 11036
rect 7101 11033 7113 11036
rect 7147 11033 7159 11067
rect 7101 11027 7159 11033
rect 7190 11024 7196 11076
rect 7248 11064 7254 11076
rect 7248 11036 7590 11064
rect 7248 11024 7254 11036
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 2869 10999 2927 11005
rect 2869 10996 2881 10999
rect 2832 10968 2881 10996
rect 2832 10956 2838 10968
rect 2869 10965 2881 10968
rect 2915 10965 2927 10999
rect 2869 10959 2927 10965
rect 5258 10956 5264 11008
rect 5316 10956 5322 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 8588 10996 8616 11104
rect 6512 10968 8616 10996
rect 6512 10956 6518 10968
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 9030 10996 9036 11008
rect 8720 10968 9036 10996
rect 8720 10956 8726 10968
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 9140 10996 9168 11104
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9490 11132 9496 11144
rect 9355 11104 9496 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9640 11104 9965 11132
rect 9640 11092 9646 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13412 11104 13457 11132
rect 13412 11092 13418 11104
rect 21082 11092 21088 11144
rect 21140 11092 21146 11144
rect 21928 11132 21956 11172
rect 22002 11132 22008 11144
rect 21915 11104 22008 11132
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 24504 11132 24532 11308
rect 24670 11296 24676 11348
rect 24728 11336 24734 11348
rect 25590 11336 25596 11348
rect 24728 11308 25596 11336
rect 24728 11296 24734 11308
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 26881 11339 26939 11345
rect 26881 11305 26893 11339
rect 26927 11336 26939 11339
rect 27338 11336 27344 11348
rect 26927 11308 27344 11336
rect 26927 11305 26939 11308
rect 26881 11299 26939 11305
rect 27338 11296 27344 11308
rect 27396 11296 27402 11348
rect 33226 11336 33232 11348
rect 33187 11308 33232 11336
rect 33226 11296 33232 11308
rect 33284 11296 33290 11348
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 24504 11104 24593 11132
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11132 25283 11135
rect 25406 11132 25412 11144
rect 25271 11104 25412 11132
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 25406 11092 25412 11104
rect 25464 11092 25470 11144
rect 26786 11132 26792 11144
rect 26747 11104 26792 11132
rect 26786 11092 26792 11104
rect 26844 11092 26850 11144
rect 29270 11092 29276 11144
rect 29328 11132 29334 11144
rect 33137 11135 33195 11141
rect 33137 11132 33149 11135
rect 29328 11104 33149 11132
rect 29328 11092 29334 11104
rect 33137 11101 33149 11104
rect 33183 11101 33195 11135
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 33137 11095 33195 11101
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 10318 11024 10324 11076
rect 10376 11064 10382 11076
rect 10870 11064 10876 11076
rect 10376 11036 10876 11064
rect 10376 11024 10382 11036
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 11330 11024 11336 11076
rect 11388 11024 11394 11076
rect 12158 11024 12164 11076
rect 12216 11064 12222 11076
rect 12216 11036 15042 11064
rect 12216 11024 12222 11036
rect 17310 11024 17316 11076
rect 17368 11024 17374 11076
rect 19058 11024 19064 11076
rect 19116 11064 19122 11076
rect 19116 11036 20392 11064
rect 19116 11024 19122 11036
rect 10962 10996 10968 11008
rect 9140 10968 10968 10996
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 17034 10996 17040 11008
rect 14792 10968 17040 10996
rect 14792 10956 14798 10968
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 20364 10996 20392 11036
rect 21284 11036 22232 11064
rect 21284 10996 21312 11036
rect 20364 10968 21312 10996
rect 22204 10996 22232 11036
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22336 11036 22381 11064
rect 22336 11024 22342 11036
rect 22738 11024 22744 11076
rect 22796 11024 22802 11076
rect 25317 11067 25375 11073
rect 25317 11064 25329 11067
rect 23584 11036 25329 11064
rect 23584 10996 23612 11036
rect 25317 11033 25329 11036
rect 25363 11033 25375 11067
rect 25317 11027 25375 11033
rect 23750 10996 23756 11008
rect 22204 10968 23612 10996
rect 23711 10968 23756 10996
rect 23750 10956 23756 10968
rect 23808 10956 23814 11008
rect 23842 10956 23848 11008
rect 23900 10996 23906 11008
rect 24673 10999 24731 11005
rect 24673 10996 24685 10999
rect 23900 10968 24685 10996
rect 23900 10956 23906 10968
rect 24673 10965 24685 10968
rect 24719 10965 24731 10999
rect 24673 10959 24731 10965
rect 38010 10956 38016 11008
rect 38068 10996 38074 11008
rect 38105 10999 38163 11005
rect 38105 10996 38117 10999
rect 38068 10968 38117 10996
rect 38068 10956 38074 10968
rect 38105 10965 38117 10968
rect 38151 10965 38163 10999
rect 38105 10959 38163 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4614 10792 4620 10804
rect 4295 10764 4620 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5810 10792 5816 10804
rect 5307 10764 5816 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 6546 10752 6552 10804
rect 6604 10752 6610 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6730 10792 6736 10804
rect 6687 10764 6736 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 8018 10792 8024 10804
rect 6972 10764 8024 10792
rect 6972 10752 6978 10764
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 12802 10792 12808 10804
rect 12759 10764 12808 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13262 10792 13268 10804
rect 13004 10764 13268 10792
rect 6564 10724 6592 10752
rect 6564 10696 8602 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2774 10656 2780 10668
rect 2731 10628 2780 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 4157 10659 4215 10665
rect 4157 10656 4169 10659
rect 3200 10628 4169 10656
rect 3200 10616 3206 10628
rect 4157 10625 4169 10628
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 5169 10659 5227 10665
rect 5169 10656 5181 10659
rect 4672 10628 5181 10656
rect 4672 10616 4678 10628
rect 5169 10625 5181 10628
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5684 10628 5825 10656
rect 5684 10616 5690 10628
rect 5813 10625 5825 10628
rect 5859 10656 5871 10659
rect 6270 10656 6276 10668
rect 5859 10628 6276 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6270 10616 6276 10628
rect 6328 10656 6334 10668
rect 6454 10656 6460 10668
rect 6328 10628 6460 10656
rect 6328 10616 6334 10628
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6914 10656 6920 10668
rect 6595 10628 6920 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7185 10659 7243 10665
rect 7185 10656 7197 10659
rect 7024 10628 7197 10656
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 1946 10588 1952 10600
rect 1811 10560 1952 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2556 10560 2881 10588
rect 2556 10548 2562 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 7024 10588 7052 10628
rect 7185 10625 7197 10628
rect 7231 10625 7243 10659
rect 7185 10619 7243 10625
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7844 10659 7902 10665
rect 7432 10646 7788 10656
rect 7844 10646 7856 10659
rect 7432 10628 7856 10646
rect 7432 10616 7438 10628
rect 7760 10625 7856 10628
rect 7890 10625 7902 10659
rect 7760 10619 7902 10625
rect 7760 10618 7880 10619
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 9456 10628 10149 10656
rect 9456 10616 9462 10628
rect 10137 10625 10149 10628
rect 10183 10656 10195 10659
rect 10226 10656 10232 10668
rect 10183 10628 10232 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10226 10616 10232 10628
rect 10284 10616 10290 10668
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10560 10628 10793 10656
rect 10560 10616 10566 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 10962 10616 10968 10668
rect 11020 10656 11026 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11020 10628 11805 10656
rect 11020 10616 11026 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 12621 10659 12679 10665
rect 12621 10625 12633 10659
rect 12667 10656 12679 10659
rect 12894 10656 12900 10668
rect 12667 10628 12900 10656
rect 12667 10625 12679 10628
rect 12621 10619 12679 10625
rect 6788 10560 7052 10588
rect 8113 10591 8171 10597
rect 6788 10548 6794 10560
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 11606 10588 11612 10600
rect 8159 10560 11612 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11808 10588 11836 10619
rect 12894 10616 12900 10628
rect 12952 10656 12958 10668
rect 13004 10656 13032 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 13872 10764 15025 10792
rect 13872 10752 13878 10764
rect 15013 10761 15025 10764
rect 15059 10761 15071 10795
rect 15013 10755 15071 10761
rect 16209 10795 16267 10801
rect 16209 10761 16221 10795
rect 16255 10792 16267 10795
rect 17770 10792 17776 10804
rect 16255 10764 17776 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 18601 10795 18659 10801
rect 18601 10761 18613 10795
rect 18647 10792 18659 10795
rect 19334 10792 19340 10804
rect 18647 10764 19340 10792
rect 18647 10761 18659 10764
rect 18601 10755 18659 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 21266 10792 21272 10804
rect 19904 10764 21272 10792
rect 13446 10724 13452 10736
rect 12952 10628 13032 10656
rect 13096 10696 13452 10724
rect 12952 10616 12958 10628
rect 13096 10588 13124 10696
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 14274 10684 14280 10736
rect 14332 10684 14338 10736
rect 16482 10684 16488 10736
rect 16540 10724 16546 10736
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 16540 10696 17141 10724
rect 16540 10684 16546 10696
rect 17129 10693 17141 10696
rect 17175 10693 17187 10727
rect 19150 10724 19156 10736
rect 18354 10696 19156 10724
rect 17129 10687 17187 10693
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 19904 10724 19932 10764
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 22646 10752 22652 10804
rect 22704 10792 22710 10804
rect 26694 10792 26700 10804
rect 22704 10764 26700 10792
rect 22704 10752 22710 10764
rect 26694 10752 26700 10764
rect 26752 10792 26758 10804
rect 26752 10764 27200 10792
rect 26752 10752 26758 10764
rect 21450 10724 21456 10736
rect 19260 10696 19932 10724
rect 20746 10696 21456 10724
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 14752 10628 16129 10656
rect 13262 10588 13268 10600
rect 11808 10560 13124 10588
rect 13223 10560 13268 10588
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 13998 10588 14004 10600
rect 13587 10560 14004 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 10229 10523 10287 10529
rect 9180 10492 9628 10520
rect 9180 10480 9186 10492
rect 9600 10464 9628 10492
rect 10229 10489 10241 10523
rect 10275 10520 10287 10523
rect 12618 10520 12624 10532
rect 10275 10492 12624 10520
rect 10275 10489 10287 10492
rect 10229 10483 10287 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 2096 10424 2237 10452
rect 2096 10412 2102 10424
rect 2225 10421 2237 10424
rect 2271 10452 2283 10455
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2271 10424 3065 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 5902 10452 5908 10464
rect 5863 10424 5908 10452
rect 3053 10415 3111 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7190 10452 7196 10464
rect 6972 10424 7196 10452
rect 6972 10412 6978 10424
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7558 10452 7564 10464
rect 7331 10424 7564 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8294 10452 8300 10464
rect 8260 10424 8300 10452
rect 8260 10412 8266 10424
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 9398 10452 9404 10464
rect 8352 10424 9404 10452
rect 8352 10412 8358 10424
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 10870 10452 10876 10464
rect 10831 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11664 10424 11897 10452
rect 11664 10412 11670 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 11885 10415 11943 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 14752 10452 14780 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 19260 10656 19288 10696
rect 21450 10684 21456 10696
rect 21508 10684 21514 10736
rect 21910 10684 21916 10736
rect 21968 10724 21974 10736
rect 21968 10696 22770 10724
rect 21968 10684 21974 10696
rect 22002 10656 22008 10668
rect 16117 10619 16175 10625
rect 19076 10628 19288 10656
rect 21963 10628 22008 10656
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 15712 10560 16865 10588
rect 15712 10548 15718 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 19076 10588 19104 10628
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 27172 10665 27200 10764
rect 27249 10727 27307 10733
rect 27249 10693 27261 10727
rect 27295 10724 27307 10727
rect 27985 10727 28043 10733
rect 27985 10724 27997 10727
rect 27295 10696 27997 10724
rect 27295 10693 27307 10696
rect 27249 10687 27307 10693
rect 27985 10693 27997 10696
rect 28031 10693 28043 10727
rect 27985 10687 28043 10693
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 37826 10616 37832 10668
rect 37884 10656 37890 10668
rect 38013 10659 38071 10665
rect 38013 10656 38025 10659
rect 37884 10628 38025 10656
rect 37884 10616 37890 10628
rect 38013 10625 38025 10628
rect 38059 10625 38071 10659
rect 38013 10619 38071 10625
rect 19242 10588 19248 10600
rect 17184 10560 19104 10588
rect 19203 10560 19248 10588
rect 17184 10548 17190 10560
rect 19242 10548 19248 10560
rect 19300 10548 19306 10600
rect 19521 10591 19579 10597
rect 19521 10557 19533 10591
rect 19567 10588 19579 10591
rect 20070 10588 20076 10600
rect 19567 10560 20076 10588
rect 19567 10557 19579 10560
rect 19521 10551 19579 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 21174 10548 21180 10600
rect 21232 10588 21238 10600
rect 21269 10591 21327 10597
rect 21269 10588 21281 10591
rect 21232 10560 21281 10588
rect 21232 10548 21238 10560
rect 21269 10557 21281 10560
rect 21315 10557 21327 10591
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 21269 10551 21327 10557
rect 22066 10560 22293 10588
rect 21818 10480 21824 10532
rect 21876 10520 21882 10532
rect 22066 10520 22094 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 22922 10548 22928 10600
rect 22980 10588 22986 10600
rect 22980 10560 23428 10588
rect 22980 10548 22986 10560
rect 23400 10532 23428 10560
rect 23566 10548 23572 10600
rect 23624 10588 23630 10600
rect 23753 10591 23811 10597
rect 23753 10588 23765 10591
rect 23624 10560 23765 10588
rect 23624 10548 23630 10560
rect 23753 10557 23765 10560
rect 23799 10557 23811 10591
rect 23753 10551 23811 10557
rect 27893 10591 27951 10597
rect 27893 10557 27905 10591
rect 27939 10588 27951 10591
rect 28074 10588 28080 10600
rect 27939 10560 28080 10588
rect 27939 10557 27951 10560
rect 27893 10551 27951 10557
rect 28074 10548 28080 10560
rect 28132 10588 28138 10600
rect 28534 10588 28540 10600
rect 28132 10560 28540 10588
rect 28132 10548 28138 10560
rect 28534 10548 28540 10560
rect 28592 10548 28598 10600
rect 21876 10492 22094 10520
rect 21876 10480 21882 10492
rect 23382 10480 23388 10532
rect 23440 10480 23446 10532
rect 28442 10520 28448 10532
rect 23676 10492 28448 10520
rect 12768 10424 14780 10452
rect 12768 10412 12774 10424
rect 16482 10412 16488 10464
rect 16540 10452 16546 10464
rect 17126 10452 17132 10464
rect 16540 10424 17132 10452
rect 16540 10412 16546 10424
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17586 10412 17592 10464
rect 17644 10452 17650 10464
rect 23676 10452 23704 10492
rect 28442 10480 28448 10492
rect 28500 10480 28506 10532
rect 38194 10452 38200 10464
rect 17644 10424 23704 10452
rect 38155 10424 38200 10452
rect 17644 10412 17650 10424
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 8573 10251 8631 10257
rect 6319 10220 8524 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 8496 10180 8524 10220
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 10042 10248 10048 10260
rect 8619 10220 10048 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 23750 10248 23756 10260
rect 11164 10220 23756 10248
rect 8496 10152 8616 10180
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 8294 10112 8300 10124
rect 5675 10084 8300 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 1946 10044 1952 10056
rect 1903 10016 1952 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2682 10044 2688 10056
rect 2643 10016 2688 10044
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3329 10047 3387 10053
rect 3329 10044 3341 10047
rect 3016 10016 3341 10044
rect 3016 10004 3022 10016
rect 3329 10013 3341 10016
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3786 10004 3792 10056
rect 3844 10044 3850 10056
rect 4062 10044 4068 10056
rect 3844 10016 4068 10044
rect 3844 10004 3850 10016
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4890 10044 4896 10056
rect 4203 10016 4896 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5583 10016 6193 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 6181 10013 6193 10016
rect 6227 10044 6239 10047
rect 6270 10044 6276 10056
rect 6227 10016 6276 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7101 9979 7159 9985
rect 7101 9945 7113 9979
rect 7147 9945 7159 9979
rect 7101 9939 7159 9945
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 3973 9911 4031 9917
rect 3973 9908 3985 9911
rect 3844 9880 3985 9908
rect 3844 9868 3850 9880
rect 3973 9877 3985 9880
rect 4019 9877 4031 9911
rect 3973 9871 4031 9877
rect 4982 9868 4988 9920
rect 5040 9908 5046 9920
rect 5258 9908 5264 9920
rect 5040 9880 5264 9908
rect 5040 9868 5046 9880
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 7116 9908 7144 9939
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 7374 9976 7380 9988
rect 7248 9948 7380 9976
rect 7248 9936 7254 9948
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 7558 9936 7564 9988
rect 7616 9936 7622 9988
rect 8588 9976 8616 10152
rect 9953 10115 10011 10121
rect 9953 10081 9965 10115
rect 9999 10112 10011 10115
rect 11164 10112 11192 10220
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 37826 10248 37832 10260
rect 37787 10220 37832 10248
rect 37826 10208 37832 10220
rect 37884 10208 37890 10260
rect 11238 10140 11244 10192
rect 11296 10180 11302 10192
rect 11425 10183 11483 10189
rect 11425 10180 11437 10183
rect 11296 10152 11437 10180
rect 11296 10140 11302 10152
rect 11425 10149 11437 10152
rect 11471 10149 11483 10183
rect 11425 10143 11483 10149
rect 13262 10140 13268 10192
rect 13320 10180 13326 10192
rect 13320 10152 14872 10180
rect 13320 10140 13326 10152
rect 9999 10084 11192 10112
rect 11885 10115 11943 10121
rect 9999 10081 10011 10084
rect 9953 10075 10011 10081
rect 11885 10081 11897 10115
rect 11931 10112 11943 10115
rect 13280 10112 13308 10140
rect 11931 10084 13308 10112
rect 14844 10112 14872 10152
rect 15194 10140 15200 10192
rect 15252 10180 15258 10192
rect 17681 10183 17739 10189
rect 15252 10152 16068 10180
rect 15252 10140 15258 10152
rect 15013 10115 15071 10121
rect 15013 10112 15025 10115
rect 14844 10084 15025 10112
rect 11931 10081 11943 10084
rect 11885 10075 11943 10081
rect 15013 10081 15025 10084
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 15712 10084 15945 10112
rect 15712 10072 15718 10084
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 16040 10112 16068 10152
rect 17681 10149 17693 10183
rect 17727 10180 17739 10183
rect 18138 10180 18144 10192
rect 17727 10152 18144 10180
rect 17727 10149 17739 10152
rect 17681 10143 17739 10149
rect 18138 10140 18144 10152
rect 18196 10140 18202 10192
rect 18233 10183 18291 10189
rect 18233 10149 18245 10183
rect 18279 10180 18291 10183
rect 19426 10180 19432 10192
rect 18279 10152 19432 10180
rect 18279 10149 18291 10152
rect 18233 10143 18291 10149
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 21266 10140 21272 10192
rect 21324 10180 21330 10192
rect 21361 10183 21419 10189
rect 21361 10180 21373 10183
rect 21324 10152 21373 10180
rect 21324 10140 21330 10152
rect 21361 10149 21373 10152
rect 21407 10149 21419 10183
rect 21361 10143 21419 10149
rect 23198 10140 23204 10192
rect 23256 10180 23262 10192
rect 23256 10152 23336 10180
rect 23256 10140 23262 10152
rect 18156 10112 18184 10140
rect 19889 10115 19947 10121
rect 19889 10112 19901 10115
rect 16040 10084 17448 10112
rect 18156 10084 19901 10112
rect 15933 10075 15991 10081
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 17420 10044 17448 10084
rect 19889 10081 19901 10084
rect 19935 10081 19947 10115
rect 23106 10112 23112 10124
rect 19889 10075 19947 10081
rect 21008 10084 23112 10112
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 13780 10016 15240 10044
rect 17420 10016 18153 10044
rect 13780 10004 13786 10016
rect 9950 9976 9956 9988
rect 8588 9948 9956 9976
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 12161 9979 12219 9985
rect 10060 9948 10442 9976
rect 7926 9908 7932 9920
rect 7116 9880 7932 9908
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 10060 9908 10088 9948
rect 12161 9945 12173 9979
rect 12207 9976 12219 9979
rect 12207 9948 12434 9976
rect 12207 9945 12219 9948
rect 12161 9939 12219 9945
rect 8168 9880 10088 9908
rect 12406 9908 12434 9948
rect 12618 9936 12624 9988
rect 12676 9936 12682 9988
rect 14277 9979 14335 9985
rect 14277 9945 14289 9979
rect 14323 9976 14335 9979
rect 14734 9976 14740 9988
rect 14323 9948 14740 9976
rect 14323 9945 14335 9948
rect 14277 9939 14335 9945
rect 14734 9936 14740 9948
rect 14792 9976 14798 9988
rect 15102 9976 15108 9988
rect 14792 9948 15108 9976
rect 14792 9936 14798 9948
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 15212 9976 15240 10016
rect 18141 10013 18153 10016
rect 18187 10044 18199 10047
rect 18690 10044 18696 10056
rect 18187 10016 18696 10044
rect 18187 10013 18199 10016
rect 18141 10007 18199 10013
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19484 10016 19625 10044
rect 19484 10004 19490 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 21008 10030 21036 10084
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 23308 10121 23336 10152
rect 28442 10140 28448 10192
rect 28500 10180 28506 10192
rect 30377 10183 30435 10189
rect 30377 10180 30389 10183
rect 28500 10152 30389 10180
rect 28500 10140 28506 10152
rect 30377 10149 30389 10152
rect 30423 10149 30435 10183
rect 30377 10143 30435 10149
rect 23293 10115 23351 10121
rect 23293 10081 23305 10115
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23440 10084 23980 10112
rect 23440 10072 23446 10084
rect 19613 10007 19671 10013
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 22557 10047 22615 10053
rect 22557 10044 22569 10047
rect 22060 10016 22569 10044
rect 22060 10004 22066 10016
rect 22557 10013 22569 10016
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 15212 9948 16221 9976
rect 16209 9945 16221 9948
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 16666 9936 16672 9988
rect 16724 9936 16730 9988
rect 21821 9979 21879 9985
rect 21821 9945 21833 9979
rect 21867 9976 21879 9979
rect 21910 9976 21916 9988
rect 21867 9948 21916 9976
rect 21867 9945 21879 9948
rect 21821 9939 21879 9945
rect 21910 9936 21916 9948
rect 21968 9936 21974 9988
rect 23385 9979 23443 9985
rect 23385 9945 23397 9979
rect 23431 9976 23443 9979
rect 23750 9976 23756 9988
rect 23431 9948 23756 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 23750 9936 23756 9948
rect 23808 9936 23814 9988
rect 23952 9985 23980 10084
rect 24394 10004 24400 10056
rect 24452 10044 24458 10056
rect 24581 10047 24639 10053
rect 24581 10044 24593 10047
rect 24452 10016 24593 10044
rect 24452 10004 24458 10016
rect 24581 10013 24593 10016
rect 24627 10013 24639 10047
rect 25222 10044 25228 10056
rect 25183 10016 25228 10044
rect 24581 10007 24639 10013
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 38010 10044 38016 10056
rect 37971 10016 38016 10044
rect 38010 10004 38016 10016
rect 38068 10004 38074 10056
rect 23937 9979 23995 9985
rect 23937 9945 23949 9979
rect 23983 9976 23995 9979
rect 23983 9948 27568 9976
rect 23983 9945 23995 9948
rect 23937 9939 23995 9945
rect 12526 9908 12532 9920
rect 12406 9880 12532 9908
rect 8168 9868 8174 9880
rect 12526 9868 12532 9880
rect 12584 9908 12590 9920
rect 13538 9908 13544 9920
rect 12584 9880 13544 9908
rect 12584 9868 12590 9880
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 15286 9908 15292 9920
rect 13679 9880 15292 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 21174 9908 21180 9920
rect 15436 9880 21180 9908
rect 15436 9868 15442 9880
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 23658 9868 23664 9920
rect 23716 9908 23722 9920
rect 24673 9911 24731 9917
rect 24673 9908 24685 9911
rect 23716 9880 24685 9908
rect 23716 9868 23722 9880
rect 24673 9877 24685 9880
rect 24719 9877 24731 9911
rect 24673 9871 24731 9877
rect 24854 9868 24860 9920
rect 24912 9908 24918 9920
rect 25317 9911 25375 9917
rect 25317 9908 25329 9911
rect 24912 9880 25329 9908
rect 24912 9868 24918 9880
rect 25317 9877 25329 9880
rect 25363 9877 25375 9911
rect 27430 9908 27436 9920
rect 27391 9880 27436 9908
rect 25317 9871 25375 9877
rect 27430 9868 27436 9880
rect 27488 9868 27494 9920
rect 27540 9908 27568 9948
rect 29178 9936 29184 9988
rect 29236 9976 29242 9988
rect 29822 9976 29828 9988
rect 29236 9948 29828 9976
rect 29236 9936 29242 9948
rect 29822 9936 29828 9948
rect 29880 9936 29886 9988
rect 29914 9936 29920 9988
rect 29972 9976 29978 9988
rect 29972 9948 30017 9976
rect 29972 9936 29978 9948
rect 30006 9908 30012 9920
rect 27540 9880 30012 9908
rect 30006 9868 30012 9880
rect 30064 9868 30070 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2682 9704 2688 9716
rect 1903 9676 2688 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 4908 9676 5856 9704
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 2004 9608 3004 9636
rect 2004 9596 2010 9608
rect 2056 9577 2084 9608
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2774 9568 2780 9580
rect 2547 9540 2780 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 1854 9460 1860 9512
rect 1912 9500 1918 9512
rect 2593 9503 2651 9509
rect 2593 9500 2605 9503
rect 1912 9472 2605 9500
rect 1912 9460 1918 9472
rect 2593 9469 2605 9472
rect 2639 9469 2651 9503
rect 2976 9500 3004 9608
rect 3050 9596 3056 9648
rect 3108 9636 3114 9648
rect 4908 9636 4936 9676
rect 3108 9608 4936 9636
rect 3108 9596 3114 9608
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 5828 9636 5856 9676
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 9214 9704 9220 9716
rect 6328 9676 9220 9704
rect 6328 9664 6334 9676
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 9674 9704 9680 9716
rect 9416 9676 9680 9704
rect 5828 9608 7958 9636
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 6822 9568 6828 9580
rect 5920 9540 6828 9568
rect 3326 9500 3332 9512
rect 2976 9472 3332 9500
rect 2593 9463 2651 9469
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4982 9500 4988 9512
rect 4571 9472 4988 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 3234 9364 3240 9376
rect 3195 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 4264 9364 4292 9463
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5920 9364 5948 9540
rect 6822 9528 6828 9540
rect 6880 9568 6886 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 6880 9540 7205 9568
rect 6880 9528 6886 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 8662 9500 8668 9512
rect 7515 9472 8668 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 9416 9509 9444 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 12342 9704 12348 9716
rect 11388 9676 12348 9704
rect 11388 9664 11394 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 17494 9704 17500 9716
rect 13832 9676 17500 9704
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9636 13507 9639
rect 13832 9636 13860 9676
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20622 9704 20628 9716
rect 20220 9676 20628 9704
rect 20220 9664 20226 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 25222 9704 25228 9716
rect 22704 9676 25228 9704
rect 22704 9664 22710 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 29914 9704 29920 9716
rect 29875 9676 29920 9704
rect 29914 9664 29920 9676
rect 29972 9664 29978 9716
rect 30006 9664 30012 9716
rect 30064 9704 30070 9716
rect 34514 9704 34520 9716
rect 30064 9676 34520 9704
rect 30064 9664 30070 9676
rect 34514 9664 34520 9676
rect 34572 9664 34578 9716
rect 13495 9608 13860 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 13906 9596 13912 9648
rect 13964 9596 13970 9648
rect 15838 9636 15844 9648
rect 14752 9608 15844 9636
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11112 9540 11713 9568
rect 11112 9528 11118 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12986 9568 12992 9580
rect 12575 9540 12992 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13170 9568 13176 9580
rect 13131 9540 13176 9568
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9469 9459 9503
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 9401 9463 9459 9469
rect 9508 9472 9689 9500
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 6914 9432 6920 9444
rect 6043 9404 6920 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 8941 9435 8999 9441
rect 8941 9432 8953 9435
rect 8904 9404 8953 9432
rect 8904 9392 8910 9404
rect 8941 9401 8953 9404
rect 8987 9432 8999 9435
rect 9508 9432 9536 9472
rect 9677 9469 9689 9472
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 14752 9500 14780 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 16209 9639 16267 9645
rect 16209 9605 16221 9639
rect 16255 9636 16267 9639
rect 19889 9639 19947 9645
rect 16255 9608 17618 9636
rect 16255 9605 16267 9608
rect 16209 9599 16267 9605
rect 19889 9605 19901 9639
rect 19935 9636 19947 9639
rect 19978 9636 19984 9648
rect 19935 9608 19984 9636
rect 19935 9605 19947 9608
rect 19889 9599 19947 9605
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 24121 9639 24179 9645
rect 24121 9636 24133 9639
rect 21114 9608 24133 9636
rect 24121 9605 24133 9608
rect 24167 9605 24179 9639
rect 24762 9636 24768 9648
rect 24723 9608 24768 9636
rect 24121 9599 24179 9605
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 27430 9636 27436 9648
rect 24912 9608 24957 9636
rect 27391 9608 27436 9636
rect 24912 9596 24918 9608
rect 27430 9596 27436 9608
rect 27488 9596 27494 9648
rect 27525 9639 27583 9645
rect 27525 9605 27537 9639
rect 27571 9636 27583 9639
rect 28350 9636 28356 9648
rect 27571 9608 28356 9636
rect 27571 9605 27583 9608
rect 27525 9599 27583 9605
rect 28350 9596 28356 9608
rect 28408 9596 28414 9648
rect 28810 9596 28816 9648
rect 28868 9636 28874 9648
rect 28868 9608 29868 9636
rect 28868 9596 28874 9608
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 15473 9571 15531 9577
rect 15473 9568 15485 9571
rect 15068 9540 15485 9568
rect 15068 9528 15074 9540
rect 15473 9537 15485 9540
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16298 9568 16304 9580
rect 16163 9540 16304 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9568 22523 9571
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22511 9540 23121 9568
rect 22511 9537 22523 9540
rect 22465 9531 22523 9537
rect 23109 9537 23121 9540
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 9824 9472 14780 9500
rect 15565 9503 15623 9509
rect 9824 9460 9830 9472
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 16666 9500 16672 9512
rect 15611 9472 16672 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9469 16911 9503
rect 17126 9500 17132 9512
rect 17087 9472 17132 9500
rect 16853 9463 16911 9469
rect 8987 9404 9536 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 16868 9432 16896 9463
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 17494 9460 17500 9512
rect 17552 9500 17558 9512
rect 17552 9472 19104 9500
rect 17552 9460 17558 9472
rect 16172 9404 16896 9432
rect 16172 9392 16178 9404
rect 4264 9336 5948 9364
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 9306 9364 9312 9376
rect 8076 9336 9312 9364
rect 8076 9324 8082 9336
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 12621 9367 12679 9373
rect 12621 9364 12633 9367
rect 11388 9336 12633 9364
rect 11388 9324 11394 9336
rect 12621 9333 12633 9336
rect 12667 9333 12679 9367
rect 12621 9327 12679 9333
rect 14921 9367 14979 9373
rect 14921 9333 14933 9367
rect 14967 9364 14979 9367
rect 17218 9364 17224 9376
rect 14967 9336 17224 9364
rect 14967 9333 14979 9336
rect 14921 9327 14979 9333
rect 17218 9324 17224 9336
rect 17276 9364 17282 9376
rect 17586 9364 17592 9376
rect 17276 9336 17592 9364
rect 17276 9324 17282 9336
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 18598 9364 18604 9376
rect 18559 9336 18604 9364
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 18966 9364 18972 9376
rect 18748 9336 18972 9364
rect 18748 9324 18754 9336
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 19076 9364 19104 9472
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19484 9472 19625 9500
rect 19484 9460 19490 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 21361 9503 21419 9509
rect 21361 9500 21373 9503
rect 19613 9463 19671 9469
rect 19720 9472 21373 9500
rect 19150 9392 19156 9444
rect 19208 9432 19214 9444
rect 19720 9432 19748 9472
rect 21361 9469 21373 9472
rect 21407 9500 21419 9503
rect 21634 9500 21640 9512
rect 21407 9472 21640 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 21634 9460 21640 9472
rect 21692 9460 21698 9512
rect 23124 9500 23152 9531
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 24029 9571 24087 9577
rect 24029 9568 24041 9571
rect 23440 9540 24041 9568
rect 23440 9528 23446 9540
rect 24029 9537 24041 9540
rect 24075 9568 24087 9571
rect 24210 9568 24216 9580
rect 24075 9540 24216 9568
rect 24075 9537 24087 9540
rect 24029 9531 24087 9537
rect 24210 9528 24216 9540
rect 24268 9528 24274 9580
rect 25406 9528 25412 9580
rect 25464 9568 25470 9580
rect 25866 9568 25872 9580
rect 25464 9540 25872 9568
rect 25464 9528 25470 9540
rect 25866 9528 25872 9540
rect 25924 9528 25930 9580
rect 28905 9571 28963 9577
rect 28905 9537 28917 9571
rect 28951 9568 28963 9571
rect 29638 9568 29644 9580
rect 28951 9540 29644 9568
rect 28951 9537 28963 9540
rect 28905 9531 28963 9537
rect 29638 9528 29644 9540
rect 29696 9528 29702 9580
rect 29840 9577 29868 9608
rect 29825 9571 29883 9577
rect 29825 9537 29837 9571
rect 29871 9568 29883 9571
rect 32398 9568 32404 9580
rect 29871 9540 32404 9568
rect 29871 9537 29883 9540
rect 29825 9531 29883 9537
rect 32398 9528 32404 9540
rect 32456 9528 32462 9580
rect 24762 9500 24768 9512
rect 23124 9472 24768 9500
rect 24762 9460 24768 9472
rect 24820 9460 24826 9512
rect 27982 9500 27988 9512
rect 27943 9472 27988 9500
rect 27982 9460 27988 9472
rect 28040 9460 28046 9512
rect 19208 9404 19748 9432
rect 19208 9392 19214 9404
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 23201 9435 23259 9441
rect 23201 9432 23213 9435
rect 20956 9404 23213 9432
rect 20956 9392 20962 9404
rect 23201 9401 23213 9404
rect 23247 9401 23259 9435
rect 24946 9432 24952 9444
rect 23201 9395 23259 9401
rect 23308 9404 24952 9432
rect 21358 9364 21364 9376
rect 19076 9336 21364 9364
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 22554 9364 22560 9376
rect 22515 9336 22560 9364
rect 22554 9324 22560 9336
rect 22612 9324 22618 9376
rect 23106 9324 23112 9376
rect 23164 9364 23170 9376
rect 23308 9364 23336 9404
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 25317 9435 25375 9441
rect 25317 9401 25329 9435
rect 25363 9432 25375 9435
rect 29270 9432 29276 9444
rect 25363 9404 29276 9432
rect 25363 9401 25375 9404
rect 25317 9395 25375 9401
rect 29270 9392 29276 9404
rect 29328 9392 29334 9444
rect 23164 9336 23336 9364
rect 23164 9324 23170 9336
rect 24486 9324 24492 9376
rect 24544 9364 24550 9376
rect 25961 9367 26019 9373
rect 25961 9364 25973 9367
rect 24544 9336 25973 9364
rect 24544 9324 24550 9336
rect 25961 9333 25973 9336
rect 26007 9333 26019 9367
rect 25961 9327 26019 9333
rect 28997 9367 29055 9373
rect 28997 9333 29009 9367
rect 29043 9364 29055 9367
rect 29914 9364 29920 9376
rect 29043 9336 29920 9364
rect 29043 9333 29055 9336
rect 28997 9327 29055 9333
rect 29914 9324 29920 9336
rect 29972 9324 29978 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2685 9163 2743 9169
rect 2685 9129 2697 9163
rect 2731 9160 2743 9163
rect 4614 9160 4620 9172
rect 2731 9132 4620 9160
rect 2731 9129 2743 9132
rect 2685 9123 2743 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 4982 9160 4988 9172
rect 4943 9132 4988 9160
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 9398 9160 9404 9172
rect 6840 9132 9404 9160
rect 3234 9052 3240 9104
rect 3292 9092 3298 9104
rect 6840 9092 6868 9132
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 11146 9160 11152 9172
rect 9508 9132 11152 9160
rect 3292 9064 6868 9092
rect 3292 9052 3298 9064
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 9508 9092 9536 9132
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 14182 9160 14188 9172
rect 11471 9132 14188 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14332 9132 14381 9160
rect 14332 9120 14338 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 15470 9160 15476 9172
rect 14369 9123 14427 9129
rect 14476 9132 15476 9160
rect 8076 9064 9536 9092
rect 8076 9052 8082 9064
rect 13446 9052 13452 9104
rect 13504 9092 13510 9104
rect 13633 9095 13691 9101
rect 13633 9092 13645 9095
rect 13504 9064 13645 9092
rect 13504 9052 13510 9064
rect 13633 9061 13645 9064
rect 13679 9092 13691 9095
rect 14476 9092 14504 9132
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 16574 9160 16580 9172
rect 15620 9132 16580 9160
rect 15620 9120 15626 9132
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 16850 9160 16856 9172
rect 16811 9132 16856 9160
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18509 9163 18567 9169
rect 18509 9160 18521 9163
rect 17920 9132 18521 9160
rect 17920 9120 17926 9132
rect 18509 9129 18521 9132
rect 18555 9129 18567 9163
rect 18509 9123 18567 9129
rect 18984 9132 21128 9160
rect 18984 9104 19012 9132
rect 13679 9064 14504 9092
rect 13679 9061 13691 9064
rect 13633 9055 13691 9061
rect 18414 9052 18420 9104
rect 18472 9092 18478 9104
rect 18966 9092 18972 9104
rect 18472 9064 18972 9092
rect 18472 9052 18478 9064
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 19702 9092 19708 9104
rect 19076 9064 19708 9092
rect 3142 8984 3148 9036
rect 3200 9024 3206 9036
rect 8386 9024 8392 9036
rect 3200 8996 8392 9024
rect 3200 8984 3206 8996
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 10410 9024 10416 9036
rect 9692 8996 10416 9024
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3936 8928 3985 8956
rect 3936 8916 3942 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4764 8928 4905 8956
rect 4764 8916 4770 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 6454 8956 6460 8968
rect 5767 8928 6460 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6730 8956 6736 8968
rect 6691 8928 6736 8956
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9692 8965 9720 8996
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 15105 9027 15163 9033
rect 12952 8996 14320 9024
rect 12952 8984 12958 8996
rect 14292 8965 14320 8996
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 16114 9024 16120 9036
rect 15151 8996 16120 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 19076 9024 19104 9064
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 21100 9092 21128 9132
rect 21174 9120 21180 9172
rect 21232 9160 21238 9172
rect 24670 9160 24676 9172
rect 21232 9132 24676 9160
rect 21232 9120 21238 9132
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 24762 9120 24768 9172
rect 24820 9160 24826 9172
rect 32122 9160 32128 9172
rect 24820 9132 32128 9160
rect 24820 9120 24826 9132
rect 32122 9120 32128 9132
rect 32180 9120 32186 9172
rect 21100 9064 22416 9092
rect 16448 8996 19104 9024
rect 16448 8984 16454 8996
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 19392 8996 19809 9024
rect 19392 8984 19398 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19797 8987 19855 8993
rect 20073 9027 20131 9033
rect 20073 8993 20085 9027
rect 20119 9024 20131 9027
rect 21818 9024 21824 9036
rect 20119 8996 21824 9024
rect 20119 8993 20131 8996
rect 20073 8987 20131 8993
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 22060 8996 22293 9024
rect 22060 8984 22066 8996
rect 22281 8993 22293 8996
rect 22327 8993 22339 9027
rect 22388 9024 22416 9064
rect 23750 9052 23756 9104
rect 23808 9092 23814 9104
rect 24029 9095 24087 9101
rect 24029 9092 24041 9095
rect 23808 9064 24041 9092
rect 23808 9052 23814 9064
rect 24029 9061 24041 9064
rect 24075 9092 24087 9095
rect 25774 9092 25780 9104
rect 24075 9064 25780 9092
rect 24075 9061 24087 9064
rect 24029 9055 24087 9061
rect 25774 9052 25780 9064
rect 25832 9052 25838 9104
rect 25866 9052 25872 9104
rect 25924 9092 25930 9104
rect 26142 9092 26148 9104
rect 25924 9064 26148 9092
rect 25924 9052 25930 9064
rect 26142 9052 26148 9064
rect 26200 9092 26206 9104
rect 26200 9064 26556 9092
rect 26200 9052 26206 9064
rect 22557 9027 22615 9033
rect 22557 9024 22569 9027
rect 22388 8996 22569 9024
rect 22281 8987 22339 8993
rect 22557 8993 22569 8996
rect 22603 9024 22615 9027
rect 26418 9024 26424 9036
rect 22603 8996 26424 9024
rect 22603 8993 22615 8996
rect 22557 8987 22615 8993
rect 26418 8984 26424 8996
rect 26476 8984 26482 9036
rect 26528 9033 26556 9064
rect 27982 9052 27988 9104
rect 28040 9092 28046 9104
rect 33042 9092 33048 9104
rect 28040 9064 33048 9092
rect 28040 9052 28046 9064
rect 33042 9052 33048 9064
rect 33100 9052 33106 9104
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 8993 26571 9027
rect 26513 8987 26571 8993
rect 9684 8959 9742 8965
rect 8628 8928 8892 8956
rect 8628 8916 8634 8928
rect 7009 8891 7067 8897
rect 7009 8857 7021 8891
rect 7055 8857 7067 8891
rect 8754 8888 8760 8900
rect 8234 8860 8760 8888
rect 7009 8851 7067 8857
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 2133 8823 2191 8829
rect 2133 8820 2145 8823
rect 2096 8792 2145 8820
rect 2096 8780 2102 8792
rect 2133 8789 2145 8792
rect 2179 8789 2191 8823
rect 2133 8783 2191 8789
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 3108 8792 4077 8820
rect 3108 8780 3114 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 4065 8783 4123 8789
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 5040 8792 5549 8820
rect 5040 8780 5046 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 7024 8820 7052 8851
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 8864 8888 8892 8928
rect 9684 8925 9696 8959
rect 9730 8925 9742 8959
rect 9684 8919 9742 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 18414 8956 18420 8968
rect 16724 8928 17816 8956
rect 18375 8928 18420 8956
rect 16724 8916 16730 8928
rect 9953 8891 10011 8897
rect 8864 8860 9904 8888
rect 7742 8820 7748 8832
rect 7024 8792 7748 8820
rect 5537 8783 5595 8789
rect 7742 8780 7748 8792
rect 7800 8820 7806 8832
rect 8018 8820 8024 8832
rect 7800 8792 8024 8820
rect 7800 8780 7806 8792
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 9674 8820 9680 8832
rect 8527 8792 9680 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9876 8820 9904 8860
rect 9953 8857 9965 8891
rect 9999 8888 10011 8891
rect 10042 8888 10048 8900
rect 9999 8860 10048 8888
rect 9999 8857 10011 8860
rect 9953 8851 10011 8857
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 12158 8888 12164 8900
rect 10244 8860 10442 8888
rect 12119 8860 12164 8888
rect 10244 8820 10272 8860
rect 12158 8848 12164 8860
rect 12216 8848 12222 8900
rect 12250 8848 12256 8900
rect 12308 8888 12314 8900
rect 15381 8891 15439 8897
rect 12308 8860 12650 8888
rect 12308 8848 12314 8860
rect 15381 8857 15393 8891
rect 15427 8888 15439 8891
rect 15470 8888 15476 8900
rect 15427 8860 15476 8888
rect 15427 8857 15439 8860
rect 15381 8851 15439 8857
rect 15470 8848 15476 8860
rect 15528 8848 15534 8900
rect 17678 8888 17684 8900
rect 16606 8860 17684 8888
rect 17678 8848 17684 8860
rect 17736 8848 17742 8900
rect 17788 8888 17816 8928
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 24486 8956 24492 8968
rect 21508 8928 22094 8956
rect 23690 8928 24492 8956
rect 21508 8916 21514 8928
rect 20162 8888 20168 8900
rect 17788 8860 20168 8888
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 21818 8888 21824 8900
rect 21298 8860 21404 8888
rect 21779 8860 21824 8888
rect 9876 8792 10272 8820
rect 13722 8780 13728 8832
rect 13780 8820 13786 8832
rect 21082 8820 21088 8832
rect 13780 8792 21088 8820
rect 13780 8780 13786 8792
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 21376 8820 21404 8860
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 22066 8888 22094 8928
rect 24486 8916 24492 8928
rect 24544 8916 24550 8968
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 24670 8956 24676 8968
rect 24627 8928 24676 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 24670 8916 24676 8928
rect 24728 8916 24734 8968
rect 25225 8959 25283 8965
rect 25225 8925 25237 8959
rect 25271 8956 25283 8959
rect 25406 8956 25412 8968
rect 25271 8928 25412 8956
rect 25271 8925 25283 8928
rect 25225 8919 25283 8925
rect 25406 8916 25412 8928
rect 25464 8916 25470 8968
rect 34514 8916 34520 8968
rect 34572 8956 34578 8968
rect 34885 8959 34943 8965
rect 34885 8956 34897 8959
rect 34572 8928 34897 8956
rect 34572 8916 34578 8928
rect 34885 8925 34897 8928
rect 34931 8925 34943 8959
rect 34885 8919 34943 8925
rect 36078 8916 36084 8968
rect 36136 8956 36142 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 36136 8928 38025 8956
rect 36136 8916 36142 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 22462 8888 22468 8900
rect 22066 8860 22468 8888
rect 22462 8848 22468 8860
rect 22520 8848 22526 8900
rect 25317 8891 25375 8897
rect 25317 8888 25329 8891
rect 23860 8860 25329 8888
rect 23860 8820 23888 8860
rect 25317 8857 25329 8860
rect 25363 8857 25375 8891
rect 26142 8888 26148 8900
rect 26103 8860 26148 8888
rect 25317 8851 25375 8857
rect 26142 8848 26148 8860
rect 26200 8848 26206 8900
rect 26234 8848 26240 8900
rect 26292 8888 26298 8900
rect 26292 8860 26337 8888
rect 26292 8848 26298 8860
rect 21376 8792 23888 8820
rect 24673 8823 24731 8829
rect 24673 8789 24685 8823
rect 24719 8820 24731 8823
rect 25222 8820 25228 8832
rect 24719 8792 25228 8820
rect 24719 8789 24731 8792
rect 24673 8783 24731 8789
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 34977 8823 35035 8829
rect 34977 8789 34989 8823
rect 35023 8820 35035 8823
rect 36262 8820 36268 8832
rect 35023 8792 36268 8820
rect 35023 8789 35035 8792
rect 34977 8783 35035 8789
rect 36262 8780 36268 8792
rect 36320 8780 36326 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 5994 8616 6000 8628
rect 3660 8588 4752 8616
rect 5955 8588 6000 8616
rect 3660 8576 3666 8588
rect 2133 8551 2191 8557
rect 2133 8517 2145 8551
rect 2179 8548 2191 8551
rect 3142 8548 3148 8560
rect 2179 8520 3148 8548
rect 2179 8517 2191 8520
rect 2133 8511 2191 8517
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 4614 8548 4620 8560
rect 3436 8520 4620 8548
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2682 8480 2688 8492
rect 2363 8452 2688 8480
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 3436 8489 3464 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 4724 8548 4752 8588
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 9674 8616 9680 8628
rect 7208 8588 9680 8616
rect 4724 8520 5014 8548
rect 7208 8489 7236 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 14366 8616 14372 8628
rect 10560 8588 14372 8616
rect 10560 8576 10566 8588
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 16666 8616 16672 8628
rect 15068 8588 16672 8616
rect 15068 8576 15074 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 19426 8616 19432 8628
rect 17236 8588 19432 8616
rect 11606 8548 11612 8560
rect 8694 8520 11612 8548
rect 11606 8508 11612 8520
rect 11664 8508 11670 8560
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 11940 8520 12449 8548
rect 11940 8508 11946 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 13446 8548 13452 8560
rect 13407 8520 13452 8548
rect 12437 8511 12495 8517
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 13596 8520 13938 8548
rect 13596 8508 13602 8520
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 7193 8483 7251 8489
rect 7193 8449 7205 8483
rect 7239 8449 7251 8483
rect 9398 8480 9404 8492
rect 9359 8452 9404 8480
rect 7193 8443 7251 8449
rect 2976 8412 3004 8443
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 10284 8452 11161 8480
rect 10284 8440 10290 8452
rect 11149 8449 11161 8452
rect 11195 8480 11207 8483
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11195 8452 11713 8480
rect 11195 8449 11207 8452
rect 11149 8443 11207 8449
rect 11701 8449 11713 8452
rect 11747 8480 11759 8483
rect 12342 8480 12348 8492
rect 11747 8452 12348 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 13170 8480 13176 8492
rect 13131 8452 13176 8480
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 17236 8489 17264 8588
rect 19426 8576 19432 8588
rect 19484 8616 19490 8628
rect 19518 8616 19524 8628
rect 19484 8588 19524 8616
rect 19484 8576 19490 8588
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 23198 8616 23204 8628
rect 20180 8588 23204 8616
rect 20180 8548 20208 8588
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 28350 8616 28356 8628
rect 28311 8588 28356 8616
rect 28350 8576 28356 8588
rect 28408 8576 28414 8628
rect 28534 8576 28540 8628
rect 28592 8616 28598 8628
rect 29641 8619 29699 8625
rect 29641 8616 29653 8619
rect 28592 8588 29653 8616
rect 28592 8576 28598 8588
rect 29641 8585 29653 8588
rect 29687 8585 29699 8619
rect 36078 8616 36084 8628
rect 36039 8588 36084 8616
rect 29641 8579 29699 8585
rect 36078 8576 36084 8588
rect 36136 8576 36142 8628
rect 21634 8548 21640 8560
rect 18722 8520 20208 8548
rect 21022 8520 21640 8548
rect 21634 8508 21640 8520
rect 21692 8508 21698 8560
rect 23658 8548 23664 8560
rect 23619 8520 23664 8548
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 25222 8548 25228 8560
rect 25183 8520 25228 8548
rect 25222 8508 25228 8520
rect 25280 8508 25286 8560
rect 25314 8508 25320 8560
rect 25372 8548 25378 8560
rect 26145 8551 26203 8557
rect 26145 8548 26157 8551
rect 25372 8520 26157 8548
rect 25372 8508 25378 8520
rect 26145 8517 26157 8520
rect 26191 8517 26203 8551
rect 26145 8511 26203 8517
rect 17221 8483 17279 8489
rect 17221 8480 17233 8483
rect 16172 8452 17233 8480
rect 16172 8440 16178 8452
rect 17221 8449 17233 8452
rect 17267 8449 17279 8483
rect 19518 8480 19524 8492
rect 19479 8452 19524 8480
rect 17221 8443 17279 8449
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 23106 8480 23112 8492
rect 21284 8452 23112 8480
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 2976 8384 3525 8412
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3513 8375 3571 8381
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 6822 8412 6828 8424
rect 4571 8384 6828 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 2777 8347 2835 8353
rect 2777 8344 2789 8347
rect 2372 8316 2789 8344
rect 2372 8304 2378 8316
rect 2777 8313 2789 8316
rect 2823 8313 2835 8347
rect 2777 8307 2835 8313
rect 4264 8276 4292 8375
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8412 7527 8415
rect 13538 8412 13544 8424
rect 7515 8384 13544 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 17497 8415 17555 8421
rect 17497 8412 17509 8415
rect 17000 8384 17509 8412
rect 17000 8372 17006 8384
rect 17497 8381 17509 8384
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 17586 8372 17592 8424
rect 17644 8412 17650 8424
rect 17644 8384 18552 8412
rect 17644 8372 17650 8384
rect 8570 8304 8576 8356
rect 8628 8344 8634 8356
rect 12158 8344 12164 8356
rect 8628 8316 12164 8344
rect 8628 8304 8634 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 4614 8276 4620 8288
rect 4264 8248 4620 8276
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 8941 8279 8999 8285
rect 8941 8276 8953 8279
rect 8812 8248 8953 8276
rect 8812 8236 8818 8248
rect 8941 8245 8953 8248
rect 8987 8276 8999 8279
rect 9122 8276 9128 8288
rect 8987 8248 9128 8276
rect 8987 8245 8999 8248
rect 8941 8239 8999 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 14918 8276 14924 8288
rect 11296 8248 14924 8276
rect 11296 8236 11302 8248
rect 14918 8236 14924 8248
rect 14976 8236 14982 8288
rect 18524 8276 18552 8384
rect 18616 8384 21036 8412
rect 18616 8356 18644 8384
rect 18598 8304 18604 8356
rect 18656 8304 18662 8356
rect 21008 8344 21036 8384
rect 21082 8372 21088 8424
rect 21140 8412 21146 8424
rect 21284 8421 21312 8452
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 26050 8440 26056 8492
rect 26108 8480 26114 8492
rect 28261 8483 28319 8489
rect 28261 8480 28273 8483
rect 26108 8452 28273 8480
rect 26108 8440 26114 8452
rect 28261 8449 28273 8452
rect 28307 8449 28319 8483
rect 28261 8443 28319 8449
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 28905 8483 28963 8489
rect 28905 8480 28917 8483
rect 28408 8452 28917 8480
rect 28408 8440 28414 8452
rect 28905 8449 28917 8452
rect 28951 8480 28963 8483
rect 29086 8480 29092 8492
rect 28951 8452 29092 8480
rect 28951 8449 28963 8452
rect 28905 8443 28963 8449
rect 29086 8440 29092 8452
rect 29144 8440 29150 8492
rect 29549 8483 29607 8489
rect 29549 8449 29561 8483
rect 29595 8480 29607 8483
rect 35802 8480 35808 8492
rect 29595 8452 35808 8480
rect 29595 8449 29607 8452
rect 29549 8443 29607 8449
rect 35802 8440 35808 8452
rect 35860 8440 35866 8492
rect 36262 8480 36268 8492
rect 36223 8452 36268 8480
rect 36262 8440 36268 8452
rect 36320 8440 36326 8492
rect 21269 8415 21327 8421
rect 21269 8412 21281 8415
rect 21140 8384 21281 8412
rect 21140 8372 21146 8384
rect 21269 8381 21281 8384
rect 21315 8381 21327 8415
rect 21269 8375 21327 8381
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 23014 8412 23020 8424
rect 21416 8384 23020 8412
rect 21416 8372 21422 8384
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 23569 8415 23627 8421
rect 23569 8412 23581 8415
rect 23492 8384 23581 8412
rect 23492 8356 23520 8384
rect 23569 8381 23581 8384
rect 23615 8381 23627 8415
rect 24026 8412 24032 8424
rect 23987 8384 24032 8412
rect 23569 8375 23627 8381
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 25133 8415 25191 8421
rect 25133 8412 25145 8415
rect 24912 8384 25145 8412
rect 24912 8372 24918 8384
rect 25133 8381 25145 8384
rect 25179 8412 25191 8415
rect 25958 8412 25964 8424
rect 25179 8384 25964 8412
rect 25179 8381 25191 8384
rect 25133 8375 25191 8381
rect 25958 8372 25964 8384
rect 26016 8372 26022 8424
rect 26602 8372 26608 8424
rect 26660 8412 26666 8424
rect 27157 8415 27215 8421
rect 27157 8412 27169 8415
rect 26660 8384 27169 8412
rect 26660 8372 26666 8384
rect 27157 8381 27169 8384
rect 27203 8381 27215 8415
rect 27157 8375 27215 8381
rect 27341 8415 27399 8421
rect 27341 8381 27353 8415
rect 27387 8412 27399 8415
rect 28997 8415 29055 8421
rect 28997 8412 29009 8415
rect 27387 8384 29009 8412
rect 27387 8381 27399 8384
rect 27341 8375 27399 8381
rect 28997 8381 29009 8384
rect 29043 8381 29055 8415
rect 28997 8375 29055 8381
rect 18708 8316 19656 8344
rect 21008 8316 23152 8344
rect 18708 8276 18736 8316
rect 18966 8276 18972 8288
rect 18524 8248 18736 8276
rect 18927 8248 18972 8276
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19628 8276 19656 8316
rect 19778 8279 19836 8285
rect 19778 8276 19790 8279
rect 19628 8248 19790 8276
rect 19778 8245 19790 8248
rect 19824 8245 19836 8279
rect 23124 8276 23152 8316
rect 23474 8304 23480 8356
rect 23532 8304 23538 8356
rect 27801 8347 27859 8353
rect 27801 8313 27813 8347
rect 27847 8344 27859 8347
rect 28442 8344 28448 8356
rect 27847 8316 28448 8344
rect 27847 8313 27859 8316
rect 27801 8307 27859 8313
rect 28442 8304 28448 8316
rect 28500 8304 28506 8356
rect 28350 8276 28356 8288
rect 23124 8248 28356 8276
rect 19778 8239 19836 8245
rect 28350 8236 28356 8248
rect 28408 8236 28414 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 2501 8075 2559 8081
rect 2501 8072 2513 8075
rect 2464 8044 2513 8072
rect 2464 8032 2470 8044
rect 2501 8041 2513 8044
rect 2547 8041 2559 8075
rect 2501 8035 2559 8041
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 4028 8044 4077 8072
rect 4028 8032 4034 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4880 8075 4938 8081
rect 4880 8041 4892 8075
rect 4926 8072 4938 8075
rect 5994 8072 6000 8084
rect 4926 8044 6000 8072
rect 4926 8041 4938 8044
rect 4880 8035 4938 8041
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6362 8072 6368 8084
rect 6323 8044 6368 8072
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 10134 8072 10140 8084
rect 6472 8044 10140 8072
rect 6086 7964 6092 8016
rect 6144 8004 6150 8016
rect 6472 8004 6500 8044
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 15102 8072 15108 8084
rect 10244 8044 15108 8072
rect 6144 7976 6500 8004
rect 6144 7964 6150 7976
rect 4614 7936 4620 7948
rect 4575 7908 4620 7936
rect 4614 7896 4620 7908
rect 4672 7936 4678 7948
rect 5626 7936 5632 7948
rect 4672 7908 5632 7936
rect 4672 7896 4678 7908
rect 5626 7896 5632 7908
rect 5684 7936 5690 7948
rect 6730 7936 6736 7948
rect 5684 7908 6736 7936
rect 5684 7896 5690 7908
rect 6730 7896 6736 7908
rect 6788 7936 6794 7948
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 6788 7908 6837 7936
rect 6788 7896 6794 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 10244 7936 10272 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 17126 8072 17132 8084
rect 15212 8044 17132 8072
rect 12713 8007 12771 8013
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 12802 8004 12808 8016
rect 12759 7976 12808 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 12802 7964 12808 7976
rect 12860 8004 12866 8016
rect 15212 8004 15240 8044
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17678 8032 17684 8084
rect 17736 8072 17742 8084
rect 17736 8044 21036 8072
rect 17736 8032 17742 8044
rect 12860 7976 15240 8004
rect 17957 8007 18015 8013
rect 12860 7964 12866 7976
rect 17957 7973 17969 8007
rect 18003 8004 18015 8007
rect 18138 8004 18144 8016
rect 18003 7976 18144 8004
rect 18003 7973 18015 7976
rect 17957 7967 18015 7973
rect 18138 7964 18144 7976
rect 18196 8004 18202 8016
rect 18690 8004 18696 8016
rect 18196 7976 18696 8004
rect 18196 7964 18202 7976
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 21008 8004 21036 8044
rect 21174 8032 21180 8084
rect 21232 8072 21238 8084
rect 24394 8072 24400 8084
rect 21232 8044 24400 8072
rect 21232 8032 21238 8044
rect 24394 8032 24400 8044
rect 24452 8032 24458 8084
rect 26326 8032 26332 8084
rect 26384 8072 26390 8084
rect 27614 8072 27620 8084
rect 26384 8044 27620 8072
rect 26384 8032 26390 8044
rect 27614 8032 27620 8044
rect 27672 8032 27678 8084
rect 21008 7976 21588 8004
rect 7147 7908 10272 7936
rect 10965 7939 11023 7945
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 13170 7936 13176 7948
rect 11011 7908 13176 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 16172 7908 16221 7936
rect 16172 7896 16178 7908
rect 16209 7905 16221 7908
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 18966 7936 18972 7948
rect 16531 7908 18972 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 19518 7936 19524 7948
rect 19479 7908 19524 7936
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 20806 7936 20812 7948
rect 19843 7908 20812 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 20806 7896 20812 7908
rect 20864 7896 20870 7948
rect 21560 7945 21588 7976
rect 24762 7964 24768 8016
rect 24820 8004 24826 8016
rect 24820 7976 35894 8004
rect 24820 7964 24826 7976
rect 21545 7939 21603 7945
rect 21545 7905 21557 7939
rect 21591 7936 21603 7939
rect 22738 7936 22744 7948
rect 21591 7908 22744 7936
rect 21591 7905 21603 7908
rect 21545 7899 21603 7905
rect 22738 7896 22744 7908
rect 22796 7896 22802 7948
rect 24210 7896 24216 7948
rect 24268 7936 24274 7948
rect 25774 7936 25780 7948
rect 24268 7908 25780 7936
rect 24268 7896 24274 7908
rect 25774 7896 25780 7908
rect 25832 7896 25838 7948
rect 26142 7896 26148 7948
rect 26200 7936 26206 7948
rect 27525 7939 27583 7945
rect 27525 7936 27537 7939
rect 26200 7908 27537 7936
rect 26200 7896 26206 7908
rect 27525 7905 27537 7908
rect 27571 7905 27583 7939
rect 28534 7936 28540 7948
rect 28495 7908 28540 7936
rect 27525 7899 27583 7905
rect 28534 7896 28540 7908
rect 28592 7896 28598 7948
rect 29181 7939 29239 7945
rect 29181 7905 29193 7939
rect 29227 7936 29239 7939
rect 29270 7936 29276 7948
rect 29227 7908 29276 7936
rect 29227 7905 29239 7908
rect 29181 7899 29239 7905
rect 29270 7896 29276 7908
rect 29328 7896 29334 7948
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 2774 7868 2780 7880
rect 2731 7840 2780 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 3326 7868 3332 7880
rect 3287 7840 3332 7868
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12952 7840 13277 7868
rect 12952 7828 12958 7840
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 18506 7868 18512 7880
rect 18467 7840 18512 7868
rect 13265 7831 13323 7837
rect 18506 7828 18512 7840
rect 18564 7868 18570 7880
rect 18564 7840 19334 7868
rect 18564 7828 18570 7840
rect 5902 7760 5908 7812
rect 5960 7760 5966 7812
rect 6178 7760 6184 7812
rect 6236 7800 6242 7812
rect 11238 7800 11244 7812
rect 6236 7772 7590 7800
rect 11199 7772 11244 7800
rect 6236 7760 6242 7772
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 11882 7760 11888 7812
rect 11940 7760 11946 7812
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13357 7803 13415 7809
rect 13357 7800 13369 7803
rect 12584 7772 13369 7800
rect 12584 7760 12590 7772
rect 13357 7769 13369 7772
rect 13403 7769 13415 7803
rect 14734 7800 14740 7812
rect 14695 7772 14740 7800
rect 13357 7763 13415 7769
rect 14734 7760 14740 7772
rect 14792 7760 14798 7812
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 15473 7803 15531 7809
rect 15473 7800 15485 7803
rect 15160 7772 15485 7800
rect 15160 7760 15166 7772
rect 15473 7769 15485 7772
rect 15519 7769 15531 7803
rect 18782 7800 18788 7812
rect 17710 7772 18788 7800
rect 15473 7763 15531 7769
rect 18782 7760 18788 7772
rect 18840 7760 18846 7812
rect 19306 7800 19334 7840
rect 22830 7828 22836 7880
rect 22888 7868 22894 7880
rect 23385 7871 23443 7877
rect 23385 7868 23397 7871
rect 22888 7840 23397 7868
rect 22888 7828 22894 7840
rect 23385 7837 23397 7840
rect 23431 7837 23443 7871
rect 35866 7868 35894 7976
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 35866 7840 38025 7868
rect 23385 7831 23443 7837
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 19886 7800 19892 7812
rect 19306 7772 19892 7800
rect 19886 7760 19892 7772
rect 19944 7760 19950 7812
rect 21082 7800 21088 7812
rect 21022 7772 21088 7800
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 24268 7772 24685 7800
rect 24268 7760 24274 7772
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 24765 7803 24823 7809
rect 24765 7769 24777 7803
rect 24811 7800 24823 7803
rect 24946 7800 24952 7812
rect 24811 7772 24952 7800
rect 24811 7769 24823 7772
rect 24765 7763 24823 7769
rect 24946 7760 24952 7772
rect 25004 7760 25010 7812
rect 25685 7803 25743 7809
rect 25685 7769 25697 7803
rect 25731 7800 25743 7803
rect 26142 7800 26148 7812
rect 25731 7772 26148 7800
rect 25731 7769 25743 7772
rect 25685 7763 25743 7769
rect 26142 7760 26148 7772
rect 26200 7760 26206 7812
rect 26421 7803 26479 7809
rect 26421 7800 26433 7803
rect 26344 7772 26433 7800
rect 26344 7744 26372 7772
rect 26421 7769 26433 7772
rect 26467 7769 26479 7803
rect 26421 7763 26479 7769
rect 26513 7803 26571 7809
rect 26513 7769 26525 7803
rect 26559 7769 26571 7803
rect 26513 7763 26571 7769
rect 27065 7803 27123 7809
rect 27065 7769 27077 7803
rect 27111 7800 27123 7803
rect 27614 7800 27620 7812
rect 27111 7772 27620 7800
rect 27111 7769 27123 7772
rect 27065 7763 27123 7769
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1728 7704 1869 7732
rect 1728 7692 1734 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 3142 7732 3148 7744
rect 3055 7704 3148 7732
rect 1857 7695 1915 7701
rect 3142 7692 3148 7704
rect 3200 7732 3206 7744
rect 3878 7732 3884 7744
rect 3200 7704 3884 7732
rect 3200 7692 3206 7704
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 8573 7735 8631 7741
rect 8573 7732 8585 7735
rect 7064 7704 8585 7732
rect 7064 7692 7070 7704
rect 8573 7701 8585 7704
rect 8619 7701 8631 7735
rect 8573 7695 8631 7701
rect 9306 7692 9312 7744
rect 9364 7732 9370 7744
rect 12066 7732 12072 7744
rect 9364 7704 12072 7732
rect 9364 7692 9370 7704
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18601 7735 18659 7741
rect 18601 7732 18613 7735
rect 18104 7704 18613 7732
rect 18104 7692 18110 7704
rect 18601 7701 18613 7704
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 21174 7732 21180 7744
rect 19024 7704 21180 7732
rect 19024 7692 19030 7704
rect 21174 7692 21180 7704
rect 21232 7692 21238 7744
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 22796 7704 23489 7732
rect 22796 7692 22802 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 26326 7692 26332 7744
rect 26384 7692 26390 7744
rect 26528 7732 26556 7763
rect 27614 7760 27620 7772
rect 27672 7760 27678 7812
rect 28629 7803 28687 7809
rect 28629 7769 28641 7803
rect 28675 7769 28687 7803
rect 28629 7763 28687 7769
rect 27890 7732 27896 7744
rect 26528 7704 27896 7732
rect 27890 7692 27896 7704
rect 27948 7692 27954 7744
rect 28644 7732 28672 7763
rect 31570 7732 31576 7744
rect 28644 7704 31576 7732
rect 31570 7692 31576 7704
rect 31628 7692 31634 7744
rect 38194 7732 38200 7744
rect 38155 7704 38200 7732
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2866 7528 2872 7540
rect 2827 7500 2872 7528
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 4525 7531 4583 7537
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 5350 7528 5356 7540
rect 4571 7500 5356 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5552 7500 9674 7528
rect 5552 7404 5580 7500
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 5684 7432 5825 7460
rect 5684 7420 5690 7432
rect 5813 7429 5825 7432
rect 5859 7429 5871 7463
rect 6638 7460 6644 7472
rect 6599 7432 6644 7460
rect 5813 7423 5871 7429
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 8021 7463 8079 7469
rect 8021 7460 8033 7463
rect 6972 7432 8033 7460
rect 6972 7420 6978 7432
rect 8021 7429 8033 7432
rect 8067 7429 8079 7463
rect 8021 7423 8079 7429
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 9646 7460 9674 7500
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 10502 7528 10508 7540
rect 9824 7500 10508 7528
rect 9824 7488 9830 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 15010 7528 15016 7540
rect 10796 7500 15016 7528
rect 10226 7460 10232 7472
rect 8352 7432 8510 7460
rect 9646 7432 10232 7460
rect 8352 7420 8358 7432
rect 10226 7420 10232 7432
rect 10284 7420 10290 7472
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 3053 7395 3111 7401
rect 3053 7392 3065 7395
rect 2004 7364 3065 7392
rect 2004 7352 2010 7364
rect 3053 7361 3065 7364
rect 3099 7361 3111 7395
rect 3786 7392 3792 7404
rect 3747 7364 3792 7392
rect 3053 7355 3111 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3936 7364 4445 7392
rect 3936 7352 3942 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5534 7392 5540 7404
rect 5123 7364 5540 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 6546 7392 6552 7404
rect 6507 7364 6552 7392
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 10134 7392 10140 7404
rect 9600 7364 10140 7392
rect 1578 7324 1584 7336
rect 1539 7296 1584 7324
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 2222 7284 2228 7336
rect 2280 7324 2286 7336
rect 6178 7324 6184 7336
rect 2280 7296 6184 7324
rect 2280 7284 2286 7296
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7064 7296 7757 7324
rect 7064 7284 7070 7296
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 9600 7324 9628 7364
rect 10134 7352 10140 7364
rect 10192 7392 10198 7404
rect 10796 7392 10824 7500
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 20438 7528 20444 7540
rect 17512 7500 20444 7528
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 11882 7460 11888 7472
rect 10928 7432 11888 7460
rect 10928 7420 10934 7432
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 13262 7460 13268 7472
rect 13223 7432 13268 7460
rect 13262 7420 13268 7432
rect 13320 7420 13326 7472
rect 17512 7460 17540 7500
rect 20438 7488 20444 7500
rect 20496 7488 20502 7540
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 21266 7488 21272 7540
rect 21324 7528 21330 7540
rect 21324 7500 24348 7528
rect 21324 7488 21330 7500
rect 19794 7460 19800 7472
rect 14490 7432 17540 7460
rect 18354 7432 19800 7460
rect 19794 7420 19800 7432
rect 19852 7420 19858 7472
rect 20990 7460 20996 7472
rect 20930 7432 20996 7460
rect 20990 7420 20996 7432
rect 21048 7420 21054 7472
rect 23201 7463 23259 7469
rect 23201 7429 23213 7463
rect 23247 7460 23259 7463
rect 24026 7460 24032 7472
rect 23247 7432 24032 7460
rect 23247 7429 23259 7432
rect 23201 7423 23259 7429
rect 24026 7420 24032 7432
rect 24084 7420 24090 7472
rect 24210 7460 24216 7472
rect 24171 7432 24216 7460
rect 24210 7420 24216 7432
rect 24268 7420 24274 7472
rect 24320 7460 24348 7500
rect 24946 7488 24952 7540
rect 25004 7528 25010 7540
rect 25004 7500 25049 7528
rect 25004 7488 25010 7500
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 27249 7531 27307 7537
rect 27249 7528 27261 7531
rect 26292 7500 27261 7528
rect 26292 7488 26298 7500
rect 27249 7497 27261 7500
rect 27295 7497 27307 7531
rect 27249 7491 27307 7497
rect 26786 7460 26792 7472
rect 24320 7432 26792 7460
rect 10192 7364 10824 7392
rect 10192 7352 10198 7364
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11204 7364 11989 7392
rect 11204 7352 11210 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 11977 7355 12035 7361
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 25516 7401 25544 7432
rect 26786 7420 26792 7432
rect 26844 7420 26850 7472
rect 24857 7395 24915 7401
rect 24857 7392 24869 7395
rect 23808 7364 24869 7392
rect 23808 7352 23814 7364
rect 24857 7361 24869 7364
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 25501 7395 25559 7401
rect 25501 7361 25513 7395
rect 25547 7361 25559 7395
rect 25501 7355 25559 7361
rect 26145 7395 26203 7401
rect 26145 7361 26157 7395
rect 26191 7361 26203 7395
rect 27154 7392 27160 7404
rect 27115 7364 27160 7392
rect 26145 7355 26203 7361
rect 9766 7324 9772 7336
rect 7745 7287 7803 7293
rect 7852 7296 9628 7324
rect 9727 7296 9772 7324
rect 2130 7216 2136 7268
rect 2188 7256 2194 7268
rect 7852 7256 7880 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10042 7284 10048 7336
rect 10100 7324 10106 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10100 7296 10977 7324
rect 10100 7284 10106 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7293 13047 7327
rect 16850 7324 16856 7336
rect 16811 7296 16856 7324
rect 12989 7287 13047 7293
rect 2188 7228 7880 7256
rect 2188 7216 2194 7228
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 11716 7256 11744 7287
rect 9916 7228 11744 7256
rect 9916 7216 9922 7228
rect 3881 7191 3939 7197
rect 3881 7157 3893 7191
rect 3927 7188 3939 7191
rect 6086 7188 6092 7200
rect 3927 7160 6092 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 6086 7148 6092 7160
rect 6144 7148 6150 7200
rect 7098 7148 7104 7200
rect 7156 7188 7162 7200
rect 11422 7188 11428 7200
rect 7156 7160 11428 7188
rect 7156 7148 7162 7160
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 13004 7188 13032 7287
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 18598 7324 18604 7336
rect 17175 7296 18604 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 19392 7296 19441 7324
rect 19392 7284 19398 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 22002 7324 22008 7336
rect 19852 7296 22008 7324
rect 19852 7284 19858 7296
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 23109 7327 23167 7333
rect 23109 7293 23121 7327
rect 23155 7324 23167 7327
rect 23474 7324 23480 7336
rect 23155 7296 23480 7324
rect 23155 7293 23167 7296
rect 23109 7287 23167 7293
rect 23474 7284 23480 7296
rect 23532 7284 23538 7336
rect 24026 7284 24032 7336
rect 24084 7324 24090 7336
rect 25593 7327 25651 7333
rect 25593 7324 25605 7327
rect 24084 7296 25605 7324
rect 24084 7284 24090 7296
rect 25593 7293 25605 7296
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 26160 7268 26188 7355
rect 27154 7352 27160 7364
rect 27212 7352 27218 7404
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 27246 7324 27252 7336
rect 26292 7296 27252 7324
rect 26292 7284 26298 7296
rect 27246 7284 27252 7296
rect 27304 7324 27310 7336
rect 31662 7324 31668 7336
rect 27304 7296 31668 7324
rect 27304 7284 27310 7296
rect 31662 7284 31668 7296
rect 31720 7284 31726 7336
rect 21910 7256 21916 7268
rect 21192 7228 21916 7256
rect 15102 7188 15108 7200
rect 13004 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 18601 7191 18659 7197
rect 18601 7188 18613 7191
rect 16816 7160 18613 7188
rect 16816 7148 16822 7160
rect 18601 7157 18613 7160
rect 18647 7188 18659 7191
rect 18782 7188 18788 7200
rect 18647 7160 18788 7188
rect 18647 7157 18659 7160
rect 18601 7151 18659 7157
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 19692 7191 19750 7197
rect 19692 7157 19704 7191
rect 19738 7188 19750 7191
rect 20714 7188 20720 7200
rect 19738 7160 20720 7188
rect 19738 7157 19750 7160
rect 19692 7151 19750 7157
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 20898 7148 20904 7200
rect 20956 7188 20962 7200
rect 21192 7188 21220 7228
rect 21910 7216 21916 7228
rect 21968 7216 21974 7268
rect 23661 7259 23719 7265
rect 23661 7225 23673 7259
rect 23707 7256 23719 7259
rect 23934 7256 23940 7268
rect 23707 7228 23940 7256
rect 23707 7225 23719 7228
rect 23661 7219 23719 7225
rect 23934 7216 23940 7228
rect 23992 7256 23998 7268
rect 24118 7256 24124 7268
rect 23992 7228 24124 7256
rect 23992 7216 23998 7228
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 25038 7216 25044 7268
rect 25096 7256 25102 7268
rect 26142 7256 26148 7268
rect 25096 7228 26148 7256
rect 25096 7216 25102 7228
rect 26142 7216 26148 7228
rect 26200 7216 26206 7268
rect 20956 7160 21220 7188
rect 20956 7148 20962 7160
rect 22094 7148 22100 7200
rect 22152 7188 22158 7200
rect 26237 7191 26295 7197
rect 26237 7188 26249 7191
rect 22152 7160 26249 7188
rect 22152 7148 22158 7160
rect 26237 7157 26249 7160
rect 26283 7157 26295 7191
rect 26237 7151 26295 7157
rect 34514 7148 34520 7200
rect 34572 7188 34578 7200
rect 38105 7191 38163 7197
rect 38105 7188 38117 7191
rect 34572 7160 38117 7188
rect 34572 7148 34578 7160
rect 38105 7157 38117 7160
rect 38151 7157 38163 7191
rect 38105 7151 38163 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 4880 6987 4938 6993
rect 4880 6953 4892 6987
rect 4926 6984 4938 6987
rect 9306 6984 9312 6996
rect 4926 6956 9312 6984
rect 4926 6953 4938 6956
rect 4880 6947 4938 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 15368 6987 15426 6993
rect 15368 6953 15380 6987
rect 15414 6984 15426 6987
rect 18690 6984 18696 6996
rect 15414 6956 18696 6984
rect 15414 6953 15426 6956
rect 15368 6947 15426 6953
rect 18690 6944 18696 6956
rect 18748 6944 18754 6996
rect 19968 6987 20026 6993
rect 19968 6953 19980 6987
rect 20014 6984 20026 6987
rect 20346 6984 20352 6996
rect 20014 6956 20352 6984
rect 20014 6953 20026 6956
rect 19968 6947 20026 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 20438 6944 20444 6996
rect 20496 6984 20502 6996
rect 27246 6984 27252 6996
rect 20496 6956 27252 6984
rect 20496 6944 20502 6956
rect 27246 6944 27252 6956
rect 27304 6944 27310 6996
rect 28997 6987 29055 6993
rect 28997 6953 29009 6987
rect 29043 6984 29055 6987
rect 29043 6956 29868 6984
rect 29043 6953 29055 6956
rect 28997 6947 29055 6953
rect 2225 6919 2283 6925
rect 2225 6885 2237 6919
rect 2271 6914 2283 6919
rect 16853 6919 16911 6925
rect 2271 6886 2305 6914
rect 2271 6885 2283 6886
rect 2225 6879 2283 6885
rect 16853 6885 16865 6919
rect 16899 6916 16911 6919
rect 16899 6888 18092 6916
rect 16899 6885 16911 6888
rect 16853 6879 16911 6885
rect 2240 6848 2268 6879
rect 3970 6848 3976 6860
rect 2240 6820 3976 6848
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 4304 6820 4629 6848
rect 4304 6808 4310 6820
rect 4617 6817 4629 6820
rect 4663 6848 4675 6851
rect 4663 6820 6224 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6780 1823 6783
rect 2222 6780 2228 6792
rect 1811 6752 2228 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2409 6783 2467 6789
rect 2409 6749 2421 6783
rect 2455 6749 2467 6783
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 2409 6743 2467 6749
rect 2424 6712 2452 6743
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 3234 6712 3240 6724
rect 2424 6684 3240 6712
rect 3234 6672 3240 6684
rect 3292 6672 3298 6724
rect 4172 6712 4200 6743
rect 4614 6712 4620 6724
rect 4172 6684 4620 6712
rect 4614 6672 4620 6684
rect 4672 6672 4678 6724
rect 5350 6672 5356 6724
rect 5408 6672 5414 6724
rect 6196 6712 6224 6820
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6788 6820 6837 6848
rect 6788 6808 6794 6820
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 7098 6848 7104 6860
rect 7059 6820 7104 6848
rect 6825 6811 6883 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 8168 6820 9321 6848
rect 8168 6808 8174 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10229 6851 10287 6857
rect 10229 6848 10241 6851
rect 9732 6820 10241 6848
rect 9732 6808 9738 6820
rect 10229 6817 10241 6820
rect 10275 6817 10287 6851
rect 10502 6848 10508 6860
rect 10463 6820 10508 6848
rect 10229 6811 10287 6817
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12124 6820 14688 6848
rect 12124 6808 12130 6820
rect 9214 6780 9220 6792
rect 9175 6752 9220 6780
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 12250 6740 12256 6792
rect 12308 6780 12314 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 12308 6752 13277 6780
rect 12308 6740 12314 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 14660 6780 14688 6820
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 14792 6820 18000 6848
rect 14792 6808 14798 6820
rect 15102 6780 15108 6792
rect 14660 6752 14964 6780
rect 15063 6752 15108 6780
rect 13265 6743 13323 6749
rect 7006 6712 7012 6724
rect 6196 6684 7012 6712
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7650 6672 7656 6724
rect 7708 6672 7714 6724
rect 9582 6712 9588 6724
rect 8404 6684 9588 6712
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 2869 6647 2927 6653
rect 2869 6644 2881 6647
rect 2556 6616 2881 6644
rect 2556 6604 2562 6616
rect 2869 6613 2881 6616
rect 2915 6613 2927 6647
rect 2869 6607 2927 6613
rect 3973 6647 4031 6653
rect 3973 6613 3985 6647
rect 4019 6644 4031 6647
rect 4706 6644 4712 6656
rect 4019 6616 4712 6644
rect 4019 6613 4031 6616
rect 3973 6607 4031 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 5684 6616 6377 6644
rect 5684 6604 5690 6616
rect 6365 6613 6377 6616
rect 6411 6644 6423 6647
rect 7282 6644 7288 6656
rect 6411 6616 7288 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 8404 6644 8432 6684
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 9950 6672 9956 6724
rect 10008 6712 10014 6724
rect 10008 6684 10994 6712
rect 10008 6672 10014 6684
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 12529 6715 12587 6721
rect 12529 6712 12541 6715
rect 12492 6684 12541 6712
rect 12492 6672 12498 6684
rect 12529 6681 12541 6684
rect 12575 6712 12587 6715
rect 14734 6712 14740 6724
rect 12575 6684 14740 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 14734 6672 14740 6684
rect 14792 6672 14798 6724
rect 8570 6644 8576 6656
rect 7432 6616 8432 6644
rect 8531 6616 8576 6644
rect 7432 6604 7438 6616
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 11422 6604 11428 6656
rect 11480 6644 11486 6656
rect 12342 6644 12348 6656
rect 11480 6616 12348 6644
rect 11480 6604 11486 6616
rect 12342 6604 12348 6616
rect 12400 6644 12406 6656
rect 13722 6644 13728 6656
rect 12400 6616 13728 6644
rect 12400 6604 12406 6616
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14936 6644 14964 6752
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 17972 6789 18000 6820
rect 17959 6783 18017 6789
rect 17959 6749 17971 6783
rect 18005 6749 18017 6783
rect 17959 6743 18017 6749
rect 16666 6712 16672 6724
rect 16606 6684 16672 6712
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 17972 6656 18000 6743
rect 18064 6712 18092 6888
rect 21082 6876 21088 6928
rect 21140 6916 21146 6928
rect 21140 6888 22048 6916
rect 21140 6876 21146 6888
rect 18785 6851 18843 6857
rect 18785 6817 18797 6851
rect 18831 6848 18843 6851
rect 19426 6848 19432 6860
rect 18831 6820 19432 6848
rect 18831 6817 18843 6820
rect 18785 6811 18843 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 19705 6851 19763 6857
rect 19705 6817 19717 6851
rect 19751 6848 19763 6851
rect 21174 6848 21180 6860
rect 19751 6820 21180 6848
rect 19751 6817 19763 6820
rect 19705 6811 19763 6817
rect 21174 6808 21180 6820
rect 21232 6848 21238 6860
rect 21913 6851 21971 6857
rect 21913 6848 21925 6851
rect 21232 6820 21925 6848
rect 21232 6808 21238 6820
rect 21913 6817 21925 6820
rect 21959 6817 21971 6851
rect 22020 6848 22048 6888
rect 23474 6876 23480 6928
rect 23532 6916 23538 6928
rect 25314 6916 25320 6928
rect 23532 6888 25320 6916
rect 23532 6876 23538 6888
rect 25314 6876 25320 6888
rect 25372 6876 25378 6928
rect 29733 6919 29791 6925
rect 29733 6885 29745 6919
rect 29779 6885 29791 6919
rect 29733 6879 29791 6885
rect 27798 6848 27804 6860
rect 22020 6820 27200 6848
rect 27759 6820 27804 6848
rect 21913 6811 21971 6817
rect 26142 6740 26148 6792
rect 26200 6780 26206 6792
rect 27172 6789 27200 6820
rect 27798 6808 27804 6820
rect 27856 6808 27862 6860
rect 27985 6851 28043 6857
rect 27985 6817 27997 6851
rect 28031 6848 28043 6851
rect 29748 6848 29776 6879
rect 28031 6820 29776 6848
rect 28031 6817 28043 6820
rect 27985 6811 28043 6817
rect 26513 6783 26571 6789
rect 26513 6780 26525 6783
rect 26200 6752 26525 6780
rect 26200 6740 26206 6752
rect 26513 6749 26525 6752
rect 26559 6749 26571 6783
rect 26513 6743 26571 6749
rect 27157 6783 27215 6789
rect 27157 6749 27169 6783
rect 27203 6749 27215 6783
rect 28442 6780 28448 6792
rect 28403 6752 28448 6780
rect 27157 6743 27215 6749
rect 28442 6740 28448 6752
rect 28500 6740 28506 6792
rect 29086 6740 29092 6792
rect 29144 6780 29150 6792
rect 29181 6783 29239 6789
rect 29181 6780 29193 6783
rect 29144 6752 29193 6780
rect 29144 6740 29150 6752
rect 29181 6749 29193 6752
rect 29227 6749 29239 6783
rect 29840 6780 29868 6956
rect 34330 6848 34336 6860
rect 30024 6820 34336 6848
rect 29917 6783 29975 6789
rect 29917 6780 29929 6783
rect 29840 6752 29929 6780
rect 29181 6743 29239 6749
rect 29917 6749 29929 6752
rect 29963 6749 29975 6783
rect 29917 6743 29975 6749
rect 19886 6712 19892 6724
rect 18064 6684 19892 6712
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 22186 6712 22192 6724
rect 21206 6684 21772 6712
rect 22147 6684 22192 6712
rect 17678 6644 17684 6656
rect 14936 6616 17684 6644
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 20898 6644 20904 6656
rect 18012 6616 20904 6644
rect 18012 6604 18018 6616
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 21450 6644 21456 6656
rect 21411 6616 21456 6644
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 21744 6644 21772 6684
rect 22186 6672 22192 6684
rect 22244 6672 22250 6724
rect 24670 6712 24676 6724
rect 23414 6684 24676 6712
rect 24670 6672 24676 6684
rect 24728 6672 24734 6724
rect 24762 6672 24768 6724
rect 24820 6712 24826 6724
rect 25041 6715 25099 6721
rect 25041 6712 25053 6715
rect 24820 6684 25053 6712
rect 24820 6672 24826 6684
rect 25041 6681 25053 6684
rect 25087 6681 25099 6715
rect 25041 6675 25099 6681
rect 25133 6715 25191 6721
rect 25133 6681 25145 6715
rect 25179 6712 25191 6715
rect 25179 6684 25360 6712
rect 25179 6681 25191 6684
rect 25133 6675 25191 6681
rect 22094 6644 22100 6656
rect 21744 6616 22100 6644
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 22278 6604 22284 6656
rect 22336 6644 22342 6656
rect 23661 6647 23719 6653
rect 23661 6644 23673 6647
rect 22336 6616 23673 6644
rect 22336 6604 22342 6616
rect 23661 6613 23673 6616
rect 23707 6613 23719 6647
rect 25332 6644 25360 6684
rect 25958 6672 25964 6724
rect 26016 6712 26022 6724
rect 26053 6715 26111 6721
rect 26053 6712 26065 6715
rect 26016 6684 26065 6712
rect 26016 6672 26022 6684
rect 26053 6681 26065 6684
rect 26099 6681 26111 6715
rect 27249 6715 27307 6721
rect 27249 6712 27261 6715
rect 26053 6675 26111 6681
rect 26160 6684 27261 6712
rect 26160 6644 26188 6684
rect 27249 6681 27261 6684
rect 27295 6681 27307 6715
rect 27249 6675 27307 6681
rect 26602 6644 26608 6656
rect 25332 6616 26188 6644
rect 26563 6616 26608 6644
rect 23661 6607 23719 6613
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 27798 6604 27804 6656
rect 27856 6644 27862 6656
rect 30024 6644 30052 6820
rect 34330 6808 34336 6820
rect 34388 6808 34394 6860
rect 33229 6783 33287 6789
rect 33229 6749 33241 6783
rect 33275 6780 33287 6783
rect 34514 6780 34520 6792
rect 33275 6752 34520 6780
rect 33275 6749 33287 6752
rect 33229 6743 33287 6749
rect 34514 6740 34520 6752
rect 34572 6740 34578 6792
rect 27856 6616 30052 6644
rect 27856 6604 27862 6616
rect 30650 6604 30656 6656
rect 30708 6644 30714 6656
rect 33321 6647 33379 6653
rect 33321 6644 33333 6647
rect 30708 6616 33333 6644
rect 30708 6604 30714 6616
rect 33321 6613 33333 6616
rect 33367 6613 33379 6647
rect 33321 6607 33379 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 5350 6440 5356 6452
rect 3476 6412 5356 6440
rect 3476 6400 3482 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6914 6440 6920 6452
rect 6043 6412 6920 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6914 6400 6920 6412
rect 6972 6440 6978 6452
rect 9030 6440 9036 6452
rect 6972 6412 9036 6440
rect 6972 6400 6978 6412
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 12250 6440 12256 6452
rect 9508 6412 12256 6440
rect 4522 6372 4528 6384
rect 4483 6344 4528 6372
rect 4522 6332 4528 6344
rect 4580 6332 4586 6384
rect 5166 6332 5172 6384
rect 5224 6332 5230 6384
rect 7006 6372 7012 6384
rect 6840 6344 7012 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 1670 6304 1676 6316
rect 1627 6276 1676 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3513 6307 3571 6313
rect 3513 6304 3525 6307
rect 3283 6276 3525 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3513 6273 3525 6276
rect 3559 6304 3571 6307
rect 3602 6304 3608 6316
rect 3559 6276 3608 6304
rect 3559 6273 3571 6276
rect 3513 6267 3571 6273
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4246 6304 4252 6316
rect 4028 6276 4252 6304
rect 4028 6264 4034 6276
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 6840 6313 6868 6344
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 9508 6372 9536 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 15930 6440 15936 6452
rect 12492 6412 15936 6440
rect 12492 6400 12498 6412
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6409 16175 6443
rect 16117 6403 16175 6409
rect 9416 6344 9536 6372
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 8202 6264 8208 6316
rect 8260 6264 8266 6316
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9416 6313 9444 6344
rect 14090 6332 14096 6384
rect 14148 6372 14154 6384
rect 14277 6375 14335 6381
rect 14277 6372 14289 6375
rect 14148 6344 14289 6372
rect 14148 6332 14154 6344
rect 14277 6341 14289 6344
rect 14323 6341 14335 6375
rect 14277 6335 14335 6341
rect 16132 6316 16160 6403
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 19334 6440 19340 6452
rect 16908 6412 19340 6440
rect 16908 6400 16914 6412
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 21542 6440 21548 6452
rect 20128 6412 21548 6440
rect 20128 6400 20134 6412
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 26602 6440 26608 6452
rect 22066 6412 26608 6440
rect 17218 6372 17224 6384
rect 16316 6344 17224 6372
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 9180 6276 9413 6304
rect 9180 6264 9186 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 10778 6264 10784 6316
rect 10836 6264 10842 6316
rect 12250 6304 12256 6316
rect 12211 6276 12256 6304
rect 12250 6264 12256 6276
rect 12308 6264 12314 6316
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 15286 6264 15292 6316
rect 15344 6304 15350 6316
rect 15838 6304 15844 6316
rect 15344 6276 15844 6304
rect 15344 6264 15350 6276
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 16114 6264 16120 6316
rect 16172 6264 16178 6316
rect 16316 6313 16344 6344
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 22066 6372 22094 6412
rect 26602 6400 26608 6412
rect 26660 6400 26666 6452
rect 27246 6440 27252 6452
rect 27207 6412 27252 6440
rect 27246 6400 27252 6412
rect 27304 6400 27310 6452
rect 27890 6440 27896 6452
rect 27851 6412 27896 6440
rect 27890 6400 27896 6412
rect 27948 6400 27954 6452
rect 29178 6440 29184 6452
rect 29139 6412 29184 6440
rect 29178 6400 29184 6412
rect 29236 6400 29242 6452
rect 29822 6440 29828 6452
rect 29783 6412 29828 6440
rect 29822 6400 29828 6412
rect 29880 6400 29886 6452
rect 23014 6372 23020 6384
rect 20930 6344 22094 6372
rect 22975 6344 23020 6372
rect 23014 6332 23020 6344
rect 23072 6332 23078 6384
rect 23109 6375 23167 6381
rect 23109 6341 23121 6375
rect 23155 6372 23167 6375
rect 28537 6375 28595 6381
rect 28537 6372 28549 6375
rect 23155 6344 28549 6372
rect 23155 6341 23167 6344
rect 23109 6335 23167 6341
rect 28537 6341 28549 6344
rect 28583 6341 28595 6375
rect 28537 6335 28595 6341
rect 28902 6332 28908 6384
rect 28960 6372 28966 6384
rect 30374 6372 30380 6384
rect 28960 6344 30380 6372
rect 28960 6332 28966 6344
rect 30374 6332 30380 6344
rect 30432 6372 30438 6384
rect 30432 6344 30604 6372
rect 30432 6332 30438 6344
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6273 16359 6307
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 16301 6267 16359 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 18230 6264 18236 6316
rect 18288 6264 18294 6316
rect 20990 6264 20996 6316
rect 21048 6304 21054 6316
rect 21453 6308 21511 6313
rect 21284 6307 21511 6308
rect 21284 6304 21465 6307
rect 21048 6280 21465 6304
rect 21048 6276 21312 6280
rect 21048 6264 21054 6276
rect 21453 6273 21465 6280
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 22281 6307 22339 6313
rect 22281 6273 22293 6307
rect 22327 6304 22339 6307
rect 22462 6304 22468 6316
rect 22327 6276 22468 6304
rect 22327 6273 22339 6276
rect 22281 6267 22339 6273
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 24486 6304 24492 6316
rect 24447 6276 24492 6304
rect 24486 6264 24492 6276
rect 24544 6264 24550 6316
rect 24854 6264 24860 6316
rect 24912 6264 24918 6316
rect 25038 6264 25044 6316
rect 25096 6304 25102 6316
rect 25133 6307 25191 6313
rect 25133 6304 25145 6307
rect 25096 6276 25145 6304
rect 25096 6264 25102 6276
rect 25133 6273 25145 6276
rect 25179 6273 25191 6307
rect 25133 6267 25191 6273
rect 25777 6307 25835 6313
rect 25777 6273 25789 6307
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 6546 6236 6552 6248
rect 2280 6208 6552 6236
rect 2280 6196 2286 6208
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 7098 6236 7104 6248
rect 7011 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6236 7162 6248
rect 9677 6239 9735 6245
rect 7156 6208 8708 6236
rect 7156 6196 7162 6208
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2774 6168 2780 6180
rect 1811 6140 2780 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2774 6128 2780 6140
rect 2832 6128 2838 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 8352 6140 8585 6168
rect 8352 6128 8358 6140
rect 8573 6137 8585 6140
rect 8619 6137 8631 6171
rect 8573 6131 8631 6137
rect 2501 6103 2559 6109
rect 2501 6069 2513 6103
rect 2547 6100 2559 6103
rect 2866 6100 2872 6112
rect 2547 6072 2872 6100
rect 2547 6069 2559 6072
rect 2501 6063 2559 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 5166 6100 5172 6112
rect 3743 6072 5172 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 8202 6100 8208 6112
rect 6696 6072 8208 6100
rect 6696 6060 6702 6072
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8680 6100 8708 6208
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 10686 6236 10692 6248
rect 9723 6208 10692 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 16758 6236 16764 6248
rect 12575 6208 16764 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 17126 6236 17132 6248
rect 17087 6208 17132 6236
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 19242 6236 19248 6248
rect 17276 6208 19248 6236
rect 17276 6196 17282 6208
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 19392 6208 19441 6236
rect 19392 6196 19398 6208
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19429 6199 19487 6205
rect 19705 6239 19763 6245
rect 19705 6205 19717 6239
rect 19751 6236 19763 6239
rect 23566 6236 23572 6248
rect 19751 6208 23572 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 23566 6196 23572 6208
rect 23624 6196 23630 6248
rect 24029 6239 24087 6245
rect 24029 6205 24041 6239
rect 24075 6236 24087 6239
rect 24872 6236 24900 6264
rect 24075 6208 24900 6236
rect 25792 6236 25820 6267
rect 25866 6264 25872 6316
rect 25924 6304 25930 6316
rect 26418 6304 26424 6316
rect 25924 6276 25969 6304
rect 26379 6276 26424 6304
rect 25924 6264 25930 6276
rect 26418 6264 26424 6276
rect 26476 6264 26482 6316
rect 27157 6307 27215 6313
rect 27157 6304 27169 6307
rect 26620 6276 27169 6304
rect 26142 6236 26148 6248
rect 25792 6208 26148 6236
rect 24075 6205 24087 6208
rect 24029 6199 24087 6205
rect 26142 6196 26148 6208
rect 26200 6196 26206 6248
rect 12158 6168 12164 6180
rect 10704 6140 12164 6168
rect 10704 6100 10732 6140
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 18322 6128 18328 6180
rect 18380 6168 18386 6180
rect 18601 6171 18659 6177
rect 18601 6168 18613 6171
rect 18380 6140 18613 6168
rect 18380 6128 18386 6140
rect 18601 6137 18613 6140
rect 18647 6137 18659 6171
rect 18601 6131 18659 6137
rect 20714 6128 20720 6180
rect 20772 6168 20778 6180
rect 21174 6168 21180 6180
rect 20772 6140 21180 6168
rect 20772 6128 20778 6140
rect 21174 6128 21180 6140
rect 21232 6168 21238 6180
rect 22094 6168 22100 6180
rect 21232 6140 22100 6168
rect 21232 6128 21238 6140
rect 22094 6128 22100 6140
rect 22152 6128 22158 6180
rect 22186 6128 22192 6180
rect 22244 6168 22250 6180
rect 22244 6140 22508 6168
rect 22244 6128 22250 6140
rect 11146 6100 11152 6112
rect 8680 6072 10732 6100
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 16666 6100 16672 6112
rect 14700 6072 16672 6100
rect 14700 6060 14706 6072
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22373 6103 22431 6109
rect 22373 6100 22385 6103
rect 22060 6072 22385 6100
rect 22060 6060 22066 6072
rect 22373 6069 22385 6072
rect 22419 6069 22431 6103
rect 22480 6100 22508 6140
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 24854 6168 24860 6180
rect 23072 6140 24860 6168
rect 23072 6128 23078 6140
rect 24854 6128 24860 6140
rect 24912 6128 24918 6180
rect 25774 6128 25780 6180
rect 25832 6168 25838 6180
rect 26418 6168 26424 6180
rect 25832 6140 26424 6168
rect 25832 6128 25838 6140
rect 26418 6128 26424 6140
rect 26476 6168 26482 6180
rect 26620 6168 26648 6276
rect 27157 6273 27169 6276
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 27801 6307 27859 6313
rect 27801 6304 27813 6307
rect 27304 6276 27813 6304
rect 27304 6264 27310 6276
rect 27801 6273 27813 6276
rect 27847 6273 27859 6307
rect 27801 6267 27859 6273
rect 28445 6307 28503 6313
rect 28445 6273 28457 6307
rect 28491 6273 28503 6307
rect 28445 6267 28503 6273
rect 29089 6307 29147 6313
rect 29089 6273 29101 6307
rect 29135 6304 29147 6307
rect 29454 6304 29460 6316
rect 29135 6276 29460 6304
rect 29135 6273 29147 6276
rect 29089 6267 29147 6273
rect 26694 6196 26700 6248
rect 26752 6236 26758 6248
rect 28460 6236 28488 6267
rect 29454 6264 29460 6276
rect 29512 6264 29518 6316
rect 30576 6313 30604 6344
rect 29733 6307 29791 6313
rect 29733 6273 29745 6307
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 30561 6307 30619 6313
rect 30561 6273 30573 6307
rect 30607 6273 30619 6307
rect 30561 6267 30619 6273
rect 26752 6208 28488 6236
rect 26752 6196 26758 6208
rect 29086 6168 29092 6180
rect 26476 6140 29092 6168
rect 26476 6128 26482 6140
rect 29086 6128 29092 6140
rect 29144 6128 29150 6180
rect 29748 6168 29776 6267
rect 36722 6168 36728 6180
rect 29748 6140 36728 6168
rect 36722 6128 36728 6140
rect 36780 6128 36786 6180
rect 24581 6103 24639 6109
rect 24581 6100 24593 6103
rect 22480 6072 24593 6100
rect 22373 6063 22431 6069
rect 24581 6069 24593 6072
rect 24627 6069 24639 6103
rect 24581 6063 24639 6069
rect 24762 6060 24768 6112
rect 24820 6100 24826 6112
rect 25225 6103 25283 6109
rect 25225 6100 25237 6103
rect 24820 6072 25237 6100
rect 24820 6060 24826 6072
rect 25225 6069 25237 6072
rect 25271 6069 25283 6103
rect 26510 6100 26516 6112
rect 26471 6072 26516 6100
rect 25225 6063 25283 6069
rect 26510 6060 26516 6072
rect 26568 6060 26574 6112
rect 30377 6103 30435 6109
rect 30377 6069 30389 6103
rect 30423 6100 30435 6103
rect 32490 6100 32496 6112
rect 30423 6072 32496 6100
rect 30423 6069 30435 6072
rect 30377 6063 30435 6069
rect 32490 6060 32496 6072
rect 32548 6060 32554 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 6270 5896 6276 5908
rect 3200 5868 6276 5896
rect 3200 5856 3206 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 8570 5896 8576 5908
rect 6564 5868 8576 5896
rect 2869 5763 2927 5769
rect 2869 5729 2881 5763
rect 2915 5760 2927 5763
rect 3878 5760 3884 5772
rect 2915 5732 3884 5760
rect 2915 5729 2927 5732
rect 2869 5723 2927 5729
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 6564 5760 6592 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 8904 5868 10456 5896
rect 8904 5856 8910 5868
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 10428 5828 10456 5868
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10836 5868 13492 5896
rect 10836 5856 10842 5868
rect 11054 5828 11060 5840
rect 8260 5800 9260 5828
rect 10428 5800 11060 5828
rect 8260 5788 8266 5800
rect 4295 5732 6592 5760
rect 6641 5763 6699 5769
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 7006 5760 7012 5772
rect 6687 5732 7012 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7340 5732 8156 5760
rect 7340 5720 7346 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 2498 5692 2504 5704
rect 1627 5664 2504 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 2593 5655 2651 5661
rect 14 5516 20 5568
rect 72 5556 78 5568
rect 1765 5559 1823 5565
rect 1765 5556 1777 5559
rect 72 5528 1777 5556
rect 72 5516 78 5528
rect 1765 5525 1777 5528
rect 1811 5525 1823 5559
rect 2608 5556 2636 5655
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 5994 5692 6000 5704
rect 5776 5664 6000 5692
rect 5776 5652 5782 5664
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 8128 5692 8156 5732
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 9122 5760 9128 5772
rect 8444 5732 9128 5760
rect 8444 5720 8450 5732
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9232 5760 9260 5800
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 10410 5760 10416 5772
rect 9232 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 10962 5760 10968 5772
rect 10919 5732 10968 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5760 11483 5763
rect 11471 5732 13400 5760
rect 11471 5729 11483 5732
rect 11425 5723 11483 5729
rect 8128 5664 8616 5692
rect 3988 5624 4016 5652
rect 4246 5624 4252 5636
rect 3988 5596 4252 5624
rect 4246 5584 4252 5596
rect 4304 5584 4310 5636
rect 4798 5584 4804 5636
rect 4856 5584 4862 5636
rect 6638 5624 6644 5636
rect 5644 5596 6644 5624
rect 5644 5556 5672 5596
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 6917 5627 6975 5633
rect 6917 5593 6929 5627
rect 6963 5593 6975 5627
rect 8478 5624 8484 5636
rect 8142 5596 8484 5624
rect 6917 5587 6975 5593
rect 2608 5528 5672 5556
rect 5721 5559 5779 5565
rect 1765 5519 1823 5525
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 6730 5556 6736 5568
rect 5767 5528 6736 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 6932 5556 6960 5587
rect 8478 5584 8484 5596
rect 8536 5584 8542 5636
rect 8588 5624 8616 5664
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 8588 5596 9413 5624
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9401 5587 9459 5593
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 11701 5627 11759 5633
rect 9548 5596 9890 5624
rect 9548 5584 9554 5596
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 11974 5624 11980 5636
rect 11747 5596 11980 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 7834 5556 7840 5568
rect 6932 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 11790 5556 11796 5568
rect 8435 5528 11796 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 13372 5556 13400 5732
rect 13464 5633 13492 5868
rect 13630 5856 13636 5908
rect 13688 5896 13694 5908
rect 22738 5896 22744 5908
rect 13688 5868 22744 5896
rect 13688 5856 13694 5868
rect 22738 5856 22744 5868
rect 22796 5856 22802 5908
rect 24670 5856 24676 5908
rect 24728 5896 24734 5908
rect 27157 5899 27215 5905
rect 27157 5896 27169 5899
rect 24728 5868 27169 5896
rect 24728 5856 24734 5868
rect 27157 5865 27169 5868
rect 27203 5865 27215 5899
rect 27157 5859 27215 5865
rect 28994 5856 29000 5908
rect 29052 5896 29058 5908
rect 29089 5899 29147 5905
rect 29089 5896 29101 5899
rect 29052 5868 29101 5896
rect 29052 5856 29058 5868
rect 29089 5865 29101 5868
rect 29135 5865 29147 5899
rect 29089 5859 29147 5865
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 13596 5800 15240 5828
rect 13596 5788 13602 5800
rect 15212 5760 15240 5800
rect 16758 5788 16764 5840
rect 16816 5828 16822 5840
rect 17681 5831 17739 5837
rect 17681 5828 17693 5831
rect 16816 5800 17693 5828
rect 16816 5788 16822 5800
rect 17681 5797 17693 5800
rect 17727 5797 17739 5831
rect 17681 5791 17739 5797
rect 18417 5831 18475 5837
rect 18417 5797 18429 5831
rect 18463 5797 18475 5831
rect 18417 5791 18475 5797
rect 15838 5760 15844 5772
rect 15212 5732 15844 5760
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 15930 5720 15936 5772
rect 15988 5760 15994 5772
rect 16853 5763 16911 5769
rect 15988 5732 16620 5760
rect 15988 5720 15994 5732
rect 14642 5692 14648 5704
rect 14603 5664 14648 5692
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 15102 5692 15108 5704
rect 15063 5664 15108 5692
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 16482 5652 16488 5704
rect 16540 5652 16546 5704
rect 16592 5692 16620 5732
rect 16853 5729 16865 5763
rect 16899 5760 16911 5763
rect 17034 5760 17040 5772
rect 16899 5732 17040 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 18432 5760 18460 5791
rect 21082 5788 21088 5840
rect 21140 5828 21146 5840
rect 26513 5831 26571 5837
rect 26513 5828 26525 5831
rect 21140 5800 22094 5828
rect 21140 5788 21146 5800
rect 17144 5732 18460 5760
rect 17144 5692 17172 5732
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 19392 5732 19809 5760
rect 19392 5720 19398 5732
rect 19797 5729 19809 5732
rect 19843 5760 19855 5763
rect 20714 5760 20720 5772
rect 19843 5732 20720 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 20714 5720 20720 5732
rect 20772 5720 20778 5772
rect 22066 5760 22094 5800
rect 26344 5800 26525 5828
rect 26344 5772 26372 5800
rect 26513 5797 26525 5800
rect 26559 5797 26571 5831
rect 26513 5791 26571 5797
rect 29733 5831 29791 5837
rect 29733 5797 29745 5831
rect 29779 5828 29791 5831
rect 32306 5828 32312 5840
rect 29779 5800 32312 5828
rect 29779 5797 29791 5800
rect 29733 5791 29791 5797
rect 32306 5788 32312 5800
rect 32364 5788 32370 5840
rect 24302 5760 24308 5772
rect 22066 5732 24308 5760
rect 24302 5720 24308 5732
rect 24360 5720 24366 5772
rect 24673 5763 24731 5769
rect 24673 5729 24685 5763
rect 24719 5760 24731 5763
rect 24854 5760 24860 5772
rect 24719 5732 24860 5760
rect 24719 5729 24731 5732
rect 24673 5723 24731 5729
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 24946 5720 24952 5772
rect 25004 5760 25010 5772
rect 25869 5763 25927 5769
rect 25869 5760 25881 5763
rect 25004 5732 25881 5760
rect 25004 5720 25010 5732
rect 25869 5729 25881 5732
rect 25915 5729 25927 5763
rect 25869 5723 25927 5729
rect 26326 5720 26332 5772
rect 26384 5720 26390 5772
rect 27522 5760 27528 5772
rect 26620 5732 27528 5760
rect 17494 5692 17500 5704
rect 16592 5664 17172 5692
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 15286 5624 15292 5636
rect 13495 5596 15292 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 15378 5584 15384 5636
rect 15436 5624 15442 5636
rect 18248 5624 18276 5655
rect 22002 5652 22008 5704
rect 22060 5692 22066 5704
rect 23753 5695 23811 5701
rect 22060 5664 22105 5692
rect 22664 5664 23704 5692
rect 22060 5652 22066 5664
rect 15436 5596 15481 5624
rect 16776 5596 18276 5624
rect 20073 5627 20131 5633
rect 15436 5584 15442 5596
rect 14366 5556 14372 5568
rect 13372 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 14461 5559 14519 5565
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 16776 5556 16804 5596
rect 20073 5593 20085 5627
rect 20119 5593 20131 5627
rect 22664 5624 22692 5664
rect 21298 5596 22692 5624
rect 22741 5627 22799 5633
rect 20073 5587 20131 5593
rect 22741 5593 22753 5627
rect 22787 5593 22799 5627
rect 23676 5624 23704 5664
rect 23753 5661 23765 5695
rect 23799 5692 23811 5695
rect 23842 5692 23848 5704
rect 23799 5664 23848 5692
rect 23799 5661 23811 5664
rect 23753 5655 23811 5661
rect 23842 5652 23848 5664
rect 23900 5652 23906 5704
rect 25317 5695 25375 5701
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25406 5692 25412 5704
rect 25363 5664 25412 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 25682 5652 25688 5704
rect 25740 5692 25746 5704
rect 25777 5695 25835 5701
rect 25777 5692 25789 5695
rect 25740 5664 25789 5692
rect 25740 5652 25746 5664
rect 25777 5661 25789 5664
rect 25823 5661 25835 5695
rect 25777 5655 25835 5661
rect 26421 5695 26479 5701
rect 26421 5661 26433 5695
rect 26467 5694 26479 5695
rect 26467 5692 26556 5694
rect 26620 5692 26648 5732
rect 27522 5720 27528 5732
rect 27580 5720 27586 5772
rect 27724 5732 28028 5760
rect 26467 5666 26648 5692
rect 26467 5661 26479 5666
rect 26528 5664 26648 5666
rect 26421 5655 26479 5661
rect 26786 5652 26792 5704
rect 26844 5692 26850 5704
rect 27724 5701 27752 5732
rect 28000 5704 28028 5732
rect 28258 5720 28264 5772
rect 28316 5760 28322 5772
rect 29270 5760 29276 5772
rect 28316 5732 29276 5760
rect 28316 5720 28322 5732
rect 29270 5720 29276 5732
rect 29328 5720 29334 5772
rect 27065 5695 27123 5701
rect 27065 5692 27077 5695
rect 26844 5664 27077 5692
rect 26844 5652 26850 5664
rect 27065 5661 27077 5664
rect 27111 5692 27123 5695
rect 27709 5695 27767 5701
rect 27709 5692 27721 5695
rect 27111 5664 27721 5692
rect 27111 5661 27123 5664
rect 27065 5655 27123 5661
rect 27709 5661 27721 5664
rect 27755 5661 27767 5695
rect 27709 5655 27767 5661
rect 27798 5652 27804 5704
rect 27856 5692 27862 5704
rect 27856 5664 27901 5692
rect 27856 5652 27862 5664
rect 27982 5652 27988 5704
rect 28040 5692 28046 5704
rect 28353 5695 28411 5701
rect 28353 5692 28365 5695
rect 28040 5664 28365 5692
rect 28040 5652 28046 5664
rect 28353 5661 28365 5664
rect 28399 5692 28411 5695
rect 28902 5692 28908 5704
rect 28399 5664 28908 5692
rect 28399 5661 28411 5664
rect 28353 5655 28411 5661
rect 28902 5652 28908 5664
rect 28960 5652 28966 5704
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 29086 5692 29092 5704
rect 29043 5664 29092 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 29086 5652 29092 5664
rect 29144 5692 29150 5704
rect 29638 5692 29644 5704
rect 29144 5664 29644 5692
rect 29144 5652 29150 5664
rect 29638 5652 29644 5664
rect 29696 5652 29702 5704
rect 29914 5692 29920 5704
rect 29875 5664 29920 5692
rect 29914 5652 29920 5664
rect 29972 5652 29978 5704
rect 30374 5692 30380 5704
rect 30335 5664 30380 5692
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 31018 5692 31024 5704
rect 30979 5664 31024 5692
rect 31018 5652 31024 5664
rect 31076 5652 31082 5704
rect 31846 5692 31852 5704
rect 31807 5664 31852 5692
rect 31846 5652 31852 5664
rect 31904 5652 31910 5704
rect 35529 5695 35587 5701
rect 35529 5661 35541 5695
rect 35575 5661 35587 5695
rect 38010 5692 38016 5704
rect 37971 5664 38016 5692
rect 35529 5655 35587 5661
rect 23676 5596 24716 5624
rect 22741 5587 22799 5593
rect 14507 5528 16804 5556
rect 20088 5556 20116 5587
rect 21082 5556 21088 5568
rect 20088 5528 21088 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 21542 5556 21548 5568
rect 21503 5528 21548 5556
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 22002 5516 22008 5568
rect 22060 5556 22066 5568
rect 22756 5556 22784 5587
rect 22060 5528 22784 5556
rect 22060 5516 22066 5528
rect 23658 5516 23664 5568
rect 23716 5556 23722 5568
rect 23845 5559 23903 5565
rect 23845 5556 23857 5559
rect 23716 5528 23857 5556
rect 23716 5516 23722 5528
rect 23845 5525 23857 5528
rect 23891 5525 23903 5559
rect 24688 5556 24716 5596
rect 24762 5584 24768 5636
rect 24820 5624 24826 5636
rect 24820 5596 24865 5624
rect 24820 5584 24826 5596
rect 27338 5584 27344 5636
rect 27396 5624 27402 5636
rect 28445 5627 28503 5633
rect 28445 5624 28457 5627
rect 27396 5596 28457 5624
rect 27396 5584 27402 5596
rect 28445 5593 28457 5596
rect 28491 5593 28503 5627
rect 28445 5587 28503 5593
rect 28534 5584 28540 5636
rect 28592 5624 28598 5636
rect 30469 5627 30527 5633
rect 30469 5624 30481 5627
rect 28592 5596 30481 5624
rect 28592 5584 28598 5596
rect 30469 5593 30481 5596
rect 30515 5593 30527 5627
rect 30469 5587 30527 5593
rect 31113 5627 31171 5633
rect 31113 5593 31125 5627
rect 31159 5624 31171 5627
rect 35544 5624 35572 5655
rect 38010 5652 38016 5664
rect 38068 5652 38074 5704
rect 31159 5596 35572 5624
rect 31159 5593 31171 5596
rect 31113 5587 31171 5593
rect 30558 5556 30564 5568
rect 24688 5528 30564 5556
rect 23845 5519 23903 5525
rect 30558 5516 30564 5528
rect 30616 5516 30622 5568
rect 31665 5559 31723 5565
rect 31665 5525 31677 5559
rect 31711 5556 31723 5559
rect 34606 5556 34612 5568
rect 31711 5528 34612 5556
rect 31711 5525 31723 5528
rect 31665 5519 31723 5525
rect 34606 5516 34612 5528
rect 34664 5516 34670 5568
rect 35345 5559 35403 5565
rect 35345 5525 35357 5559
rect 35391 5556 35403 5559
rect 38010 5556 38016 5568
rect 35391 5528 38016 5556
rect 35391 5525 35403 5528
rect 35345 5519 35403 5525
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 38194 5556 38200 5568
rect 38155 5528 38200 5556
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 11146 5352 11152 5364
rect 8220 5324 11152 5352
rect 2746 5256 5014 5284
rect 1578 5216 1584 5228
rect 1539 5188 1584 5216
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2590 5176 2596 5228
rect 2648 5216 2654 5228
rect 2746 5216 2774 5256
rect 7006 5244 7012 5296
rect 7064 5284 7070 5296
rect 7285 5287 7343 5293
rect 7285 5284 7297 5287
rect 7064 5256 7297 5284
rect 7064 5244 7070 5256
rect 7285 5253 7297 5256
rect 7331 5253 7343 5287
rect 7285 5247 7343 5253
rect 2648 5188 2774 5216
rect 2869 5219 2927 5225
rect 2648 5176 2654 5188
rect 2869 5185 2881 5219
rect 2915 5185 2927 5219
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 2869 5179 2927 5185
rect 658 4972 664 5024
rect 716 5012 722 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 716 4984 1777 5012
rect 716 4972 722 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 2884 5012 2912 5179
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5920 5188 6561 5216
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 4062 5148 4068 5160
rect 3743 5120 4068 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4571 5120 5672 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 5644 5092 5672 5120
rect 5626 5040 5632 5092
rect 5684 5040 5690 5092
rect 5534 5012 5540 5024
rect 2884 4984 5540 5012
rect 1765 4975 1823 4981
rect 5534 4972 5540 4984
rect 5592 5012 5598 5024
rect 5920 5012 5948 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6052 5120 6097 5148
rect 6052 5108 6058 5120
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 8220 5080 8248 5324
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 14642 5352 14648 5364
rect 12544 5324 14648 5352
rect 8662 5244 8668 5296
rect 8720 5284 8726 5296
rect 8720 5256 9154 5284
rect 8720 5244 8726 5256
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 12544 5293 12572 5324
rect 14642 5312 14648 5324
rect 14700 5312 14706 5364
rect 22646 5352 22652 5364
rect 14752 5324 22652 5352
rect 10413 5287 10471 5293
rect 10413 5284 10425 5287
rect 10376 5256 10425 5284
rect 10376 5244 10382 5256
rect 10413 5253 10425 5256
rect 10459 5253 10471 5287
rect 10413 5247 10471 5253
rect 12529 5287 12587 5293
rect 12529 5253 12541 5287
rect 12575 5253 12587 5287
rect 12529 5247 12587 5253
rect 13170 5244 13176 5296
rect 13228 5244 13234 5296
rect 14752 5293 14780 5324
rect 22646 5312 22652 5324
rect 22704 5312 22710 5364
rect 23198 5312 23204 5364
rect 23256 5352 23262 5364
rect 25961 5355 26019 5361
rect 25961 5352 25973 5355
rect 23256 5324 25973 5352
rect 23256 5312 23262 5324
rect 25961 5321 25973 5324
rect 26007 5321 26019 5355
rect 25961 5315 26019 5321
rect 26602 5312 26608 5364
rect 26660 5352 26666 5364
rect 29641 5355 29699 5361
rect 29641 5352 29653 5355
rect 26660 5324 27292 5352
rect 26660 5312 26666 5324
rect 14737 5287 14795 5293
rect 14737 5253 14749 5287
rect 14783 5253 14795 5287
rect 14737 5247 14795 5253
rect 15746 5244 15752 5296
rect 15804 5244 15810 5296
rect 19058 5284 19064 5296
rect 18446 5256 19064 5284
rect 19058 5244 19064 5256
rect 19116 5244 19122 5296
rect 19334 5284 19340 5296
rect 19168 5256 19340 5284
rect 8386 5216 8392 5228
rect 8347 5188 8392 5216
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11514 5216 11520 5228
rect 11195 5188 11520 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 12250 5216 12256 5228
rect 12211 5188 12256 5216
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 19168 5225 19196 5256
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 19426 5244 19432 5296
rect 19484 5284 19490 5296
rect 22278 5284 22284 5296
rect 19484 5256 19529 5284
rect 20654 5256 22284 5284
rect 19484 5244 19490 5256
rect 22278 5244 22284 5256
rect 22336 5244 22342 5296
rect 25038 5284 25044 5296
rect 23506 5256 25044 5284
rect 25038 5244 25044 5256
rect 25096 5244 25102 5296
rect 27264 5293 27292 5324
rect 27356 5324 29653 5352
rect 27356 5293 27384 5324
rect 29641 5321 29653 5324
rect 29687 5321 29699 5355
rect 31570 5352 31576 5364
rect 31531 5324 31576 5352
rect 29641 5315 29699 5321
rect 31570 5312 31576 5324
rect 31628 5312 31634 5364
rect 27249 5287 27307 5293
rect 27249 5253 27261 5287
rect 27295 5253 27307 5287
rect 27249 5247 27307 5253
rect 27341 5287 27399 5293
rect 27341 5253 27353 5287
rect 27387 5253 27399 5287
rect 27341 5247 27399 5253
rect 27893 5287 27951 5293
rect 27893 5253 27905 5287
rect 27939 5284 27951 5287
rect 28258 5284 28264 5296
rect 27939 5256 28264 5284
rect 27939 5253 27951 5256
rect 27893 5247 27951 5253
rect 28258 5244 28264 5256
rect 28316 5244 28322 5296
rect 28534 5284 28540 5296
rect 28495 5256 28540 5284
rect 28534 5244 28540 5256
rect 28592 5244 28598 5296
rect 28810 5244 28816 5296
rect 28868 5284 28874 5296
rect 30285 5287 30343 5293
rect 30285 5284 30297 5287
rect 28868 5256 30297 5284
rect 28868 5244 28874 5256
rect 30285 5253 30297 5256
rect 30331 5253 30343 5287
rect 30285 5247 30343 5253
rect 30466 5244 30472 5296
rect 30524 5284 30530 5296
rect 32582 5284 32588 5296
rect 30524 5256 32588 5284
rect 30524 5244 30530 5256
rect 32582 5244 32588 5256
rect 32640 5244 32646 5296
rect 19153 5219 19211 5225
rect 19153 5185 19165 5219
rect 19199 5185 19211 5219
rect 21266 5216 21272 5228
rect 19153 5179 19211 5185
rect 20824 5188 21272 5216
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5148 8723 5151
rect 8711 5120 10364 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 6144 5052 8248 5080
rect 10336 5080 10364 5120
rect 12618 5108 12624 5160
rect 12676 5148 12682 5160
rect 12676 5120 13768 5148
rect 12676 5108 12682 5120
rect 10336 5052 11100 5080
rect 6144 5040 6150 5052
rect 5592 4984 5948 5012
rect 5592 4972 5598 4984
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 6604 4984 10977 5012
rect 6604 4972 6610 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 11072 5012 11100 5052
rect 13262 5012 13268 5024
rect 11072 4984 13268 5012
rect 10965 4975 11023 4981
rect 13262 4972 13268 4984
rect 13320 5012 13326 5024
rect 13630 5012 13636 5024
rect 13320 4984 13636 5012
rect 13320 4972 13326 4984
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13740 5012 13768 5120
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 14424 5120 14473 5148
rect 14424 5108 14430 5120
rect 14461 5117 14473 5120
rect 14507 5148 14519 5151
rect 15102 5148 15108 5160
rect 14507 5120 15108 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 15102 5108 15108 5120
rect 15160 5148 15166 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 15160 5120 16957 5148
rect 15160 5108 15166 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17221 5151 17279 5157
rect 17221 5117 17233 5151
rect 17267 5148 17279 5151
rect 17862 5148 17868 5160
rect 17267 5120 17868 5148
rect 17267 5117 17279 5120
rect 17221 5111 17279 5117
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 20824 5148 20852 5188
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 22002 5216 22008 5228
rect 21963 5188 22008 5216
rect 22002 5176 22008 5188
rect 22060 5176 22066 5228
rect 24486 5176 24492 5228
rect 24544 5216 24550 5228
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 24544 5188 24593 5216
rect 24544 5176 24550 5188
rect 24581 5185 24593 5188
rect 24627 5185 24639 5219
rect 24581 5179 24639 5185
rect 25225 5219 25283 5225
rect 25225 5185 25237 5219
rect 25271 5216 25283 5219
rect 25498 5216 25504 5228
rect 25271 5188 25504 5216
rect 25271 5185 25283 5188
rect 25225 5179 25283 5185
rect 25498 5176 25504 5188
rect 25556 5176 25562 5228
rect 25869 5219 25927 5225
rect 25869 5185 25881 5219
rect 25915 5216 25927 5219
rect 26418 5216 26424 5228
rect 25915 5188 26424 5216
rect 25915 5185 25927 5188
rect 25869 5179 25927 5185
rect 26418 5176 26424 5188
rect 26476 5176 26482 5228
rect 29546 5216 29552 5228
rect 29507 5188 29552 5216
rect 29546 5176 29552 5188
rect 29604 5176 29610 5228
rect 29638 5176 29644 5228
rect 29696 5216 29702 5228
rect 30193 5219 30251 5225
rect 30193 5216 30205 5219
rect 29696 5188 30205 5216
rect 29696 5176 29702 5188
rect 30193 5185 30205 5188
rect 30239 5216 30251 5219
rect 30837 5219 30895 5225
rect 30837 5216 30849 5219
rect 30239 5188 30849 5216
rect 30239 5185 30251 5188
rect 30193 5179 30251 5185
rect 30837 5185 30849 5188
rect 30883 5216 30895 5219
rect 31202 5216 31208 5228
rect 30883 5188 31208 5216
rect 30883 5185 30895 5188
rect 30837 5179 30895 5185
rect 31202 5176 31208 5188
rect 31260 5176 31266 5228
rect 31481 5219 31539 5225
rect 31481 5185 31493 5219
rect 31527 5185 31539 5219
rect 31481 5179 31539 5185
rect 18248 5120 20852 5148
rect 20901 5151 20959 5157
rect 13998 5080 14004 5092
rect 13959 5052 14004 5080
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 13740 4984 16221 5012
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 16298 4972 16304 5024
rect 16356 5012 16362 5024
rect 18248 5012 18276 5120
rect 20901 5117 20913 5151
rect 20947 5148 20959 5151
rect 21082 5148 21088 5160
rect 20947 5120 21088 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21082 5108 21088 5120
rect 21140 5108 21146 5160
rect 21174 5108 21180 5160
rect 21232 5148 21238 5160
rect 22281 5151 22339 5157
rect 22281 5148 22293 5151
rect 21232 5120 22293 5148
rect 21232 5108 21238 5120
rect 22281 5117 22293 5120
rect 22327 5148 22339 5151
rect 26142 5148 26148 5160
rect 22327 5136 25728 5148
rect 25976 5136 26148 5148
rect 22327 5120 26148 5136
rect 22327 5117 22339 5120
rect 22281 5111 22339 5117
rect 25700 5108 26004 5120
rect 26142 5108 26148 5120
rect 26200 5108 26206 5160
rect 28442 5148 28448 5160
rect 28403 5120 28448 5148
rect 28442 5108 28448 5120
rect 28500 5108 28506 5160
rect 31496 5148 31524 5179
rect 31662 5176 31668 5228
rect 31720 5216 31726 5228
rect 32309 5219 32367 5225
rect 32309 5216 32321 5219
rect 31720 5188 32321 5216
rect 31720 5176 31726 5188
rect 32309 5185 32321 5188
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 28552 5120 31524 5148
rect 18693 5083 18751 5089
rect 18693 5049 18705 5083
rect 18739 5080 18751 5083
rect 18782 5080 18788 5092
rect 18739 5052 18788 5080
rect 18739 5049 18751 5052
rect 18693 5043 18751 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 23474 5040 23480 5092
rect 23532 5080 23538 5092
rect 24673 5083 24731 5089
rect 24673 5080 24685 5083
rect 23532 5052 24685 5080
rect 23532 5040 23538 5052
rect 24673 5049 24685 5052
rect 24719 5049 24731 5083
rect 28552 5080 28580 5120
rect 24673 5043 24731 5049
rect 24780 5052 28580 5080
rect 16356 4984 18276 5012
rect 16356 4972 16362 4984
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 23566 5012 23572 5024
rect 18656 4984 23572 5012
rect 18656 4972 18662 4984
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 23750 5012 23756 5024
rect 23711 4984 23756 5012
rect 23750 4972 23756 4984
rect 23808 4972 23814 5024
rect 24026 4972 24032 5024
rect 24084 5012 24090 5024
rect 24780 5012 24808 5052
rect 28994 5040 29000 5092
rect 29052 5080 29058 5092
rect 31018 5080 31024 5092
rect 29052 5052 31024 5080
rect 29052 5040 29058 5052
rect 31018 5040 31024 5052
rect 31076 5040 31082 5092
rect 25314 5012 25320 5024
rect 24084 4984 24808 5012
rect 25275 4984 25320 5012
rect 24084 4972 24090 4984
rect 25314 4972 25320 4984
rect 25372 4972 25378 5024
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 29822 5012 29828 5024
rect 28868 4984 29828 5012
rect 28868 4972 28874 4984
rect 29822 4972 29828 4984
rect 29880 4972 29886 5024
rect 29914 4972 29920 5024
rect 29972 5012 29978 5024
rect 30929 5015 30987 5021
rect 30929 5012 30941 5015
rect 29972 4984 30941 5012
rect 29972 4972 29978 4984
rect 30929 4981 30941 4984
rect 30975 4981 30987 5015
rect 30929 4975 30987 4981
rect 32401 5015 32459 5021
rect 32401 4981 32413 5015
rect 32447 5012 32459 5015
rect 33778 5012 33784 5024
rect 32447 4984 33784 5012
rect 32447 4981 32459 4984
rect 32401 4975 32459 4981
rect 33778 4972 33784 4984
rect 33836 4972 33842 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 7926 4808 7932 4820
rect 4304 4780 7512 4808
rect 7887 4780 7932 4808
rect 4304 4768 4310 4780
rect 3421 4743 3479 4749
rect 3421 4709 3433 4743
rect 3467 4740 3479 4743
rect 3602 4740 3608 4752
rect 3467 4712 3608 4740
rect 3467 4709 3479 4712
rect 3421 4703 3479 4709
rect 3602 4700 3608 4712
rect 3660 4740 3666 4752
rect 3878 4740 3884 4752
rect 3660 4712 3884 4740
rect 3660 4700 3666 4712
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 7484 4740 7512 4780
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8352 4780 8401 4808
rect 8352 4768 8358 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 11517 4811 11575 4817
rect 11517 4777 11529 4811
rect 11563 4808 11575 4811
rect 11698 4808 11704 4820
rect 11563 4780 11704 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 21174 4808 21180 4820
rect 13372 4780 20760 4808
rect 21135 4780 21180 4808
rect 9490 4740 9496 4752
rect 7484 4712 9496 4740
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 3973 4675 4031 4681
rect 1995 4644 3924 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 3510 4536 3516 4548
rect 3174 4508 3516 4536
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 3896 4468 3924 4644
rect 3973 4641 3985 4675
rect 4019 4641 4031 4675
rect 3973 4635 4031 4641
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4672 6239 4675
rect 7006 4672 7012 4684
rect 6227 4644 7012 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 3988 4548 4016 4635
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 9766 4672 9772 4684
rect 9679 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4672 9830 4684
rect 10042 4672 10048 4684
rect 9824 4644 10048 4672
rect 9824 4632 9830 4644
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 11977 4675 12035 4681
rect 11977 4672 11989 4675
rect 11756 4644 11989 4672
rect 11756 4632 11762 4644
rect 11977 4641 11989 4644
rect 12023 4672 12035 4675
rect 12250 4672 12256 4684
rect 12023 4644 12256 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8444 4576 8585 4604
rect 8444 4564 8450 4576
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4604 9183 4607
rect 9214 4604 9220 4616
rect 9171 4576 9220 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 13372 4590 13400 4780
rect 13725 4743 13783 4749
rect 13725 4709 13737 4743
rect 13771 4740 13783 4743
rect 13814 4740 13820 4752
rect 13771 4712 13820 4740
rect 13771 4709 13783 4712
rect 13725 4703 13783 4709
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 20732 4740 20760 4780
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 28721 4811 28779 4817
rect 28721 4808 28733 4811
rect 21284 4780 28733 4808
rect 21284 4740 21312 4780
rect 28721 4777 28733 4780
rect 28767 4777 28779 4811
rect 28721 4771 28779 4777
rect 31757 4811 31815 4817
rect 31757 4777 31769 4811
rect 31803 4808 31815 4811
rect 31846 4808 31852 4820
rect 31803 4780 31852 4808
rect 31803 4777 31815 4780
rect 31757 4771 31815 4777
rect 31846 4768 31852 4780
rect 31904 4768 31910 4820
rect 20732 4712 21312 4740
rect 23566 4700 23572 4752
rect 23624 4740 23630 4752
rect 27433 4743 27491 4749
rect 27433 4740 27445 4743
rect 23624 4712 27445 4740
rect 23624 4700 23630 4712
rect 27433 4709 27445 4712
rect 27479 4709 27491 4743
rect 27433 4703 27491 4709
rect 27522 4700 27528 4752
rect 27580 4740 27586 4752
rect 32309 4743 32367 4749
rect 32309 4740 32321 4743
rect 27580 4712 32321 4740
rect 27580 4700 27586 4712
rect 32309 4709 32321 4712
rect 32355 4709 32367 4743
rect 33594 4740 33600 4752
rect 33555 4712 33600 4740
rect 32309 4703 32367 4709
rect 33594 4700 33600 4712
rect 33652 4700 33658 4752
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 16298 4672 16304 4684
rect 15335 4644 16304 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16632 4644 17049 4672
rect 16632 4632 16638 4644
rect 17037 4641 17049 4644
rect 17083 4672 17095 4675
rect 17310 4672 17316 4684
rect 17083 4644 17316 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 18598 4672 18604 4684
rect 17788 4644 18604 4672
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 14608 4576 15025 4604
rect 14608 4564 14614 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 17788 4604 17816 4644
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 18785 4675 18843 4681
rect 18785 4641 18797 4675
rect 18831 4672 18843 4675
rect 19150 4672 19156 4684
rect 18831 4644 19156 4672
rect 18831 4641 18843 4644
rect 18785 4635 18843 4641
rect 19150 4632 19156 4644
rect 19208 4672 19214 4684
rect 21637 4675 21695 4681
rect 21637 4672 21649 4675
rect 19208 4644 21649 4672
rect 19208 4632 19214 4644
rect 21637 4641 21649 4644
rect 21683 4641 21695 4675
rect 29825 4675 29883 4681
rect 29825 4672 29837 4675
rect 21637 4635 21695 4641
rect 23032 4644 29837 4672
rect 17954 4604 17960 4616
rect 16422 4576 17816 4604
rect 17915 4576 17960 4604
rect 15013 4567 15071 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 21542 4604 21548 4616
rect 20838 4576 21548 4604
rect 19429 4567 19487 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 23032 4590 23060 4644
rect 29825 4641 29837 4644
rect 29871 4641 29883 4675
rect 29825 4635 29883 4641
rect 29932 4644 33180 4672
rect 25317 4607 25375 4613
rect 25317 4573 25329 4607
rect 25363 4604 25375 4607
rect 25406 4604 25412 4616
rect 25363 4576 25412 4604
rect 25363 4573 25375 4576
rect 25317 4567 25375 4573
rect 25406 4564 25412 4576
rect 25464 4564 25470 4616
rect 25682 4564 25688 4616
rect 25740 4604 25746 4616
rect 26053 4607 26111 4613
rect 26053 4604 26065 4607
rect 25740 4576 26065 4604
rect 25740 4564 25746 4576
rect 26053 4573 26065 4576
rect 26099 4573 26111 4607
rect 26053 4567 26111 4573
rect 26142 4564 26148 4616
rect 26200 4604 26206 4616
rect 26697 4607 26755 4613
rect 26697 4604 26709 4607
rect 26200 4576 26709 4604
rect 26200 4564 26206 4576
rect 26697 4573 26709 4576
rect 26743 4573 26755 4607
rect 26697 4567 26755 4573
rect 26878 4564 26884 4616
rect 26936 4604 26942 4616
rect 27341 4607 27399 4613
rect 27341 4604 27353 4607
rect 26936 4576 27353 4604
rect 26936 4564 26942 4576
rect 27341 4573 27353 4576
rect 27387 4604 27399 4607
rect 27798 4604 27804 4616
rect 27387 4576 27804 4604
rect 27387 4573 27399 4576
rect 27341 4567 27399 4573
rect 27798 4564 27804 4576
rect 27856 4564 27862 4616
rect 27982 4604 27988 4616
rect 27943 4576 27988 4604
rect 27982 4564 27988 4576
rect 28040 4564 28046 4616
rect 28534 4564 28540 4616
rect 28592 4604 28598 4616
rect 28629 4607 28687 4613
rect 28629 4604 28641 4607
rect 28592 4576 28641 4604
rect 28592 4564 28598 4576
rect 28629 4573 28641 4576
rect 28675 4573 28687 4607
rect 28629 4567 28687 4573
rect 28902 4564 28908 4616
rect 28960 4604 28966 4616
rect 29270 4604 29276 4616
rect 28960 4576 29276 4604
rect 28960 4564 28966 4576
rect 29270 4564 29276 4576
rect 29328 4564 29334 4616
rect 29730 4604 29736 4616
rect 29691 4576 29736 4604
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 3970 4496 3976 4548
rect 4028 4496 4034 4548
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4536 4307 4539
rect 4522 4536 4528 4548
rect 4295 4508 4528 4536
rect 4295 4505 4307 4508
rect 4249 4499 4307 4505
rect 4522 4496 4528 4508
rect 4580 4496 4586 4548
rect 5258 4496 5264 4548
rect 5316 4496 5322 4548
rect 5994 4536 6000 4548
rect 5552 4508 6000 4536
rect 5552 4468 5580 4508
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 6457 4539 6515 4545
rect 6457 4536 6469 4539
rect 6420 4508 6469 4536
rect 6420 4496 6426 4508
rect 6457 4505 6469 4508
rect 6503 4505 6515 4539
rect 10042 4536 10048 4548
rect 6457 4499 6515 4505
rect 6564 4508 6946 4536
rect 10003 4508 10048 4536
rect 3896 4440 5580 4468
rect 5721 4471 5779 4477
rect 5721 4437 5733 4471
rect 5767 4468 5779 4471
rect 5902 4468 5908 4480
rect 5767 4440 5908 4468
rect 5767 4437 5779 4440
rect 5721 4431 5779 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 6564 4468 6592 4508
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 12253 4539 12311 4545
rect 11270 4508 11652 4536
rect 9214 4468 9220 4480
rect 6236 4440 6592 4468
rect 9175 4440 9220 4468
rect 6236 4428 6242 4440
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 11624 4468 11652 4508
rect 12253 4505 12265 4539
rect 12299 4536 12311 4539
rect 12342 4536 12348 4548
rect 12299 4508 12348 4536
rect 12299 4505 12311 4508
rect 12253 4499 12311 4505
rect 12342 4496 12348 4508
rect 12400 4496 12406 4548
rect 13648 4508 14964 4536
rect 13648 4468 13676 4508
rect 11624 4440 13676 4468
rect 14461 4471 14519 4477
rect 14461 4437 14473 4471
rect 14507 4468 14519 4471
rect 14826 4468 14832 4480
rect 14507 4440 14832 4468
rect 14507 4437 14519 4440
rect 14461 4431 14519 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 14936 4468 14964 4508
rect 17126 4496 17132 4548
rect 17184 4536 17190 4548
rect 18782 4536 18788 4548
rect 17184 4508 18788 4536
rect 17184 4496 17190 4508
rect 18782 4496 18788 4508
rect 18840 4496 18846 4548
rect 18966 4496 18972 4548
rect 19024 4536 19030 4548
rect 19705 4539 19763 4545
rect 19705 4536 19717 4539
rect 19024 4508 19717 4536
rect 19024 4496 19030 4508
rect 19705 4505 19717 4508
rect 19751 4536 19763 4539
rect 19978 4536 19984 4548
rect 19751 4508 19984 4536
rect 19751 4505 19763 4508
rect 19705 4499 19763 4505
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 20990 4496 20996 4548
rect 21048 4536 21054 4548
rect 21913 4539 21971 4545
rect 21913 4536 21925 4539
rect 21048 4508 21925 4536
rect 21048 4496 21054 4508
rect 21913 4505 21925 4508
rect 21959 4536 21971 4539
rect 22002 4536 22008 4548
rect 21959 4508 22008 4536
rect 21959 4505 21971 4508
rect 21913 4499 21971 4505
rect 22002 4496 22008 4508
rect 22060 4496 22066 4548
rect 24026 4536 24032 4548
rect 23400 4508 24032 4536
rect 18046 4468 18052 4480
rect 14936 4440 18052 4468
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 21082 4468 21088 4480
rect 19392 4440 21088 4468
rect 19392 4428 19398 4440
rect 21082 4428 21088 4440
rect 21140 4428 21146 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 23400 4477 23428 4508
rect 24026 4496 24032 4508
rect 24084 4496 24090 4548
rect 24670 4536 24676 4548
rect 24631 4508 24676 4536
rect 24670 4496 24676 4508
rect 24728 4496 24734 4548
rect 24765 4539 24823 4545
rect 24765 4505 24777 4539
rect 24811 4505 24823 4539
rect 26510 4536 26516 4548
rect 24765 4499 24823 4505
rect 25424 4508 26516 4536
rect 23385 4471 23443 4477
rect 23385 4468 23397 4471
rect 22152 4440 23397 4468
rect 22152 4428 22158 4440
rect 23385 4437 23397 4440
rect 23431 4437 23443 4471
rect 23842 4468 23848 4480
rect 23803 4440 23848 4468
rect 23385 4431 23443 4437
rect 23842 4428 23848 4440
rect 23900 4428 23906 4480
rect 24780 4468 24808 4499
rect 25424 4468 25452 4508
rect 26510 4496 26516 4508
rect 26568 4496 26574 4548
rect 27522 4536 27528 4548
rect 26620 4508 27528 4536
rect 26142 4468 26148 4480
rect 24780 4440 25452 4468
rect 26103 4440 26148 4468
rect 26142 4428 26148 4440
rect 26200 4428 26206 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 26620 4468 26648 4508
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
rect 27632 4508 28212 4536
rect 26786 4468 26792 4480
rect 26292 4440 26648 4468
rect 26747 4440 26792 4468
rect 26292 4428 26298 4440
rect 26786 4428 26792 4440
rect 26844 4428 26850 4480
rect 26878 4428 26884 4480
rect 26936 4468 26942 4480
rect 27632 4468 27660 4508
rect 28074 4468 28080 4480
rect 26936 4440 27660 4468
rect 28035 4440 28080 4468
rect 26936 4428 26942 4440
rect 28074 4428 28080 4440
rect 28132 4428 28138 4480
rect 28184 4468 28212 4508
rect 28258 4496 28264 4548
rect 28316 4536 28322 4548
rect 29932 4536 29960 4644
rect 30377 4607 30435 4613
rect 30377 4573 30389 4607
rect 30423 4604 30435 4607
rect 30742 4604 30748 4616
rect 30423 4576 30748 4604
rect 30423 4573 30435 4576
rect 30377 4567 30435 4573
rect 30742 4564 30748 4576
rect 30800 4564 30806 4616
rect 31021 4607 31079 4613
rect 31021 4573 31033 4607
rect 31067 4604 31079 4607
rect 31202 4604 31208 4616
rect 31067 4576 31208 4604
rect 31067 4573 31079 4576
rect 31021 4567 31079 4573
rect 31202 4564 31208 4576
rect 31260 4564 31266 4616
rect 31662 4604 31668 4616
rect 31623 4576 31668 4604
rect 31662 4564 31668 4576
rect 31720 4564 31726 4616
rect 32490 4604 32496 4616
rect 32451 4576 32496 4604
rect 32490 4564 32496 4576
rect 32548 4564 32554 4616
rect 33152 4613 33180 4644
rect 33137 4607 33195 4613
rect 33137 4573 33149 4607
rect 33183 4573 33195 4607
rect 33778 4604 33784 4616
rect 33739 4576 33784 4604
rect 33137 4567 33195 4573
rect 33778 4564 33784 4576
rect 33836 4564 33842 4616
rect 38010 4604 38016 4616
rect 37971 4576 38016 4604
rect 38010 4564 38016 4576
rect 38068 4564 38074 4616
rect 31110 4536 31116 4548
rect 28316 4508 29960 4536
rect 31071 4508 31116 4536
rect 28316 4496 28322 4508
rect 31110 4496 31116 4508
rect 31168 4496 31174 4548
rect 29914 4468 29920 4480
rect 28184 4440 29920 4468
rect 29914 4428 29920 4440
rect 29972 4428 29978 4480
rect 30466 4468 30472 4480
rect 30427 4440 30472 4468
rect 30466 4428 30472 4440
rect 30524 4428 30530 4480
rect 30650 4428 30656 4480
rect 30708 4468 30714 4480
rect 32953 4471 33011 4477
rect 32953 4468 32965 4471
rect 30708 4440 32965 4468
rect 30708 4428 30714 4440
rect 32953 4437 32965 4440
rect 32999 4437 33011 4471
rect 38194 4468 38200 4480
rect 38155 4440 38200 4468
rect 32953 4431 33011 4437
rect 38194 4428 38200 4440
rect 38252 4428 38258 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 9214 4264 9220 4276
rect 4856 4236 9220 4264
rect 4856 4224 4862 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 26142 4264 26148 4276
rect 9324 4236 26148 4264
rect 4246 4196 4252 4208
rect 3174 4168 4252 4196
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 4522 4196 4528 4208
rect 4483 4168 4528 4196
rect 4522 4156 4528 4168
rect 4580 4156 4586 4208
rect 5810 4196 5816 4208
rect 5750 4168 5816 4196
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 5902 4156 5908 4208
rect 5960 4196 5966 4208
rect 7098 4196 7104 4208
rect 5960 4168 7104 4196
rect 5960 4156 5966 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 9324 4196 9352 4236
rect 26142 4224 26148 4236
rect 26200 4224 26206 4276
rect 26234 4224 26240 4276
rect 26292 4264 26298 4276
rect 28994 4264 29000 4276
rect 26292 4236 29000 4264
rect 26292 4224 26298 4236
rect 28994 4224 29000 4236
rect 29052 4224 29058 4276
rect 29454 4224 29460 4276
rect 29512 4264 29518 4276
rect 33597 4267 33655 4273
rect 33597 4264 33609 4267
rect 29512 4236 33609 4264
rect 29512 4224 29518 4236
rect 33597 4233 33609 4236
rect 33643 4233 33655 4267
rect 33597 4227 33655 4233
rect 9766 4196 9772 4208
rect 8050 4168 9352 4196
rect 9416 4168 9772 4196
rect 9416 4137 9444 4168
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 10962 4196 10968 4208
rect 10902 4168 10968 4196
rect 10962 4156 10968 4168
rect 11020 4156 11026 4208
rect 13262 4196 13268 4208
rect 13202 4168 13268 4196
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 14829 4199 14887 4205
rect 14829 4165 14841 4199
rect 14875 4196 14887 4199
rect 14918 4196 14924 4208
rect 14875 4168 14924 4196
rect 14875 4165 14887 4168
rect 14829 4159 14887 4165
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 16390 4196 16396 4208
rect 16054 4168 16396 4196
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 17126 4196 17132 4208
rect 17087 4168 17132 4196
rect 17126 4156 17132 4168
rect 17184 4156 17190 4208
rect 19334 4196 19340 4208
rect 18354 4168 19340 4196
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 19426 4156 19432 4208
rect 19484 4196 19490 4208
rect 19484 4168 19529 4196
rect 19484 4156 19490 4168
rect 20162 4156 20168 4208
rect 20220 4156 20226 4208
rect 22094 4196 22100 4208
rect 20824 4168 22100 4196
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4097 9459 4131
rect 11698 4128 11704 4140
rect 11659 4100 11704 4128
rect 9401 4091 9459 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 1670 4060 1676 4072
rect 1631 4032 1676 4060
rect 1670 4020 1676 4032
rect 1728 4020 1734 4072
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4060 2007 4063
rect 3418 4060 3424 4072
rect 1995 4032 3424 4060
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4120 4032 4261 4060
rect 4120 4020 4126 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 6546 4060 6552 4072
rect 4249 4023 4307 4029
rect 4356 4032 5580 4060
rect 6507 4032 6552 4060
rect 4356 3992 4384 4032
rect 3712 3964 4384 3992
rect 5552 3992 5580 4032
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6656 4032 6837 4060
rect 6656 3992 6684 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 8260 4032 9689 4060
rect 8260 4020 8266 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 11330 4060 11336 4072
rect 10192 4032 11336 4060
rect 10192 4020 10198 4032
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11974 4060 11980 4072
rect 11440 4032 11980 4060
rect 5552 3964 6684 3992
rect 8220 3964 9536 3992
rect 3712 3936 3740 3964
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 3694 3924 3700 3936
rect 3467 3896 3700 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4890 3924 4896 3936
rect 3936 3896 4896 3924
rect 3936 3884 3942 3896
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 8220 3924 8248 3964
rect 6043 3896 8248 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 9508 3924 9536 3964
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11440 3992 11468 4032
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 13538 4060 13544 4072
rect 12676 4032 13544 4060
rect 12676 4020 12682 4032
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 13722 4060 13728 4072
rect 13683 4032 13728 4060
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 16850 4060 16856 4072
rect 14660 4032 16712 4060
rect 16811 4032 16856 4060
rect 14660 3992 14688 4032
rect 11112 3964 11468 3992
rect 13004 3964 14688 3992
rect 16684 3992 16712 4032
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 18966 4060 18972 4072
rect 16960 4032 18972 4060
rect 16960 3992 16988 4032
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 19058 4020 19064 4072
rect 19116 4060 19122 4072
rect 20824 4060 20852 4168
rect 22094 4156 22100 4168
rect 22152 4156 22158 4208
rect 22465 4199 22523 4205
rect 22465 4165 22477 4199
rect 22511 4196 22523 4199
rect 24029 4199 24087 4205
rect 22511 4168 23244 4196
rect 22511 4165 22523 4168
rect 22465 4159 22523 4165
rect 21358 4128 21364 4140
rect 20916 4100 21364 4128
rect 20916 4069 20944 4100
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 19116 4032 20852 4060
rect 20901 4063 20959 4069
rect 19116 4020 19122 4032
rect 20901 4029 20913 4063
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 22373 4063 22431 4069
rect 22373 4029 22385 4063
rect 22419 4060 22431 4063
rect 23014 4060 23020 4072
rect 22419 4032 23020 4060
rect 22419 4029 22431 4032
rect 22373 4023 22431 4029
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 22646 3992 22652 4004
rect 16684 3964 16988 3992
rect 18156 3964 18736 3992
rect 11112 3952 11118 3964
rect 10042 3924 10048 3936
rect 8352 3896 8397 3924
rect 9508 3896 10048 3924
rect 8352 3884 8358 3896
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 13004 3924 13032 3964
rect 11195 3896 13032 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 13136 3896 16313 3924
rect 13136 3884 13142 3896
rect 16301 3893 16313 3896
rect 16347 3924 16359 3927
rect 18156 3924 18184 3964
rect 18598 3924 18604 3936
rect 16347 3896 18184 3924
rect 18559 3896 18604 3924
rect 16347 3893 16359 3896
rect 16301 3887 16359 3893
rect 18598 3884 18604 3896
rect 18656 3884 18662 3936
rect 18708 3924 18736 3964
rect 21284 3964 22652 3992
rect 20438 3924 20444 3936
rect 18708 3896 20444 3924
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 21284 3924 21312 3964
rect 22646 3952 22652 3964
rect 22704 3952 22710 4004
rect 23216 3992 23244 4168
rect 24029 4165 24041 4199
rect 24075 4196 24087 4199
rect 26786 4196 26792 4208
rect 24075 4168 26792 4196
rect 24075 4165 24087 4168
rect 24029 4159 24087 4165
rect 26786 4156 26792 4168
rect 26844 4156 26850 4208
rect 27430 4196 27436 4208
rect 26896 4168 27436 4196
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24946 4128 24952 4140
rect 24627 4100 24952 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 25038 4088 25044 4140
rect 25096 4128 25102 4140
rect 25096 4100 25141 4128
rect 25096 4088 25102 4100
rect 25590 4088 25596 4140
rect 25648 4128 25654 4140
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25648 4100 25789 4128
rect 25648 4088 25654 4100
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 25777 4091 25835 4097
rect 26421 4131 26479 4137
rect 26421 4097 26433 4131
rect 26467 4128 26479 4131
rect 26896 4128 26924 4168
rect 27430 4156 27436 4168
rect 27488 4196 27494 4208
rect 28534 4196 28540 4208
rect 27488 4168 28540 4196
rect 27488 4156 27494 4168
rect 28534 4156 28540 4168
rect 28592 4156 28598 4208
rect 31662 4196 31668 4208
rect 29196 4168 31668 4196
rect 27154 4128 27160 4140
rect 26467 4100 26924 4128
rect 27115 4100 27160 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 27798 4128 27804 4140
rect 27759 4100 27804 4128
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 27982 4088 27988 4140
rect 28040 4128 28046 4140
rect 28445 4131 28503 4137
rect 28445 4128 28457 4131
rect 28040 4100 28457 4128
rect 28040 4088 28046 4100
rect 28445 4097 28457 4100
rect 28491 4128 28503 4131
rect 28902 4128 28908 4140
rect 28491 4100 28908 4128
rect 28491 4097 28503 4100
rect 28445 4091 28503 4097
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 29086 4128 29092 4140
rect 29047 4100 29092 4128
rect 29086 4088 29092 4100
rect 29144 4088 29150 4140
rect 23382 4060 23388 4072
rect 23343 4032 23388 4060
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 23934 4060 23940 4072
rect 23895 4032 23940 4060
rect 23934 4020 23940 4032
rect 23992 4020 23998 4072
rect 27893 4063 27951 4069
rect 27893 4060 27905 4063
rect 24044 4032 27905 4060
rect 24044 3992 24072 4032
rect 27893 4029 27905 4032
rect 27939 4029 27951 4063
rect 27893 4023 27951 4029
rect 28350 4020 28356 4072
rect 28408 4060 28414 4072
rect 29196 4060 29224 4168
rect 31662 4156 31668 4168
rect 31720 4156 31726 4208
rect 32876 4168 33088 4196
rect 29270 4088 29276 4140
rect 29328 4128 29334 4140
rect 29733 4131 29791 4137
rect 29733 4128 29745 4131
rect 29328 4100 29745 4128
rect 29328 4088 29334 4100
rect 29733 4097 29745 4100
rect 29779 4097 29791 4131
rect 29733 4091 29791 4097
rect 30377 4131 30435 4137
rect 30377 4097 30389 4131
rect 30423 4097 30435 4131
rect 30377 4091 30435 4097
rect 30469 4131 30527 4137
rect 30469 4097 30481 4131
rect 30515 4128 30527 4131
rect 30558 4128 30564 4140
rect 30515 4100 30564 4128
rect 30515 4097 30527 4100
rect 30469 4091 30527 4097
rect 28408 4032 29224 4060
rect 28408 4020 28414 4032
rect 29638 4020 29644 4072
rect 29696 4060 29702 4072
rect 30392 4060 30420 4091
rect 30558 4088 30564 4100
rect 30616 4088 30622 4140
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 31021 4131 31079 4137
rect 31021 4128 31033 4131
rect 30800 4100 31033 4128
rect 30800 4088 30806 4100
rect 31021 4097 31033 4100
rect 31067 4128 31079 4131
rect 31570 4128 31576 4140
rect 31067 4100 31576 4128
rect 31067 4097 31079 4100
rect 31021 4091 31079 4097
rect 31570 4088 31576 4100
rect 31628 4088 31634 4140
rect 32309 4131 32367 4137
rect 32309 4097 32321 4131
rect 32355 4128 32367 4131
rect 32398 4128 32404 4140
rect 32355 4100 32404 4128
rect 32355 4097 32367 4100
rect 32309 4091 32367 4097
rect 32398 4088 32404 4100
rect 32456 4088 32462 4140
rect 29696 4032 30420 4060
rect 29696 4020 29702 4032
rect 31110 4020 31116 4072
rect 31168 4060 31174 4072
rect 32876 4060 32904 4168
rect 32953 4131 33011 4137
rect 32953 4097 32965 4131
rect 32999 4097 33011 4131
rect 33060 4128 33088 4168
rect 33781 4131 33839 4137
rect 33781 4128 33793 4131
rect 33060 4100 33793 4128
rect 32953 4091 33011 4097
rect 33781 4097 33793 4100
rect 33827 4097 33839 4131
rect 33781 4091 33839 4097
rect 34241 4131 34299 4137
rect 34241 4097 34253 4131
rect 34287 4097 34299 4131
rect 38286 4128 38292 4140
rect 38247 4100 38292 4128
rect 34241 4091 34299 4097
rect 31168 4032 32904 4060
rect 31168 4020 31174 4032
rect 23216 3964 24072 3992
rect 24854 3952 24860 4004
rect 24912 3992 24918 4004
rect 25133 3995 25191 4001
rect 25133 3992 25145 3995
rect 24912 3964 25145 3992
rect 24912 3952 24918 3964
rect 25133 3961 25145 3964
rect 25179 3961 25191 3995
rect 25133 3955 25191 3961
rect 25314 3952 25320 4004
rect 25372 3992 25378 4004
rect 29181 3995 29239 4001
rect 29181 3992 29193 3995
rect 25372 3964 29193 3992
rect 25372 3952 25378 3964
rect 29181 3961 29193 3964
rect 29227 3961 29239 3995
rect 29181 3955 29239 3961
rect 29270 3952 29276 4004
rect 29328 3992 29334 4004
rect 32401 3995 32459 4001
rect 32401 3992 32413 3995
rect 29328 3964 32413 3992
rect 29328 3952 29334 3964
rect 32401 3961 32413 3964
rect 32447 3961 32459 3995
rect 32968 3992 32996 4091
rect 33042 4020 33048 4072
rect 33100 4060 33106 4072
rect 34256 4060 34284 4091
rect 38286 4088 38292 4100
rect 38344 4088 38350 4140
rect 33100 4032 34284 4060
rect 33100 4020 33106 4032
rect 32401 3955 32459 3961
rect 32508 3964 32996 3992
rect 20588 3896 21312 3924
rect 20588 3884 20594 3896
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 22370 3924 22376 3936
rect 21416 3896 22376 3924
rect 21416 3884 21422 3896
rect 22370 3884 22376 3896
rect 22428 3884 22434 3936
rect 22554 3884 22560 3936
rect 22612 3924 22618 3936
rect 23934 3924 23940 3936
rect 22612 3896 23940 3924
rect 22612 3884 22618 3896
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 25222 3884 25228 3936
rect 25280 3924 25286 3936
rect 25869 3927 25927 3933
rect 25869 3924 25881 3927
rect 25280 3896 25881 3924
rect 25280 3884 25286 3896
rect 25869 3893 25881 3896
rect 25915 3893 25927 3927
rect 26510 3924 26516 3936
rect 26471 3896 26516 3924
rect 25869 3887 25927 3893
rect 26510 3884 26516 3896
rect 26568 3884 26574 3936
rect 26786 3884 26792 3936
rect 26844 3924 26850 3936
rect 27249 3927 27307 3933
rect 27249 3924 27261 3927
rect 26844 3896 27261 3924
rect 26844 3884 26850 3896
rect 27249 3893 27261 3896
rect 27295 3893 27307 3927
rect 27249 3887 27307 3893
rect 27614 3884 27620 3936
rect 27672 3924 27678 3936
rect 28350 3924 28356 3936
rect 27672 3896 28356 3924
rect 27672 3884 27678 3896
rect 28350 3884 28356 3896
rect 28408 3884 28414 3936
rect 28534 3924 28540 3936
rect 28495 3896 28540 3924
rect 28534 3884 28540 3896
rect 28592 3884 28598 3936
rect 29362 3884 29368 3936
rect 29420 3924 29426 3936
rect 29825 3927 29883 3933
rect 29825 3924 29837 3927
rect 29420 3896 29837 3924
rect 29420 3884 29426 3896
rect 29825 3893 29837 3896
rect 29871 3893 29883 3927
rect 29825 3887 29883 3893
rect 30558 3884 30564 3936
rect 30616 3924 30622 3936
rect 31113 3927 31171 3933
rect 31113 3924 31125 3927
rect 30616 3896 31125 3924
rect 30616 3884 30622 3896
rect 31113 3893 31125 3896
rect 31159 3893 31171 3927
rect 31113 3887 31171 3893
rect 31294 3884 31300 3936
rect 31352 3924 31358 3936
rect 32508 3924 32536 3964
rect 35802 3952 35808 4004
rect 35860 3992 35866 4004
rect 38105 3995 38163 4001
rect 38105 3992 38117 3995
rect 35860 3964 38117 3992
rect 35860 3952 35866 3964
rect 38105 3961 38117 3964
rect 38151 3961 38163 3995
rect 38105 3955 38163 3961
rect 33042 3924 33048 3936
rect 31352 3896 32536 3924
rect 33003 3896 33048 3924
rect 31352 3884 31358 3896
rect 33042 3884 33048 3896
rect 33100 3884 33106 3936
rect 34333 3927 34391 3933
rect 34333 3893 34345 3927
rect 34379 3924 34391 3927
rect 35710 3924 35716 3936
rect 34379 3896 35716 3924
rect 34379 3893 34391 3896
rect 34333 3887 34391 3893
rect 35710 3884 35716 3896
rect 35768 3884 35774 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3200 3692 3433 3720
rect 3200 3680 3206 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 4982 3720 4988 3732
rect 3421 3683 3479 3689
rect 3988 3692 4988 3720
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2038 3584 2044 3596
rect 1995 3556 2044 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 3988 3525 4016 3692
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 6365 3723 6423 3729
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 6822 3720 6828 3732
rect 6411 3692 6828 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 9398 3720 9404 3732
rect 7156 3692 9404 3720
rect 7156 3680 7162 3692
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 11882 3720 11888 3732
rect 9508 3692 11888 3720
rect 8478 3612 8484 3664
rect 8536 3652 8542 3664
rect 9508 3652 9536 3692
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12802 3720 12808 3732
rect 12084 3692 12808 3720
rect 8536 3624 9536 3652
rect 8536 3612 8542 3624
rect 11054 3612 11060 3664
rect 11112 3652 11118 3664
rect 12084 3652 12112 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 20990 3720 20996 3732
rect 12952 3692 18092 3720
rect 12952 3680 12958 3692
rect 11112 3624 12112 3652
rect 11112 3612 11118 3624
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 17589 3655 17647 3661
rect 13780 3624 15976 3652
rect 13780 3612 13786 3624
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3584 4675 3587
rect 6546 3584 6552 3596
rect 4663 3556 6552 3584
rect 4663 3553 4675 3556
rect 4617 3547 4675 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 9766 3584 9772 3596
rect 6871 3556 9772 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10778 3584 10784 3596
rect 10091 3556 10784 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11977 3587 12035 3593
rect 11977 3553 11989 3587
rect 12023 3584 12035 3587
rect 14550 3584 14556 3596
rect 12023 3556 14556 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 14550 3544 14556 3556
rect 14608 3584 14614 3596
rect 15197 3587 15255 3593
rect 15197 3584 15209 3587
rect 14608 3556 15209 3584
rect 14608 3544 14614 3556
rect 15197 3553 15209 3556
rect 15243 3584 15255 3587
rect 15841 3587 15899 3593
rect 15841 3584 15853 3587
rect 15243 3556 15853 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 15841 3553 15853 3556
rect 15887 3553 15899 3587
rect 15948 3584 15976 3624
rect 17589 3621 17601 3655
rect 17635 3652 17647 3655
rect 17770 3652 17776 3664
rect 17635 3624 17776 3652
rect 17635 3621 17647 3624
rect 17589 3615 17647 3621
rect 17770 3612 17776 3624
rect 17828 3612 17834 3664
rect 16574 3584 16580 3596
rect 15948 3556 16580 3584
rect 15841 3547 15899 3553
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 18064 3593 18092 3692
rect 19076 3692 20996 3720
rect 18049 3587 18107 3593
rect 16724 3556 17632 3584
rect 16724 3544 16730 3556
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 9309 3519 9367 3525
rect 6026 3488 6868 3516
rect 3973 3479 4031 3485
rect 6840 3460 6868 3488
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14734 3516 14740 3528
rect 14507 3488 14740 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 4798 3448 4804 3460
rect 3174 3420 4804 3448
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 4890 3408 4896 3460
rect 4948 3448 4954 3460
rect 4948 3420 4993 3448
rect 4948 3408 4954 3420
rect 6822 3408 6828 3460
rect 6880 3408 6886 3460
rect 7006 3408 7012 3460
rect 7064 3448 7070 3460
rect 7101 3451 7159 3457
rect 7101 3448 7113 3451
rect 7064 3420 7113 3448
rect 7064 3408 7070 3420
rect 7101 3417 7113 3420
rect 7147 3417 7159 3451
rect 7101 3411 7159 3417
rect 7190 3408 7196 3460
rect 7248 3448 7254 3460
rect 7248 3420 7590 3448
rect 7248 3408 7254 3420
rect 4065 3383 4123 3389
rect 4065 3349 4077 3383
rect 4111 3380 4123 3383
rect 5258 3380 5264 3392
rect 4111 3352 5264 3380
rect 4111 3349 4123 3352
rect 4065 3343 4123 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 8478 3380 8484 3392
rect 5592 3352 8484 3380
rect 5592 3340 5598 3352
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9122 3380 9128 3392
rect 8628 3352 8673 3380
rect 9083 3352 9128 3380
rect 8628 3340 8634 3352
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9324 3380 9352 3479
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 17604 3516 17632 3556
rect 18049 3553 18061 3587
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 17770 3516 17776 3528
rect 17604 3488 17776 3516
rect 17770 3476 17776 3488
rect 17828 3516 17834 3528
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 17828 3488 18337 3516
rect 17828 3476 17834 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 10134 3448 10140 3460
rect 9456 3420 10140 3448
rect 9456 3408 9462 3420
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 12158 3448 12164 3460
rect 11270 3420 12164 3448
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 12253 3451 12311 3457
rect 12253 3417 12265 3451
rect 12299 3448 12311 3451
rect 12526 3448 12532 3460
rect 12299 3420 12532 3448
rect 12299 3417 12311 3420
rect 12253 3411 12311 3417
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 13538 3448 13544 3460
rect 13478 3420 13544 3448
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 16114 3448 16120 3460
rect 13648 3420 15976 3448
rect 16075 3420 16120 3448
rect 10870 3380 10876 3392
rect 9324 3352 10876 3380
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 11517 3383 11575 3389
rect 11517 3349 11529 3383
rect 11563 3380 11575 3383
rect 13648 3380 13676 3420
rect 11563 3352 13676 3380
rect 11563 3349 11575 3352
rect 11517 3343 11575 3349
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 15948 3380 15976 3420
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 17954 3448 17960 3460
rect 17342 3420 17960 3448
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 19076 3448 19104 3692
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 28534 3720 28540 3732
rect 21100 3692 28540 3720
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19429 3587 19487 3593
rect 19429 3584 19441 3587
rect 19208 3556 19441 3584
rect 19208 3544 19214 3556
rect 19429 3553 19441 3556
rect 19475 3553 19487 3587
rect 19429 3547 19487 3553
rect 21100 3516 21128 3692
rect 28534 3680 28540 3692
rect 28592 3680 28598 3732
rect 28718 3680 28724 3732
rect 28776 3720 28782 3732
rect 29638 3720 29644 3732
rect 28776 3692 29644 3720
rect 28776 3680 28782 3692
rect 29638 3680 29644 3692
rect 29696 3680 29702 3732
rect 29822 3720 29828 3732
rect 29783 3692 29828 3720
rect 29822 3680 29828 3692
rect 29880 3680 29886 3732
rect 30374 3680 30380 3732
rect 30432 3720 30438 3732
rect 31757 3723 31815 3729
rect 31757 3720 31769 3723
rect 30432 3692 31769 3720
rect 30432 3680 30438 3692
rect 31757 3689 31769 3692
rect 31803 3689 31815 3723
rect 36722 3720 36728 3732
rect 36683 3692 36728 3720
rect 31757 3683 31815 3689
rect 36722 3680 36728 3692
rect 36780 3680 36786 3732
rect 21177 3655 21235 3661
rect 21177 3621 21189 3655
rect 21223 3652 21235 3655
rect 21266 3652 21272 3664
rect 21223 3624 21272 3652
rect 21223 3621 21235 3624
rect 21177 3615 21235 3621
rect 21266 3612 21272 3624
rect 21324 3612 21330 3664
rect 24946 3652 24952 3664
rect 22066 3624 24952 3652
rect 22066 3584 22094 3624
rect 24946 3612 24952 3624
rect 25004 3612 25010 3664
rect 25682 3612 25688 3664
rect 25740 3652 25746 3664
rect 29270 3652 29276 3664
rect 25740 3624 29276 3652
rect 25740 3612 25746 3624
rect 29270 3612 29276 3624
rect 29328 3612 29334 3664
rect 30650 3612 30656 3664
rect 30708 3652 30714 3664
rect 32309 3655 32367 3661
rect 32309 3652 32321 3655
rect 30708 3624 32321 3652
rect 30708 3612 30714 3624
rect 32309 3621 32321 3624
rect 32355 3621 32367 3655
rect 32309 3615 32367 3621
rect 21192 3556 22094 3584
rect 22833 3587 22891 3593
rect 21192 3528 21220 3556
rect 22833 3553 22845 3587
rect 22879 3584 22891 3587
rect 23842 3584 23848 3596
rect 22879 3556 23848 3584
rect 22879 3553 22891 3556
rect 22833 3547 22891 3553
rect 23842 3544 23848 3556
rect 23900 3544 23906 3596
rect 23934 3544 23940 3596
rect 23992 3584 23998 3596
rect 28534 3584 28540 3596
rect 23992 3556 28540 3584
rect 23992 3544 23998 3556
rect 28534 3544 28540 3556
rect 28592 3544 28598 3596
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 30469 3587 30527 3593
rect 30469 3584 30481 3587
rect 28960 3556 30481 3584
rect 28960 3544 28966 3556
rect 30469 3553 30481 3556
rect 30515 3553 30527 3587
rect 30760 3584 31156 3596
rect 32766 3584 32772 3596
rect 30469 3547 30527 3553
rect 30576 3568 32772 3584
rect 30576 3556 30788 3568
rect 31128 3556 32772 3568
rect 20838 3488 21128 3516
rect 21174 3476 21180 3528
rect 21232 3476 21238 3528
rect 21729 3519 21787 3525
rect 21729 3485 21741 3519
rect 21775 3516 21787 3519
rect 21775 3488 22094 3516
rect 21775 3485 21787 3488
rect 21729 3479 21787 3485
rect 18064 3420 19104 3448
rect 18064 3380 18092 3420
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 19705 3451 19763 3457
rect 19705 3448 19717 3451
rect 19484 3420 19717 3448
rect 19484 3408 19490 3420
rect 19705 3417 19717 3420
rect 19751 3448 19763 3451
rect 19978 3448 19984 3460
rect 19751 3420 19984 3448
rect 19751 3417 19763 3420
rect 19705 3411 19763 3417
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 13780 3352 13825 3380
rect 15948 3352 18092 3380
rect 13780 3340 13786 3352
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 21913 3383 21971 3389
rect 21913 3380 21925 3383
rect 18196 3352 21925 3380
rect 18196 3340 18202 3352
rect 21913 3349 21925 3352
rect 21959 3349 21971 3383
rect 22066 3380 22094 3488
rect 24486 3476 24492 3528
rect 24544 3476 24550 3528
rect 26142 3516 26148 3528
rect 25516 3488 26148 3516
rect 22925 3451 22983 3457
rect 22925 3417 22937 3451
rect 22971 3448 22983 3451
rect 23290 3448 23296 3460
rect 22971 3420 23296 3448
rect 22971 3417 22983 3420
rect 22925 3411 22983 3417
rect 23290 3408 23296 3420
rect 23348 3408 23354 3460
rect 23477 3451 23535 3457
rect 23477 3417 23489 3451
rect 23523 3448 23535 3451
rect 24504 3448 24532 3476
rect 24673 3451 24731 3457
rect 24673 3448 24685 3451
rect 23523 3420 24440 3448
rect 24504 3420 24685 3448
rect 23523 3417 23535 3420
rect 23477 3411 23535 3417
rect 24302 3380 24308 3392
rect 22066 3352 24308 3380
rect 21913 3343 21971 3349
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 24412 3380 24440 3420
rect 24673 3417 24685 3420
rect 24719 3417 24731 3451
rect 24673 3411 24731 3417
rect 24762 3408 24768 3460
rect 24820 3448 24826 3460
rect 24820 3420 24865 3448
rect 24820 3408 24826 3420
rect 25516 3380 25544 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26326 3516 26332 3528
rect 26287 3488 26332 3516
rect 26326 3476 26332 3488
rect 26384 3476 26390 3528
rect 26418 3476 26424 3528
rect 26476 3516 26482 3528
rect 26789 3519 26847 3525
rect 26789 3516 26801 3519
rect 26476 3488 26801 3516
rect 26476 3476 26482 3488
rect 26789 3485 26801 3488
rect 26835 3485 26847 3519
rect 26789 3479 26847 3485
rect 26878 3476 26884 3528
rect 26936 3516 26942 3528
rect 27893 3519 27951 3525
rect 27893 3516 27905 3519
rect 26936 3488 27905 3516
rect 26936 3476 26942 3488
rect 27893 3485 27905 3488
rect 27939 3485 27951 3519
rect 27893 3479 27951 3485
rect 28169 3519 28227 3525
rect 28169 3485 28181 3519
rect 28215 3516 28227 3519
rect 28258 3516 28264 3528
rect 28215 3488 28264 3516
rect 28215 3485 28227 3488
rect 28169 3479 28227 3485
rect 28258 3476 28264 3488
rect 28316 3476 28322 3528
rect 28442 3476 28448 3528
rect 28500 3516 28506 3528
rect 28629 3519 28687 3525
rect 28629 3516 28641 3519
rect 28500 3488 28641 3516
rect 28500 3476 28506 3488
rect 28629 3485 28641 3488
rect 28675 3516 28687 3519
rect 28718 3516 28724 3528
rect 28675 3488 28724 3516
rect 28675 3485 28687 3488
rect 28629 3479 28687 3485
rect 28718 3476 28724 3488
rect 28776 3476 28782 3528
rect 29086 3476 29092 3528
rect 29144 3516 29150 3528
rect 29733 3519 29791 3525
rect 29733 3516 29745 3519
rect 29144 3488 29745 3516
rect 29144 3476 29150 3488
rect 29733 3485 29745 3488
rect 29779 3516 29791 3519
rect 30377 3519 30435 3525
rect 30377 3516 30389 3519
rect 29779 3488 30389 3516
rect 29779 3485 29791 3488
rect 29733 3479 29791 3485
rect 30377 3485 30389 3488
rect 30423 3516 30435 3519
rect 30576 3516 30604 3556
rect 32766 3544 32772 3556
rect 32824 3544 32830 3596
rect 30423 3488 30604 3516
rect 31021 3519 31079 3525
rect 30423 3485 30435 3488
rect 30377 3479 30435 3485
rect 31021 3485 31033 3519
rect 31067 3516 31079 3519
rect 31202 3516 31208 3528
rect 31067 3488 31208 3516
rect 31067 3485 31079 3488
rect 31021 3479 31079 3485
rect 31202 3476 31208 3488
rect 31260 3476 31266 3528
rect 31386 3476 31392 3528
rect 31444 3516 31450 3528
rect 31665 3519 31723 3525
rect 31665 3516 31677 3519
rect 31444 3488 31677 3516
rect 31444 3476 31450 3488
rect 31665 3485 31677 3488
rect 31711 3485 31723 3519
rect 32490 3516 32496 3528
rect 32451 3488 32496 3516
rect 31665 3479 31723 3485
rect 32490 3476 32496 3488
rect 32548 3476 32554 3528
rect 32582 3476 32588 3528
rect 32640 3516 32646 3528
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 32640 3488 32965 3516
rect 32640 3476 32646 3488
rect 32953 3485 32965 3488
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 35069 3519 35127 3525
rect 35069 3516 35081 3519
rect 34756 3488 35081 3516
rect 34756 3476 34762 3488
rect 35069 3485 35081 3488
rect 35115 3485 35127 3519
rect 35710 3516 35716 3528
rect 35671 3488 35716 3516
rect 35069 3479 35127 3485
rect 35710 3476 35716 3488
rect 35768 3476 35774 3528
rect 36909 3519 36967 3525
rect 36909 3485 36921 3519
rect 36955 3516 36967 3519
rect 37366 3516 37372 3528
rect 36955 3488 37372 3516
rect 36955 3485 36967 3488
rect 36909 3479 36967 3485
rect 37366 3476 37372 3488
rect 37424 3476 37430 3528
rect 37918 3476 37924 3528
rect 37976 3516 37982 3528
rect 38013 3519 38071 3525
rect 38013 3516 38025 3519
rect 37976 3488 38025 3516
rect 37976 3476 37982 3488
rect 38013 3485 38025 3488
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 25685 3451 25743 3457
rect 25685 3417 25697 3451
rect 25731 3448 25743 3451
rect 25958 3448 25964 3460
rect 25731 3420 25964 3448
rect 25731 3417 25743 3420
rect 25685 3411 25743 3417
rect 25958 3408 25964 3420
rect 26016 3408 26022 3460
rect 33045 3451 33103 3457
rect 33045 3448 33057 3451
rect 26068 3420 33057 3448
rect 24412 3352 25544 3380
rect 25590 3340 25596 3392
rect 25648 3380 25654 3392
rect 26068 3380 26096 3420
rect 33045 3417 33057 3420
rect 33091 3417 33103 3451
rect 34422 3448 34428 3460
rect 33045 3411 33103 3417
rect 33152 3420 34428 3448
rect 25648 3352 26096 3380
rect 25648 3340 25654 3352
rect 26142 3340 26148 3392
rect 26200 3380 26206 3392
rect 26200 3352 26245 3380
rect 26200 3340 26206 3352
rect 26418 3340 26424 3392
rect 26476 3380 26482 3392
rect 26881 3383 26939 3389
rect 26881 3380 26893 3383
rect 26476 3352 26893 3380
rect 26476 3340 26482 3352
rect 26881 3349 26893 3352
rect 26927 3349 26939 3383
rect 26881 3343 26939 3349
rect 28166 3340 28172 3392
rect 28224 3380 28230 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 28224 3352 28733 3380
rect 28224 3340 28230 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 28810 3340 28816 3392
rect 28868 3380 28874 3392
rect 30742 3380 30748 3392
rect 28868 3352 30748 3380
rect 28868 3340 28874 3352
rect 30742 3340 30748 3352
rect 30800 3340 30806 3392
rect 31110 3380 31116 3392
rect 31071 3352 31116 3380
rect 31110 3340 31116 3352
rect 31168 3340 31174 3392
rect 31202 3340 31208 3392
rect 31260 3380 31266 3392
rect 33152 3380 33180 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 33594 3380 33600 3392
rect 31260 3352 33180 3380
rect 33555 3352 33600 3380
rect 31260 3340 31266 3352
rect 33594 3340 33600 3352
rect 33652 3340 33658 3392
rect 33686 3340 33692 3392
rect 33744 3380 33750 3392
rect 34885 3383 34943 3389
rect 34885 3380 34897 3383
rect 33744 3352 34897 3380
rect 33744 3340 33750 3352
rect 34885 3349 34897 3352
rect 34931 3349 34943 3383
rect 34885 3343 34943 3349
rect 35529 3383 35587 3389
rect 35529 3349 35541 3383
rect 35575 3380 35587 3383
rect 36630 3380 36636 3392
rect 35575 3352 36636 3380
rect 35575 3349 35587 3352
rect 35529 3343 35587 3349
rect 36630 3340 36636 3352
rect 36688 3340 36694 3392
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5534 3176 5540 3188
rect 2332 3148 5540 3176
rect 2332 3117 2360 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5868 3148 6009 3176
rect 5868 3136 5874 3148
rect 5997 3145 6009 3148
rect 6043 3176 6055 3179
rect 6043 3148 16620 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 2317 3111 2375 3117
rect 2317 3077 2329 3111
rect 2363 3077 2375 3111
rect 3970 3108 3976 3120
rect 3542 3080 3976 3108
rect 2317 3071 2375 3077
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 6822 3108 6828 3120
rect 5750 3080 6828 3108
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 8110 3108 8116 3120
rect 8050 3080 8116 3108
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 8570 3108 8576 3120
rect 8531 3080 8576 3108
rect 8570 3068 8576 3080
rect 8628 3068 8634 3120
rect 9582 3108 9588 3120
rect 9416 3080 9588 3108
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 9306 3040 9312 3052
rect 8036 3012 9312 3040
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 2041 2975 2099 2981
rect 2041 2972 2053 2975
rect 1728 2944 2053 2972
rect 1728 2932 1734 2944
rect 2041 2941 2053 2944
rect 2087 2972 2099 2975
rect 4062 2972 4068 2984
rect 2087 2944 4068 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 4062 2932 4068 2944
rect 4120 2972 4126 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4120 2944 4261 2972
rect 4120 2932 4126 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 4249 2935 4307 2941
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2972 4583 2975
rect 5258 2972 5264 2984
rect 4571 2944 5264 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5552 2944 6837 2972
rect 3786 2904 3792 2916
rect 3747 2876 3792 2904
rect 3786 2864 3792 2876
rect 3844 2864 3850 2916
rect 3602 2796 3608 2848
rect 3660 2836 3666 2848
rect 5552 2836 5580 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 8036 2972 8064 3012
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9416 3049 9444 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 9677 3111 9735 3117
rect 9677 3077 9689 3111
rect 9723 3108 9735 3111
rect 9950 3108 9956 3120
rect 9723 3080 9956 3108
rect 9723 3077 9735 3080
rect 9677 3071 9735 3077
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10962 3108 10968 3120
rect 10902 3080 10968 3108
rect 10962 3068 10968 3080
rect 11020 3068 11026 3120
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 12618 3108 12624 3120
rect 11940 3080 12624 3108
rect 11940 3068 11946 3080
rect 12618 3068 12624 3080
rect 12676 3068 12682 3120
rect 14458 3108 14464 3120
rect 13924 3080 14464 3108
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 13722 3000 13728 3052
rect 13780 3000 13786 3052
rect 10686 2972 10692 2984
rect 6972 2944 8064 2972
rect 8128 2944 10692 2972
rect 6972 2932 6978 2944
rect 3660 2808 5580 2836
rect 3660 2796 3666 2808
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 8128 2836 8156 2944
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 12342 2972 12348 2984
rect 10928 2944 11928 2972
rect 12303 2944 12348 2972
rect 10928 2932 10934 2944
rect 11149 2907 11207 2913
rect 11149 2873 11161 2907
rect 11195 2904 11207 2907
rect 11606 2904 11612 2916
rect 11195 2876 11612 2904
rect 11195 2873 11207 2876
rect 11149 2867 11207 2873
rect 11606 2864 11612 2876
rect 11664 2864 11670 2916
rect 5684 2808 8156 2836
rect 5684 2796 5690 2808
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 11793 2839 11851 2845
rect 11793 2836 11805 2839
rect 9548 2808 11805 2836
rect 9548 2796 9554 2808
rect 11793 2805 11805 2808
rect 11839 2805 11851 2839
rect 11900 2836 11928 2944
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12618 2932 12624 2984
rect 12676 2972 12682 2984
rect 13924 2972 13952 3080
rect 14458 3068 14464 3080
rect 14516 3108 14522 3120
rect 14829 3111 14887 3117
rect 14829 3108 14841 3111
rect 14516 3080 14841 3108
rect 14516 3068 14522 3080
rect 14829 3077 14841 3080
rect 14875 3077 14887 3111
rect 16482 3108 16488 3120
rect 16054 3080 16488 3108
rect 14829 3071 14887 3077
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 12676 2944 13952 2972
rect 12676 2932 12682 2944
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 16298 2972 16304 2984
rect 16080 2944 16304 2972
rect 16080 2932 16086 2944
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 13354 2836 13360 2848
rect 11900 2808 13360 2836
rect 11793 2799 11851 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 14093 2839 14151 2845
rect 14093 2805 14105 2839
rect 14139 2836 14151 2839
rect 14918 2836 14924 2848
rect 14139 2808 14924 2836
rect 14139 2805 14151 2808
rect 14093 2799 14151 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 16592 2836 16620 3148
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 19886 3176 19892 3188
rect 17828 3148 19892 3176
rect 17828 3136 17834 3148
rect 19886 3136 19892 3148
rect 19944 3136 19950 3188
rect 26418 3176 26424 3188
rect 19996 3148 26424 3176
rect 19996 3108 20024 3148
rect 26418 3136 26424 3148
rect 26476 3136 26482 3188
rect 33042 3176 33048 3188
rect 27349 3148 33048 3176
rect 21910 3108 21916 3120
rect 18630 3080 20024 3108
rect 20838 3080 21916 3108
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 22465 3111 22523 3117
rect 22465 3077 22477 3111
rect 22511 3108 22523 3111
rect 25314 3108 25320 3120
rect 22511 3080 25320 3108
rect 22511 3077 22523 3080
rect 22465 3071 22523 3077
rect 25314 3068 25320 3080
rect 25372 3068 25378 3120
rect 25590 3108 25596 3120
rect 25551 3080 25596 3108
rect 25590 3068 25596 3080
rect 25648 3068 25654 3120
rect 25682 3068 25688 3120
rect 25740 3108 25746 3120
rect 26602 3108 26608 3120
rect 25740 3080 25785 3108
rect 26563 3080 26608 3108
rect 25740 3068 25746 3080
rect 26602 3068 26608 3080
rect 26660 3068 26666 3120
rect 27349 3117 27377 3148
rect 33042 3136 33048 3148
rect 33100 3136 33106 3188
rect 34330 3176 34336 3188
rect 34291 3148 34336 3176
rect 34330 3136 34336 3148
rect 34388 3136 34394 3188
rect 35618 3176 35624 3188
rect 35579 3148 35624 3176
rect 35618 3136 35624 3148
rect 35676 3136 35682 3188
rect 27341 3111 27399 3117
rect 27341 3077 27353 3111
rect 27387 3077 27399 3111
rect 27341 3071 27399 3077
rect 27430 3068 27436 3120
rect 27488 3108 27494 3120
rect 33686 3108 33692 3120
rect 27488 3080 29224 3108
rect 27488 3068 27494 3080
rect 16850 3000 16856 3052
rect 16908 3040 16914 3052
rect 17126 3040 17132 3052
rect 16908 3012 17132 3040
rect 16908 3000 16914 3012
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 19208 3012 19349 3040
rect 19208 3000 19214 3012
rect 19337 3009 19349 3012
rect 19383 3009 19395 3043
rect 23842 3040 23848 3052
rect 23803 3012 23848 3040
rect 19337 3003 19395 3009
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 24578 3000 24584 3052
rect 24636 3040 24642 3052
rect 24673 3043 24731 3049
rect 24673 3040 24685 3043
rect 24636 3012 24685 3040
rect 24636 3000 24642 3012
rect 24673 3009 24685 3012
rect 24719 3009 24731 3043
rect 28534 3040 28540 3052
rect 28495 3012 28540 3040
rect 24673 3003 24731 3009
rect 28534 3000 28540 3012
rect 28592 3000 28598 3052
rect 29196 3049 29224 3080
rect 29656 3080 33692 3108
rect 29656 3049 29684 3080
rect 33686 3068 33692 3080
rect 33744 3068 33750 3120
rect 29181 3043 29239 3049
rect 29181 3009 29193 3043
rect 29227 3009 29239 3043
rect 29181 3003 29239 3009
rect 29641 3043 29699 3049
rect 29641 3009 29653 3043
rect 29687 3009 29699 3043
rect 29641 3003 29699 3009
rect 30285 3043 30343 3049
rect 30285 3009 30297 3043
rect 30331 3009 30343 3043
rect 30285 3003 30343 3009
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 19058 2972 19064 2984
rect 17451 2944 19064 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19613 2975 19671 2981
rect 19613 2941 19625 2975
rect 19659 2972 19671 2975
rect 20990 2972 20996 2984
rect 19659 2944 20996 2972
rect 19659 2941 19671 2944
rect 19613 2935 19671 2941
rect 20990 2932 20996 2944
rect 21048 2932 21054 2984
rect 22370 2972 22376 2984
rect 21836 2960 22048 2972
rect 22112 2960 22232 2972
rect 21836 2944 22232 2960
rect 22331 2944 22376 2972
rect 21085 2907 21143 2913
rect 21085 2873 21097 2907
rect 21131 2904 21143 2907
rect 21358 2904 21364 2916
rect 21131 2876 21364 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 18414 2836 18420 2848
rect 16592 2808 18420 2836
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 18877 2839 18935 2845
rect 18877 2805 18889 2839
rect 18923 2836 18935 2839
rect 21836 2836 21864 2944
rect 22020 2932 22140 2944
rect 21910 2864 21916 2916
rect 21968 2904 21974 2916
rect 22204 2904 22232 2944
rect 22370 2932 22376 2944
rect 22428 2932 22434 2984
rect 22646 2972 22652 2984
rect 22607 2944 22652 2972
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 25866 2972 25872 2984
rect 23768 2944 25872 2972
rect 23768 2904 23796 2944
rect 25866 2932 25872 2944
rect 25924 2932 25930 2984
rect 27246 2972 27252 2984
rect 27207 2944 27252 2972
rect 27246 2932 27252 2944
rect 27304 2932 27310 2984
rect 29730 2972 29736 2984
rect 27349 2944 29040 2972
rect 29691 2944 29736 2972
rect 23934 2904 23940 2916
rect 21968 2876 22140 2904
rect 22204 2876 23796 2904
rect 23895 2876 23940 2904
rect 21968 2864 21974 2876
rect 18923 2808 21864 2836
rect 22112 2836 22140 2876
rect 23934 2864 23940 2876
rect 23992 2864 23998 2916
rect 24302 2864 24308 2916
rect 24360 2904 24366 2916
rect 24489 2907 24547 2913
rect 24489 2904 24501 2907
rect 24360 2876 24501 2904
rect 24360 2864 24366 2876
rect 24489 2873 24501 2876
rect 24535 2873 24547 2907
rect 24489 2867 24547 2873
rect 25038 2864 25044 2916
rect 25096 2904 25102 2916
rect 27349 2904 27377 2944
rect 25096 2876 27377 2904
rect 25096 2864 25102 2876
rect 27614 2864 27620 2916
rect 27672 2904 27678 2916
rect 27801 2907 27859 2913
rect 27801 2904 27813 2907
rect 27672 2876 27813 2904
rect 27672 2864 27678 2876
rect 27801 2873 27813 2876
rect 27847 2873 27859 2907
rect 27801 2867 27859 2873
rect 27890 2864 27896 2916
rect 27948 2904 27954 2916
rect 29012 2913 29040 2944
rect 29730 2932 29736 2944
rect 29788 2932 29794 2984
rect 30300 2972 30328 3003
rect 30834 3000 30840 3052
rect 30892 3040 30898 3052
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30892 3012 30941 3040
rect 30892 3000 30898 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 31573 3043 31631 3049
rect 31573 3040 31585 3043
rect 30929 3003 30987 3009
rect 31496 3012 31585 3040
rect 31202 2972 31208 2984
rect 30300 2944 31208 2972
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31496 2972 31524 3012
rect 31573 3009 31585 3012
rect 31619 3009 31631 3043
rect 31573 3003 31631 3009
rect 31662 3000 31668 3052
rect 31720 3040 31726 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31720 3012 32321 3040
rect 31720 3000 31726 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 32766 3000 32772 3052
rect 32824 3040 32830 3052
rect 32953 3043 33011 3049
rect 32953 3040 32965 3043
rect 32824 3012 32965 3040
rect 32824 3000 32830 3012
rect 32953 3009 32965 3012
rect 32999 3009 33011 3043
rect 33597 3043 33655 3049
rect 33597 3040 33609 3043
rect 32953 3003 33011 3009
rect 33060 3012 33609 3040
rect 33060 2972 33088 3012
rect 33597 3009 33609 3012
rect 33643 3009 33655 3043
rect 33597 3003 33655 3009
rect 34241 3043 34299 3049
rect 34241 3009 34253 3043
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 31496 2944 33088 2972
rect 28353 2907 28411 2913
rect 28353 2904 28365 2907
rect 27948 2876 28365 2904
rect 27948 2864 27954 2876
rect 28353 2873 28365 2876
rect 28399 2873 28411 2907
rect 28353 2867 28411 2873
rect 28997 2907 29055 2913
rect 28997 2873 29009 2907
rect 29043 2873 29055 2907
rect 28997 2867 29055 2873
rect 29086 2864 29092 2916
rect 29144 2904 29150 2916
rect 30377 2907 30435 2913
rect 30377 2904 30389 2907
rect 29144 2876 30389 2904
rect 29144 2864 29150 2876
rect 30377 2873 30389 2876
rect 30423 2873 30435 2907
rect 30377 2867 30435 2873
rect 30742 2864 30748 2916
rect 30800 2904 30806 2916
rect 31021 2907 31079 2913
rect 31021 2904 31033 2907
rect 30800 2876 31033 2904
rect 30800 2864 30806 2876
rect 31021 2873 31033 2876
rect 31067 2873 31079 2907
rect 31021 2867 31079 2873
rect 28166 2836 28172 2848
rect 22112 2808 28172 2836
rect 18923 2805 18935 2808
rect 18877 2799 18935 2805
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 28718 2796 28724 2848
rect 28776 2836 28782 2848
rect 31496 2836 31524 2944
rect 33134 2932 33140 2984
rect 33192 2972 33198 2984
rect 34256 2972 34284 3003
rect 34422 3000 34428 3052
rect 34480 3040 34486 3052
rect 34885 3043 34943 3049
rect 34885 3040 34897 3043
rect 34480 3012 34897 3040
rect 34480 3000 34486 3012
rect 34885 3009 34897 3012
rect 34931 3009 34943 3043
rect 35526 3040 35532 3052
rect 35487 3012 35532 3040
rect 34885 3003 34943 3009
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 35866 3012 36369 3040
rect 33192 2944 34284 2972
rect 33192 2932 33198 2944
rect 35434 2932 35440 2984
rect 35492 2972 35498 2984
rect 35866 2972 35894 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 36357 3003 36415 3009
rect 36630 3000 36636 3052
rect 36688 3040 36694 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 36688 3012 38025 3040
rect 36688 3000 36694 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 35492 2944 35894 2972
rect 35492 2932 35498 2944
rect 33226 2864 33232 2916
rect 33284 2904 33290 2916
rect 33689 2907 33747 2913
rect 33689 2904 33701 2907
rect 33284 2876 33701 2904
rect 33284 2864 33290 2876
rect 33689 2873 33701 2876
rect 33735 2873 33747 2907
rect 33689 2867 33747 2873
rect 31662 2836 31668 2848
rect 28776 2808 31524 2836
rect 31623 2808 31668 2836
rect 28776 2796 28782 2808
rect 31662 2796 31668 2808
rect 31720 2796 31726 2848
rect 32398 2836 32404 2848
rect 32359 2808 32404 2836
rect 32398 2796 32404 2808
rect 32456 2796 32462 2848
rect 32858 2796 32864 2848
rect 32916 2836 32922 2848
rect 33045 2839 33103 2845
rect 33045 2836 33057 2839
rect 32916 2808 33057 2836
rect 32916 2796 32922 2808
rect 33045 2805 33057 2808
rect 33091 2805 33103 2839
rect 33045 2799 33103 2805
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34977 2839 35035 2845
rect 34977 2836 34989 2839
rect 34572 2808 34989 2836
rect 34572 2796 34578 2808
rect 34977 2805 34989 2808
rect 35023 2805 35035 2839
rect 36170 2836 36176 2848
rect 36131 2808 36176 2836
rect 34977 2799 35035 2805
rect 36170 2796 36176 2808
rect 36228 2796 36234 2848
rect 38197 2839 38255 2845
rect 38197 2805 38209 2839
rect 38243 2836 38255 2839
rect 38654 2836 38660 2848
rect 38243 2808 38660 2836
rect 38243 2805 38255 2808
rect 38197 2799 38255 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 3418 2592 3424 2604
rect 3476 2632 3482 2644
rect 5626 2632 5632 2644
rect 3476 2604 5632 2632
rect 3476 2592 3482 2604
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 13630 2632 13636 2644
rect 8220 2604 13636 2632
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 3786 2496 3792 2508
rect 1995 2468 3792 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4120 2468 4261 2496
rect 4120 2456 4126 2468
rect 4249 2465 4261 2468
rect 4295 2496 4307 2499
rect 6546 2496 6552 2508
rect 4295 2468 6552 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 6546 2456 6552 2468
rect 6604 2496 6610 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6604 2468 6837 2496
rect 6604 2456 6610 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 8220 2414 8248 2604
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 15470 2632 15476 2644
rect 13771 2604 15476 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 19426 2632 19432 2644
rect 18923 2604 19432 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 21174 2632 21180 2644
rect 19576 2604 21180 2632
rect 19576 2592 19582 2604
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 23474 2632 23480 2644
rect 21284 2604 23480 2632
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 11882 2564 11888 2576
rect 11195 2536 11888 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 11882 2524 11888 2536
rect 11940 2524 11946 2576
rect 18414 2524 18420 2576
rect 18472 2564 18478 2576
rect 18472 2536 19564 2564
rect 18472 2524 18478 2536
rect 9401 2499 9459 2505
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 9766 2496 9772 2508
rect 9447 2468 9772 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 9824 2468 11989 2496
rect 9824 2456 9830 2468
rect 11977 2465 11989 2468
rect 12023 2496 12035 2499
rect 12342 2496 12348 2508
rect 12023 2468 12348 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 12342 2456 12348 2468
rect 12400 2456 12406 2508
rect 14550 2496 14556 2508
rect 14511 2468 14556 2496
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 16022 2496 16028 2508
rect 14875 2468 16028 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 17126 2496 17132 2508
rect 17039 2468 17132 2496
rect 17126 2456 17132 2468
rect 17184 2496 17190 2508
rect 19150 2496 19156 2508
rect 17184 2468 19156 2496
rect 17184 2456 17190 2468
rect 19150 2456 19156 2468
rect 19208 2496 19214 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19208 2468 19441 2496
rect 19208 2456 19214 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19536 2496 19564 2536
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 19536 2468 19717 2496
rect 19429 2459 19487 2465
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 21284 2496 21312 2604
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 23842 2632 23848 2644
rect 23803 2604 23848 2632
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 24854 2592 24860 2644
rect 24912 2632 24918 2644
rect 24912 2604 25452 2632
rect 24912 2592 24918 2604
rect 25317 2567 25375 2573
rect 25317 2564 25329 2567
rect 22388 2536 25329 2564
rect 22388 2505 22416 2536
rect 25317 2533 25329 2536
rect 25363 2533 25375 2567
rect 25424 2564 25452 2604
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 26384 2604 27169 2632
rect 26384 2592 26390 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 27264 2604 31754 2632
rect 27264 2564 27292 2604
rect 25424 2536 27292 2564
rect 25317 2527 25375 2533
rect 19705 2459 19763 2465
rect 20824 2468 21312 2496
rect 22373 2499 22431 2505
rect 20824 2414 20852 2468
rect 22373 2465 22385 2499
rect 22419 2465 22431 2499
rect 22646 2496 22652 2508
rect 22607 2468 22652 2496
rect 22373 2459 22431 2465
rect 22646 2456 22652 2468
rect 22704 2456 22710 2508
rect 27890 2496 27896 2508
rect 25332 2468 27896 2496
rect 22186 2428 22192 2440
rect 22066 2400 22192 2428
rect 4062 2360 4068 2372
rect 3174 2332 4068 2360
rect 4062 2320 4068 2332
rect 4120 2320 4126 2372
rect 4525 2363 4583 2369
rect 4525 2329 4537 2363
rect 4571 2329 4583 2363
rect 5902 2360 5908 2372
rect 5750 2332 5908 2360
rect 4525 2323 4583 2329
rect 4540 2292 4568 2323
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 7101 2363 7159 2369
rect 7101 2329 7113 2363
rect 7147 2329 7159 2363
rect 8938 2360 8944 2372
rect 7101 2323 7159 2329
rect 8404 2332 8944 2360
rect 5810 2292 5816 2304
rect 4540 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 7116 2292 7144 2323
rect 8404 2292 8432 2332
rect 8938 2320 8944 2332
rect 8996 2320 9002 2372
rect 9677 2363 9735 2369
rect 9677 2329 9689 2363
rect 9723 2360 9735 2363
rect 9950 2360 9956 2372
rect 9723 2332 9956 2360
rect 9723 2329 9735 2332
rect 9677 2323 9735 2329
rect 9950 2320 9956 2332
rect 10008 2320 10014 2372
rect 12158 2360 12164 2372
rect 10902 2332 12164 2360
rect 12158 2320 12164 2332
rect 12216 2320 12222 2372
rect 12253 2363 12311 2369
rect 12253 2329 12265 2363
rect 12299 2329 12311 2363
rect 13722 2360 13728 2372
rect 13478 2332 13728 2360
rect 12253 2323 12311 2329
rect 6043 2264 8432 2292
rect 8573 2295 8631 2301
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 8573 2261 8585 2295
rect 8619 2292 8631 2295
rect 10594 2292 10600 2304
rect 8619 2264 10600 2292
rect 8619 2261 8631 2264
rect 8573 2255 8631 2261
rect 10594 2252 10600 2264
rect 10652 2292 10658 2304
rect 12268 2292 12296 2323
rect 13722 2320 13728 2332
rect 13780 2320 13786 2372
rect 17310 2360 17316 2372
rect 16054 2332 17316 2360
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 17405 2363 17463 2369
rect 17405 2329 17417 2363
rect 17451 2329 17463 2363
rect 22066 2360 22094 2400
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23348 2400 24041 2428
rect 23348 2388 23354 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24762 2428 24768 2440
rect 24723 2400 24768 2428
rect 24029 2391 24087 2397
rect 24762 2388 24768 2400
rect 24820 2388 24826 2440
rect 25225 2431 25283 2437
rect 25225 2397 25237 2431
rect 25271 2428 25283 2431
rect 25332 2428 25360 2468
rect 27890 2456 27896 2468
rect 27948 2456 27954 2508
rect 28077 2499 28135 2505
rect 28077 2465 28089 2499
rect 28123 2496 28135 2499
rect 28626 2496 28632 2508
rect 28123 2468 28632 2496
rect 28123 2465 28135 2468
rect 28077 2459 28135 2465
rect 28626 2456 28632 2468
rect 28684 2456 28690 2508
rect 30006 2496 30012 2508
rect 29967 2468 30012 2496
rect 30006 2456 30012 2468
rect 30064 2456 30070 2508
rect 25866 2428 25872 2440
rect 25271 2400 25360 2428
rect 25827 2400 25872 2428
rect 25271 2397 25283 2400
rect 25225 2391 25283 2397
rect 25866 2388 25872 2400
rect 25924 2428 25930 2440
rect 26142 2428 26148 2440
rect 25924 2400 26148 2428
rect 25924 2388 25930 2400
rect 26142 2388 26148 2400
rect 26200 2388 26206 2440
rect 27338 2428 27344 2440
rect 27299 2400 27344 2428
rect 27338 2388 27344 2400
rect 27396 2388 27402 2440
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27764 2400 27813 2428
rect 27764 2388 27770 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29052 2400 29745 2428
rect 29052 2388 29058 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 22462 2360 22468 2372
rect 18630 2332 19656 2360
rect 17405 2323 17463 2329
rect 10652 2264 12296 2292
rect 10652 2252 10658 2264
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16298 2292 16304 2304
rect 16172 2264 16304 2292
rect 16172 2252 16178 2264
rect 16298 2252 16304 2264
rect 16356 2252 16362 2304
rect 17420 2292 17448 2323
rect 19518 2292 19524 2304
rect 17420 2264 19524 2292
rect 19518 2252 19524 2264
rect 19576 2252 19582 2304
rect 19628 2292 19656 2332
rect 21008 2332 22094 2360
rect 22423 2332 22468 2360
rect 21008 2292 21036 2332
rect 22462 2320 22468 2332
rect 22520 2320 22526 2372
rect 31036 2360 31064 2391
rect 24596 2332 31064 2360
rect 31726 2360 31754 2604
rect 32122 2592 32128 2644
rect 32180 2632 32186 2644
rect 32180 2604 37780 2632
rect 32180 2592 32186 2604
rect 36081 2567 36139 2573
rect 36081 2533 36093 2567
rect 36127 2564 36139 2567
rect 37182 2564 37188 2576
rect 36127 2536 37188 2564
rect 36127 2533 36139 2536
rect 36081 2527 36139 2533
rect 37182 2524 37188 2536
rect 37240 2524 37246 2576
rect 34606 2456 34612 2508
rect 34664 2496 34670 2508
rect 37752 2505 37780 2604
rect 37737 2499 37795 2505
rect 34664 2468 36676 2496
rect 34664 2456 34670 2468
rect 32306 2428 32312 2440
rect 32267 2400 32312 2428
rect 32306 2388 32312 2400
rect 32364 2388 32370 2440
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33560 2400 33609 2428
rect 33560 2388 33566 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36648 2437 36676 2468
rect 37737 2465 37749 2499
rect 37783 2465 37795 2499
rect 37737 2459 37795 2465
rect 36633 2431 36691 2437
rect 35952 2400 35997 2428
rect 35952 2388 35958 2400
rect 36633 2397 36645 2431
rect 36679 2397 36691 2431
rect 37458 2428 37464 2440
rect 37419 2400 37464 2428
rect 36633 2391 36691 2397
rect 37458 2388 37464 2400
rect 37516 2388 37522 2440
rect 33042 2360 33048 2372
rect 31726 2332 33048 2360
rect 24596 2301 24624 2332
rect 33042 2320 33048 2332
rect 33100 2320 33106 2372
rect 19628 2264 21036 2292
rect 24581 2295 24639 2301
rect 24581 2261 24593 2295
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 26142 2252 26148 2304
rect 26200 2292 26206 2304
rect 29546 2292 29552 2304
rect 26200 2264 29552 2292
rect 26200 2252 26206 2264
rect 29546 2252 29552 2264
rect 29604 2252 29610 2304
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30340 2264 31217 2292
rect 30340 2252 30346 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32272 2264 32505 2292
rect 32272 2252 32278 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 33560 2264 33793 2292
rect 33560 2252 33566 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34204 2264 35081 2292
rect 34204 2252 34210 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 36817 2295 36875 2301
rect 36817 2292 36829 2295
rect 36780 2264 36829 2292
rect 36780 2252 36786 2264
rect 36817 2261 36829 2264
rect 36863 2261 36875 2295
rect 36817 2255 36875 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 2774 2048 2780 2100
rect 2832 2088 2838 2100
rect 4706 2088 4712 2100
rect 2832 2060 4712 2088
rect 2832 2048 2838 2060
rect 4706 2048 4712 2060
rect 4764 2048 4770 2100
rect 22462 2048 22468 2100
rect 22520 2088 22526 2100
rect 26786 2088 26792 2100
rect 22520 2060 26792 2088
rect 22520 2048 22526 2060
rect 26786 2048 26792 2060
rect 26844 2048 26850 2100
rect 17310 1980 17316 2032
rect 17368 2020 17374 2032
rect 17368 1992 24716 2020
rect 17368 1980 17374 1992
rect 13630 1912 13636 1964
rect 13688 1952 13694 1964
rect 23658 1952 23664 1964
rect 13688 1924 23664 1952
rect 13688 1912 13694 1924
rect 23658 1912 23664 1924
rect 23716 1912 23722 1964
rect 24688 1952 24716 1992
rect 24762 1980 24768 2032
rect 24820 2020 24826 2032
rect 30834 2020 30840 2032
rect 24820 1992 30840 2020
rect 24820 1980 24826 1992
rect 30834 1980 30840 1992
rect 30892 1980 30898 2032
rect 31110 1952 31116 1964
rect 24688 1924 31116 1952
rect 31110 1912 31116 1924
rect 31168 1912 31174 1964
rect 17954 1844 17960 1896
rect 18012 1884 18018 1896
rect 29086 1884 29092 1896
rect 18012 1856 29092 1884
rect 18012 1844 18018 1856
rect 29086 1844 29092 1856
rect 29144 1844 29150 1896
rect 9950 1776 9956 1828
rect 10008 1816 10014 1828
rect 18874 1816 18880 1828
rect 10008 1788 18880 1816
rect 10008 1776 10014 1788
rect 18874 1776 18880 1788
rect 18932 1776 18938 1828
rect 20990 1776 20996 1828
rect 21048 1816 21054 1828
rect 21048 1788 31754 1816
rect 21048 1776 21054 1788
rect 11790 1708 11796 1760
rect 11848 1748 11854 1760
rect 18414 1748 18420 1760
rect 11848 1720 18420 1748
rect 11848 1708 11854 1720
rect 18414 1708 18420 1720
rect 18472 1708 18478 1760
rect 27798 1748 27804 1760
rect 18524 1720 27804 1748
rect 16298 1640 16304 1692
rect 16356 1680 16362 1692
rect 18524 1680 18552 1720
rect 27798 1708 27804 1720
rect 27856 1708 27862 1760
rect 16356 1652 18552 1680
rect 16356 1640 16362 1652
rect 19978 1640 19984 1692
rect 20036 1680 20042 1692
rect 27338 1680 27344 1692
rect 20036 1652 27344 1680
rect 20036 1640 20042 1652
rect 27338 1640 27344 1652
rect 27396 1640 27402 1692
rect 31726 1680 31754 1788
rect 36170 1680 36176 1692
rect 31726 1652 36176 1680
rect 36170 1640 36176 1652
rect 36228 1640 36234 1692
rect 23198 1572 23204 1624
rect 23256 1612 23262 1624
rect 27430 1612 27436 1624
rect 23256 1584 27436 1612
rect 23256 1572 23262 1584
rect 27430 1572 27436 1584
rect 27488 1572 27494 1624
rect 21266 1504 21272 1556
rect 21324 1544 21330 1556
rect 23290 1544 23296 1556
rect 21324 1516 23296 1544
rect 21324 1504 21330 1516
rect 23290 1504 23296 1516
rect 23348 1504 23354 1556
rect 12158 1436 12164 1488
rect 12216 1476 12222 1488
rect 25222 1476 25228 1488
rect 12216 1448 25228 1476
rect 12216 1436 12222 1448
rect 25222 1436 25228 1448
rect 25280 1436 25286 1488
rect 21174 1368 21180 1420
rect 21232 1408 21238 1420
rect 25130 1408 25136 1420
rect 21232 1380 25136 1408
rect 21232 1368 21238 1380
rect 25130 1368 25136 1380
rect 25188 1368 25194 1420
rect 20438 1300 20444 1352
rect 20496 1340 20502 1352
rect 31386 1340 31392 1352
rect 20496 1312 31392 1340
rect 20496 1300 20502 1312
rect 31386 1300 31392 1312
rect 31444 1300 31450 1352
rect 10962 1232 10968 1284
rect 11020 1272 11026 1284
rect 34514 1272 34520 1284
rect 11020 1244 34520 1272
rect 11020 1232 11026 1244
rect 34514 1232 34520 1244
rect 34572 1232 34578 1284
rect 13262 1164 13268 1216
rect 13320 1204 13326 1216
rect 29270 1204 29276 1216
rect 13320 1176 29276 1204
rect 13320 1164 13326 1176
rect 29270 1164 29276 1176
rect 29328 1164 29334 1216
rect 16390 1096 16396 1148
rect 16448 1136 16454 1148
rect 32398 1136 32404 1148
rect 16448 1108 32404 1136
rect 16448 1096 16454 1108
rect 32398 1096 32404 1108
rect 32456 1096 32462 1148
rect 11974 1028 11980 1080
rect 12032 1068 12038 1080
rect 27154 1068 27160 1080
rect 12032 1040 27160 1068
rect 12032 1028 12038 1040
rect 27154 1028 27160 1040
rect 27212 1028 27218 1080
rect 4062 960 4068 1012
rect 4120 1000 4126 1012
rect 31662 1000 31668 1012
rect 4120 972 31668 1000
rect 4120 960 4126 972
rect 31662 960 31668 972
rect 31720 960 31726 1012
<< via1 >>
rect 16580 37612 16632 37664
rect 19156 37612 19208 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16580 37340 16632 37392
rect 1584 37315 1636 37324
rect 1584 37281 1593 37315
rect 1593 37281 1627 37315
rect 1627 37281 1636 37315
rect 1584 37272 1636 37281
rect 3884 37272 3936 37324
rect 5816 37272 5868 37324
rect 8392 37272 8444 37324
rect 16120 37272 16172 37324
rect 23572 37340 23624 37392
rect 22560 37272 22612 37324
rect 24860 37315 24912 37324
rect 24860 37281 24869 37315
rect 24869 37281 24903 37315
rect 24903 37281 24912 37315
rect 24860 37272 24912 37281
rect 27712 37272 27764 37324
rect 29644 37272 29696 37324
rect 1860 37247 1912 37256
rect 1860 37213 1869 37247
rect 1869 37213 1903 37247
rect 1903 37213 1912 37247
rect 1860 37204 1912 37213
rect 2780 37204 2832 37256
rect 4252 37247 4304 37256
rect 4252 37213 4261 37247
rect 4261 37213 4295 37247
rect 4295 37213 4304 37247
rect 4252 37204 4304 37213
rect 5172 37204 5224 37256
rect 6828 37247 6880 37256
rect 6828 37213 6837 37247
rect 6837 37213 6871 37247
rect 6871 37213 6880 37247
rect 6828 37204 6880 37213
rect 7104 37204 7156 37256
rect 9404 37247 9456 37256
rect 9404 37213 9413 37247
rect 9413 37213 9447 37247
rect 9447 37213 9456 37247
rect 9404 37204 9456 37213
rect 5264 37111 5316 37120
rect 5264 37077 5273 37111
rect 5273 37077 5307 37111
rect 5307 37077 5316 37111
rect 5264 37068 5316 37077
rect 11060 37136 11112 37188
rect 11612 37204 11664 37256
rect 12440 37204 12492 37256
rect 13544 37204 13596 37256
rect 14924 37247 14976 37256
rect 14924 37213 14933 37247
rect 14933 37213 14967 37247
rect 14967 37213 14976 37247
rect 14924 37204 14976 37213
rect 18052 37204 18104 37256
rect 18420 37204 18472 37256
rect 21272 37204 21324 37256
rect 16580 37136 16632 37188
rect 21088 37136 21140 37188
rect 24492 37204 24544 37256
rect 25780 37204 25832 37256
rect 26332 37247 26384 37256
rect 26332 37213 26341 37247
rect 26341 37213 26375 37247
rect 26375 37213 26384 37247
rect 26332 37204 26384 37213
rect 28080 37247 28132 37256
rect 28080 37213 28089 37247
rect 28089 37213 28123 37247
rect 28123 37213 28132 37247
rect 28080 37204 28132 37213
rect 29000 37204 29052 37256
rect 31024 37247 31076 37256
rect 31024 37213 31033 37247
rect 31033 37213 31067 37247
rect 31067 37213 31076 37247
rect 31024 37204 31076 37213
rect 32128 37204 32180 37256
rect 32404 37204 32456 37256
rect 34888 37247 34940 37256
rect 34888 37213 34897 37247
rect 34897 37213 34931 37247
rect 34931 37213 34940 37247
rect 34888 37204 34940 37213
rect 35532 37204 35584 37256
rect 37464 37247 37516 37256
rect 37464 37213 37473 37247
rect 37473 37213 37507 37247
rect 37507 37213 37516 37247
rect 37464 37204 37516 37213
rect 10324 37068 10376 37120
rect 11704 37111 11756 37120
rect 11704 37077 11713 37111
rect 11713 37077 11747 37111
rect 11747 37077 11756 37111
rect 11704 37068 11756 37077
rect 12348 37111 12400 37120
rect 12348 37077 12357 37111
rect 12357 37077 12391 37111
rect 12391 37077 12400 37111
rect 12348 37068 12400 37077
rect 12532 37068 12584 37120
rect 14096 37111 14148 37120
rect 14096 37077 14105 37111
rect 14105 37077 14139 37111
rect 14139 37077 14148 37111
rect 14096 37068 14148 37077
rect 14832 37068 14884 37120
rect 18052 37068 18104 37120
rect 19984 37068 20036 37120
rect 20352 37068 20404 37120
rect 23020 37068 23072 37120
rect 26424 37068 26476 37120
rect 27160 37068 27212 37120
rect 29828 37068 29880 37120
rect 30932 37068 30984 37120
rect 32220 37068 32272 37120
rect 33140 37068 33192 37120
rect 34520 37068 34572 37120
rect 36084 37068 36136 37120
rect 37372 37068 37424 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1768 36907 1820 36916
rect 1768 36873 1777 36907
rect 1777 36873 1811 36907
rect 1811 36873 1820 36907
rect 1768 36864 1820 36873
rect 4252 36864 4304 36916
rect 11796 36864 11848 36916
rect 18420 36864 18472 36916
rect 19340 36864 19392 36916
rect 31024 36864 31076 36916
rect 37464 36864 37516 36916
rect 9404 36796 9456 36848
rect 15568 36796 15620 36848
rect 1952 36728 2004 36780
rect 3148 36771 3200 36780
rect 3148 36737 3157 36771
rect 3157 36737 3191 36771
rect 3191 36737 3200 36771
rect 3148 36728 3200 36737
rect 9036 36728 9088 36780
rect 11796 36728 11848 36780
rect 16764 36728 16816 36780
rect 28080 36796 28132 36848
rect 38108 36839 38160 36848
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 23480 36771 23532 36780
rect 23480 36737 23489 36771
rect 23489 36737 23523 36771
rect 23523 36737 23532 36771
rect 23480 36728 23532 36737
rect 28448 36771 28500 36780
rect 28448 36737 28457 36771
rect 28457 36737 28491 36771
rect 28491 36737 28500 36771
rect 28448 36728 28500 36737
rect 38108 36805 38117 36839
rect 38117 36805 38151 36839
rect 38151 36805 38160 36839
rect 38108 36796 38160 36805
rect 35440 36728 35492 36780
rect 36360 36771 36412 36780
rect 36360 36737 36369 36771
rect 36369 36737 36403 36771
rect 36403 36737 36412 36771
rect 36360 36728 36412 36737
rect 4620 36660 4672 36712
rect 6736 36592 6788 36644
rect 34888 36592 34940 36644
rect 5816 36524 5868 36576
rect 8024 36524 8076 36576
rect 15476 36524 15528 36576
rect 21640 36524 21692 36576
rect 33140 36524 33192 36576
rect 36820 36524 36872 36576
rect 37280 36524 37332 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 39304 36320 39356 36372
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 36820 36159 36872 36168
rect 36820 36125 36829 36159
rect 36829 36125 36863 36159
rect 36863 36125 36872 36159
rect 36820 36116 36872 36125
rect 33324 36048 33376 36100
rect 2688 35980 2740 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 12532 35819 12584 35828
rect 12532 35785 12541 35819
rect 12541 35785 12575 35819
rect 12575 35785 12584 35819
rect 12532 35776 12584 35785
rect 664 35640 716 35692
rect 13912 35640 13964 35692
rect 38660 35708 38712 35760
rect 38016 35683 38068 35692
rect 38016 35649 38025 35683
rect 38025 35649 38059 35683
rect 38059 35649 38068 35683
rect 38016 35640 38068 35649
rect 5724 35436 5776 35488
rect 34520 35436 34572 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 38292 35071 38344 35080
rect 38292 35037 38301 35071
rect 38301 35037 38335 35071
rect 38335 35037 38344 35071
rect 38292 35028 38344 35037
rect 20628 34892 20680 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 33784 34552 33836 34604
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19984 33804 20036 33856
rect 37280 33804 37332 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4620 33600 4672 33652
rect 6644 33464 6696 33516
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 32404 33056 32456 33108
rect 38016 33056 38068 33108
rect 1768 32759 1820 32768
rect 1768 32725 1777 32759
rect 1777 32725 1811 32759
rect 1811 32725 1820 32759
rect 1768 32716 1820 32725
rect 5540 32852 5592 32904
rect 6828 32852 6880 32904
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 36820 32852 36872 32904
rect 38108 32827 38160 32836
rect 38108 32793 38117 32827
rect 38117 32793 38151 32827
rect 38151 32793 38160 32827
rect 38108 32784 38160 32793
rect 37832 32716 37884 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 13912 32555 13964 32564
rect 13912 32521 13921 32555
rect 13921 32521 13955 32555
rect 13955 32521 13964 32555
rect 13912 32512 13964 32521
rect 36820 32555 36872 32564
rect 36820 32521 36829 32555
rect 36829 32521 36863 32555
rect 36863 32521 36872 32555
rect 36820 32512 36872 32521
rect 12348 32444 12400 32496
rect 2596 32376 2648 32428
rect 15016 32376 15068 32428
rect 36728 32419 36780 32428
rect 36728 32385 36737 32419
rect 36737 32385 36771 32419
rect 36771 32385 36780 32419
rect 36728 32376 36780 32385
rect 38108 32419 38160 32428
rect 38108 32385 38117 32419
rect 38117 32385 38151 32419
rect 38151 32385 38160 32419
rect 38108 32376 38160 32385
rect 3424 32240 3476 32292
rect 20812 32240 20864 32292
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 15384 32215 15436 32224
rect 15384 32181 15393 32215
rect 15393 32181 15427 32215
rect 15427 32181 15436 32215
rect 15384 32172 15436 32181
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 17040 31968 17092 32020
rect 23112 31968 23164 32020
rect 11704 31900 11756 31952
rect 10416 31832 10468 31884
rect 18236 31832 18288 31884
rect 20076 31832 20128 31884
rect 5816 31807 5868 31816
rect 5816 31773 5825 31807
rect 5825 31773 5859 31807
rect 5859 31773 5868 31807
rect 5816 31764 5868 31773
rect 20352 31764 20404 31816
rect 20628 31807 20680 31816
rect 20628 31773 20637 31807
rect 20637 31773 20671 31807
rect 20671 31773 20680 31807
rect 20628 31764 20680 31773
rect 20812 31807 20864 31816
rect 20812 31773 20821 31807
rect 20821 31773 20855 31807
rect 20855 31773 20864 31807
rect 20812 31764 20864 31773
rect 21640 31807 21692 31816
rect 21640 31773 21649 31807
rect 21649 31773 21683 31807
rect 21683 31773 21692 31807
rect 21640 31764 21692 31773
rect 23020 31764 23072 31816
rect 38200 31900 38252 31952
rect 26516 31671 26568 31680
rect 26516 31637 26525 31671
rect 26525 31637 26559 31671
rect 26559 31637 26568 31671
rect 26516 31628 26568 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 33324 31467 33376 31476
rect 33324 31433 33333 31467
rect 33333 31433 33367 31467
rect 33367 31433 33376 31467
rect 33324 31424 33376 31433
rect 5724 31331 5776 31340
rect 5724 31297 5733 31331
rect 5733 31297 5767 31331
rect 5767 31297 5776 31331
rect 5724 31288 5776 31297
rect 29828 31288 29880 31340
rect 32404 31288 32456 31340
rect 6092 31084 6144 31136
rect 24032 31084 24084 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 11152 30744 11204 30796
rect 2688 30676 2740 30728
rect 8024 30719 8076 30728
rect 8024 30685 8033 30719
rect 8033 30685 8067 30719
rect 8067 30685 8076 30719
rect 8024 30676 8076 30685
rect 11060 30719 11112 30728
rect 11060 30685 11069 30719
rect 11069 30685 11103 30719
rect 11103 30685 11112 30719
rect 11060 30676 11112 30685
rect 33140 30744 33192 30796
rect 34520 30676 34572 30728
rect 38016 30719 38068 30728
rect 38016 30685 38025 30719
rect 38025 30685 38059 30719
rect 38059 30685 38068 30719
rect 38016 30676 38068 30685
rect 10968 30608 11020 30660
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 8208 30540 8260 30592
rect 13360 30540 13412 30592
rect 24952 30540 25004 30592
rect 29828 30583 29880 30592
rect 29828 30549 29837 30583
rect 29837 30549 29871 30583
rect 29871 30549 29880 30583
rect 29828 30540 29880 30549
rect 38200 30583 38252 30592
rect 38200 30549 38209 30583
rect 38209 30549 38243 30583
rect 38243 30549 38252 30583
rect 38200 30540 38252 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 23572 30336 23624 30388
rect 6644 30311 6696 30320
rect 6644 30277 6653 30311
rect 6653 30277 6687 30311
rect 6687 30277 6696 30311
rect 6644 30268 6696 30277
rect 6000 30200 6052 30252
rect 10508 30200 10560 30252
rect 17868 30200 17920 30252
rect 24860 30200 24912 30252
rect 27160 30243 27212 30252
rect 27160 30209 27169 30243
rect 27169 30209 27203 30243
rect 27203 30209 27212 30243
rect 27160 30200 27212 30209
rect 1584 30064 1636 30116
rect 11152 30064 11204 30116
rect 38016 30064 38068 30116
rect 25964 29996 26016 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 33784 29835 33836 29844
rect 33784 29801 33793 29835
rect 33793 29801 33827 29835
rect 33827 29801 33836 29835
rect 33784 29792 33836 29801
rect 5264 29656 5316 29708
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 6736 29588 6788 29640
rect 16580 29588 16632 29640
rect 26332 29588 26384 29640
rect 32496 29588 32548 29640
rect 35440 29588 35492 29640
rect 5632 29452 5684 29504
rect 7012 29452 7064 29504
rect 10692 29495 10744 29504
rect 10692 29461 10701 29495
rect 10701 29461 10735 29495
rect 10735 29461 10744 29495
rect 10692 29452 10744 29461
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 2320 29112 2372 29164
rect 14096 29112 14148 29164
rect 15476 29155 15528 29164
rect 15476 29121 15485 29155
rect 15485 29121 15519 29155
rect 15519 29121 15528 29155
rect 15476 29112 15528 29121
rect 36268 29112 36320 29164
rect 15936 29044 15988 29096
rect 1768 29019 1820 29028
rect 1768 28985 1777 29019
rect 1777 28985 1811 29019
rect 1811 28985 1820 29019
rect 1768 28976 1820 28985
rect 15200 28976 15252 29028
rect 38200 29019 38252 29028
rect 38200 28985 38209 29019
rect 38209 28985 38243 29019
rect 38243 28985 38252 29019
rect 38200 28976 38252 28985
rect 17316 28908 17368 28960
rect 23112 28908 23164 28960
rect 27712 28908 27764 28960
rect 35532 28908 35584 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 11796 28500 11848 28552
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 14096 28364 14148 28416
rect 18144 28407 18196 28416
rect 18144 28373 18153 28407
rect 18153 28373 18187 28407
rect 18187 28373 18196 28407
rect 18144 28364 18196 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 36268 28160 36320 28212
rect 15568 28024 15620 28076
rect 28080 28024 28132 28076
rect 35348 28024 35400 28076
rect 14556 27820 14608 27872
rect 22100 27820 22152 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 38292 27455 38344 27464
rect 38292 27421 38301 27455
rect 38301 27421 38335 27455
rect 38335 27421 38344 27455
rect 38292 27412 38344 27421
rect 4068 27276 4120 27328
rect 37372 27276 37424 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 6000 27072 6052 27124
rect 22468 27072 22520 27124
rect 29828 27072 29880 27124
rect 35348 27115 35400 27124
rect 35348 27081 35357 27115
rect 35357 27081 35391 27115
rect 35391 27081 35400 27115
rect 35348 27072 35400 27081
rect 16304 27004 16356 27056
rect 28448 27004 28500 27056
rect 7104 26936 7156 26988
rect 12440 26936 12492 26988
rect 15108 26936 15160 26988
rect 37740 27004 37792 27056
rect 20536 26868 20588 26920
rect 2596 26800 2648 26852
rect 12808 26775 12860 26784
rect 12808 26741 12817 26775
rect 12817 26741 12851 26775
rect 12851 26741 12860 26775
rect 12808 26732 12860 26741
rect 13728 26732 13780 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5540 26460 5592 26512
rect 1768 26367 1820 26376
rect 1768 26333 1777 26367
rect 1777 26333 1811 26367
rect 1811 26333 1820 26367
rect 1768 26324 1820 26333
rect 5724 26324 5776 26376
rect 11520 26256 11572 26308
rect 20352 26528 20404 26580
rect 35440 26528 35492 26580
rect 14004 26460 14056 26512
rect 15568 26460 15620 26512
rect 12440 26392 12492 26444
rect 13728 26367 13780 26376
rect 13728 26333 13737 26367
rect 13737 26333 13771 26367
rect 13771 26333 13780 26367
rect 13728 26324 13780 26333
rect 14372 26299 14424 26308
rect 14372 26265 14381 26299
rect 14381 26265 14415 26299
rect 14415 26265 14424 26299
rect 14372 26256 14424 26265
rect 15108 26256 15160 26308
rect 19064 26324 19116 26376
rect 29184 26324 29236 26376
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 17224 26188 17276 26240
rect 38108 26231 38160 26240
rect 38108 26197 38117 26231
rect 38117 26197 38151 26231
rect 38151 26197 38160 26231
rect 38108 26188 38160 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 32404 25984 32456 26036
rect 12808 25848 12860 25900
rect 17868 25891 17920 25900
rect 17868 25857 17877 25891
rect 17877 25857 17911 25891
rect 17911 25857 17920 25891
rect 17868 25848 17920 25857
rect 19064 25848 19116 25900
rect 27068 25848 27120 25900
rect 14464 25644 14516 25696
rect 18052 25644 18104 25696
rect 18328 25644 18380 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 32496 25440 32548 25492
rect 2688 25372 2740 25424
rect 3424 25372 3476 25424
rect 14188 25236 14240 25288
rect 21640 25304 21692 25356
rect 17224 25279 17276 25288
rect 11244 25168 11296 25220
rect 13084 25168 13136 25220
rect 17224 25245 17233 25279
rect 17233 25245 17267 25279
rect 17267 25245 17276 25279
rect 17224 25236 17276 25245
rect 27988 25279 28040 25288
rect 27988 25245 27997 25279
rect 27997 25245 28031 25279
rect 28031 25245 28040 25279
rect 27988 25236 28040 25245
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 18052 25168 18104 25220
rect 18328 25211 18380 25220
rect 18328 25177 18337 25211
rect 18337 25177 18371 25211
rect 18371 25177 18380 25211
rect 18328 25168 18380 25177
rect 19340 25168 19392 25220
rect 13912 25100 13964 25152
rect 15292 25100 15344 25152
rect 16948 25100 17000 25152
rect 17132 25100 17184 25152
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14372 24871 14424 24880
rect 14372 24837 14381 24871
rect 14381 24837 14415 24871
rect 14415 24837 14424 24871
rect 14372 24828 14424 24837
rect 16948 24828 17000 24880
rect 1584 24803 1636 24812
rect 1584 24769 1593 24803
rect 1593 24769 1627 24803
rect 1627 24769 1636 24803
rect 1584 24760 1636 24769
rect 5632 24760 5684 24812
rect 9036 24760 9088 24812
rect 15016 24760 15068 24812
rect 15384 24760 15436 24812
rect 22744 24803 22796 24812
rect 13820 24692 13872 24744
rect 15844 24692 15896 24744
rect 9588 24624 9640 24676
rect 14188 24624 14240 24676
rect 15108 24624 15160 24676
rect 22744 24769 22753 24803
rect 22753 24769 22787 24803
rect 22787 24769 22796 24803
rect 22744 24760 22796 24769
rect 18052 24692 18104 24744
rect 17960 24624 18012 24676
rect 1768 24599 1820 24608
rect 1768 24565 1777 24599
rect 1777 24565 1811 24599
rect 1811 24565 1820 24599
rect 1768 24556 1820 24565
rect 10140 24556 10192 24608
rect 10232 24556 10284 24608
rect 10692 24556 10744 24608
rect 15476 24556 15528 24608
rect 15752 24556 15804 24608
rect 16948 24556 17000 24608
rect 22836 24556 22888 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1584 24352 1636 24404
rect 30748 24352 30800 24404
rect 12164 24284 12216 24336
rect 12808 24284 12860 24336
rect 15844 24327 15896 24336
rect 8484 24216 8536 24268
rect 10876 24216 10928 24268
rect 10968 24216 11020 24268
rect 15016 24259 15068 24268
rect 15016 24225 15025 24259
rect 15025 24225 15059 24259
rect 15059 24225 15068 24259
rect 15016 24216 15068 24225
rect 2688 24148 2740 24200
rect 9036 24148 9088 24200
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 9496 24080 9548 24132
rect 11244 24191 11296 24200
rect 11244 24157 11253 24191
rect 11253 24157 11287 24191
rect 11287 24157 11296 24191
rect 11244 24148 11296 24157
rect 12348 24123 12400 24132
rect 12348 24089 12357 24123
rect 12357 24089 12391 24123
rect 12391 24089 12400 24123
rect 12348 24080 12400 24089
rect 14372 24123 14424 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 9404 24055 9456 24064
rect 9404 24021 9413 24055
rect 9413 24021 9447 24055
rect 9447 24021 9456 24055
rect 9404 24012 9456 24021
rect 11152 24012 11204 24064
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 14372 24089 14381 24123
rect 14381 24089 14415 24123
rect 14415 24089 14424 24123
rect 14372 24080 14424 24089
rect 14464 24123 14516 24132
rect 14464 24089 14473 24123
rect 14473 24089 14507 24123
rect 14507 24089 14516 24123
rect 15844 24293 15853 24327
rect 15853 24293 15887 24327
rect 15887 24293 15896 24327
rect 15844 24284 15896 24293
rect 15476 24259 15528 24268
rect 15476 24225 15485 24259
rect 15485 24225 15519 24259
rect 15519 24225 15528 24259
rect 15476 24216 15528 24225
rect 15568 24216 15620 24268
rect 23388 24284 23440 24336
rect 16948 24259 17000 24268
rect 16948 24225 16957 24259
rect 16957 24225 16991 24259
rect 16991 24225 17000 24259
rect 16948 24216 17000 24225
rect 19616 24216 19668 24268
rect 20168 24216 20220 24268
rect 20536 24259 20588 24268
rect 20536 24225 20545 24259
rect 20545 24225 20579 24259
rect 20579 24225 20588 24259
rect 20536 24216 20588 24225
rect 18880 24148 18932 24200
rect 37464 24191 37516 24200
rect 37464 24157 37473 24191
rect 37473 24157 37507 24191
rect 37507 24157 37516 24191
rect 37464 24148 37516 24157
rect 37924 24148 37976 24200
rect 14464 24080 14516 24089
rect 17960 24080 18012 24132
rect 19616 24123 19668 24132
rect 19616 24089 19625 24123
rect 19625 24089 19659 24123
rect 19659 24089 19668 24123
rect 19616 24080 19668 24089
rect 16304 24012 16356 24064
rect 18328 24012 18380 24064
rect 22652 24055 22704 24064
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 10876 23808 10928 23860
rect 15568 23808 15620 23860
rect 9404 23740 9456 23792
rect 10508 23740 10560 23792
rect 15108 23783 15160 23792
rect 15108 23749 15117 23783
rect 15117 23749 15151 23783
rect 15151 23749 15160 23783
rect 15108 23740 15160 23749
rect 5540 23672 5592 23724
rect 9496 23672 9548 23724
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 14004 23715 14056 23724
rect 14004 23681 14013 23715
rect 14013 23681 14047 23715
rect 14047 23681 14056 23715
rect 14004 23672 14056 23681
rect 16120 23715 16172 23724
rect 16120 23681 16129 23715
rect 16129 23681 16163 23715
rect 16163 23681 16172 23715
rect 16120 23672 16172 23681
rect 18880 23715 18932 23724
rect 11060 23604 11112 23656
rect 12716 23647 12768 23656
rect 12716 23613 12725 23647
rect 12725 23613 12759 23647
rect 12759 23613 12768 23647
rect 12716 23604 12768 23613
rect 13912 23604 13964 23656
rect 9404 23536 9456 23588
rect 14372 23536 14424 23588
rect 8576 23468 8628 23520
rect 13728 23468 13780 23520
rect 15384 23604 15436 23656
rect 18880 23681 18889 23715
rect 18889 23681 18923 23715
rect 18923 23681 18932 23715
rect 18880 23672 18932 23681
rect 28356 23808 28408 23860
rect 30748 23851 30800 23860
rect 30748 23817 30757 23851
rect 30757 23817 30791 23851
rect 30791 23817 30800 23851
rect 30748 23808 30800 23817
rect 22652 23715 22704 23724
rect 22652 23681 22661 23715
rect 22661 23681 22695 23715
rect 22695 23681 22704 23715
rect 22652 23672 22704 23681
rect 22836 23715 22888 23724
rect 22836 23681 22845 23715
rect 22845 23681 22879 23715
rect 22879 23681 22888 23715
rect 22836 23672 22888 23681
rect 17868 23604 17920 23656
rect 17960 23536 18012 23588
rect 20444 23604 20496 23656
rect 30104 23672 30156 23724
rect 18512 23536 18564 23588
rect 18420 23468 18472 23520
rect 23020 23511 23072 23520
rect 23020 23477 23029 23511
rect 23029 23477 23063 23511
rect 23063 23477 23072 23511
rect 23020 23468 23072 23477
rect 38016 23468 38068 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 17500 23264 17552 23316
rect 19432 23264 19484 23316
rect 10324 23196 10376 23248
rect 10232 23128 10284 23180
rect 12072 23196 12124 23248
rect 16580 23196 16632 23248
rect 24952 23196 25004 23248
rect 18512 23171 18564 23180
rect 18512 23137 18521 23171
rect 18521 23137 18555 23171
rect 18555 23137 18564 23171
rect 18512 23128 18564 23137
rect 1952 23060 2004 23112
rect 8576 23103 8628 23112
rect 8576 23069 8585 23103
rect 8585 23069 8619 23103
rect 8619 23069 8628 23103
rect 8576 23060 8628 23069
rect 9312 23060 9364 23112
rect 10692 23103 10744 23112
rect 10692 23069 10701 23103
rect 10701 23069 10735 23103
rect 10735 23069 10744 23103
rect 10692 23060 10744 23069
rect 12716 23060 12768 23112
rect 20628 23128 20680 23180
rect 22744 23128 22796 23180
rect 20812 23060 20864 23112
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 12532 22992 12584 23044
rect 18328 23035 18380 23044
rect 18328 23001 18337 23035
rect 18337 23001 18371 23035
rect 18371 23001 18380 23035
rect 18328 22992 18380 23001
rect 10784 22924 10836 22976
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 13176 22967 13228 22976
rect 13176 22933 13185 22967
rect 13185 22933 13219 22967
rect 13219 22933 13228 22967
rect 13176 22924 13228 22933
rect 14740 22967 14792 22976
rect 14740 22933 14749 22967
rect 14749 22933 14783 22967
rect 14783 22933 14792 22967
rect 14740 22924 14792 22933
rect 20260 22967 20312 22976
rect 20260 22933 20269 22967
rect 20269 22933 20303 22967
rect 20303 22933 20312 22967
rect 20260 22924 20312 22933
rect 21456 22924 21508 22976
rect 23480 22924 23532 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2320 22763 2372 22772
rect 2320 22729 2329 22763
rect 2329 22729 2363 22763
rect 2363 22729 2372 22763
rect 2320 22720 2372 22729
rect 10232 22720 10284 22772
rect 4068 22652 4120 22704
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 2504 22627 2556 22636
rect 2504 22593 2513 22627
rect 2513 22593 2547 22627
rect 2547 22593 2556 22627
rect 2504 22584 2556 22593
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 7196 22584 7248 22593
rect 9312 22584 9364 22636
rect 10692 22720 10744 22772
rect 11060 22720 11112 22772
rect 11428 22720 11480 22772
rect 15108 22720 15160 22772
rect 15660 22720 15712 22772
rect 11336 22652 11388 22704
rect 15752 22695 15804 22704
rect 9404 22516 9456 22568
rect 11888 22584 11940 22636
rect 13636 22627 13688 22636
rect 12164 22516 12216 22568
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 14648 22584 14700 22636
rect 15752 22661 15761 22695
rect 15761 22661 15795 22695
rect 15795 22661 15804 22695
rect 15752 22652 15804 22661
rect 13728 22516 13780 22568
rect 15844 22516 15896 22568
rect 23020 22720 23072 22772
rect 29184 22763 29236 22772
rect 29184 22729 29193 22763
rect 29193 22729 29227 22763
rect 29227 22729 29236 22763
rect 29184 22720 29236 22729
rect 17132 22695 17184 22704
rect 17132 22661 17141 22695
rect 17141 22661 17175 22695
rect 17175 22661 17184 22695
rect 17132 22652 17184 22661
rect 19340 22652 19392 22704
rect 20536 22652 20588 22704
rect 23480 22695 23532 22704
rect 23480 22661 23489 22695
rect 23489 22661 23523 22695
rect 23523 22661 23532 22695
rect 23480 22652 23532 22661
rect 25044 22695 25096 22704
rect 25044 22661 25053 22695
rect 25053 22661 25087 22695
rect 25087 22661 25096 22695
rect 25044 22652 25096 22661
rect 26516 22652 26568 22704
rect 20260 22584 20312 22636
rect 20628 22584 20680 22636
rect 21456 22584 21508 22636
rect 29092 22627 29144 22636
rect 29092 22593 29101 22627
rect 29101 22593 29135 22627
rect 29135 22593 29144 22627
rect 29092 22584 29144 22593
rect 2504 22448 2556 22500
rect 9128 22448 9180 22500
rect 11244 22448 11296 22500
rect 11428 22448 11480 22500
rect 20352 22516 20404 22568
rect 24032 22516 24084 22568
rect 24308 22559 24360 22568
rect 24308 22525 24317 22559
rect 24317 22525 24351 22559
rect 24351 22525 24360 22559
rect 24308 22516 24360 22525
rect 24952 22559 25004 22568
rect 24952 22525 24961 22559
rect 24961 22525 24995 22559
rect 24995 22525 25004 22559
rect 24952 22516 25004 22525
rect 1768 22423 1820 22432
rect 1768 22389 1777 22423
rect 1777 22389 1811 22423
rect 1811 22389 1820 22423
rect 1768 22380 1820 22389
rect 7288 22380 7340 22432
rect 9772 22380 9824 22432
rect 10508 22380 10560 22432
rect 17408 22448 17460 22500
rect 38200 22491 38252 22500
rect 13728 22423 13780 22432
rect 13728 22389 13737 22423
rect 13737 22389 13771 22423
rect 13771 22389 13780 22423
rect 13728 22380 13780 22389
rect 15016 22423 15068 22432
rect 15016 22389 15025 22423
rect 15025 22389 15059 22423
rect 15059 22389 15068 22423
rect 15016 22380 15068 22389
rect 16856 22380 16908 22432
rect 18328 22380 18380 22432
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 20996 22423 21048 22432
rect 20996 22389 21005 22423
rect 21005 22389 21039 22423
rect 21039 22389 21048 22423
rect 20996 22380 21048 22389
rect 22744 22380 22796 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1768 22176 1820 22228
rect 12716 22176 12768 22228
rect 13268 22176 13320 22228
rect 17684 22176 17736 22228
rect 17408 22108 17460 22160
rect 9956 22040 10008 22092
rect 1952 22015 2004 22024
rect 1952 21981 1961 22015
rect 1961 21981 1995 22015
rect 1995 21981 2004 22015
rect 1952 21972 2004 21981
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 12256 22040 12308 22092
rect 12624 22040 12676 22092
rect 13176 22040 13228 22092
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 14924 22040 14976 22092
rect 16304 22040 16356 22092
rect 18236 22083 18288 22092
rect 18236 22049 18245 22083
rect 18245 22049 18279 22083
rect 18279 22049 18288 22083
rect 18236 22040 18288 22049
rect 20076 22040 20128 22092
rect 20168 22083 20220 22092
rect 20168 22049 20177 22083
rect 20177 22049 20211 22083
rect 20211 22049 20220 22083
rect 20168 22040 20220 22049
rect 23296 22083 23348 22092
rect 23296 22049 23305 22083
rect 23305 22049 23339 22083
rect 23339 22049 23348 22083
rect 23296 22040 23348 22049
rect 27988 22040 28040 22092
rect 12532 21972 12584 22024
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 24584 21972 24636 22024
rect 38108 21972 38160 22024
rect 38292 22015 38344 22024
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 7196 21904 7248 21956
rect 1584 21836 1636 21888
rect 7288 21836 7340 21888
rect 7380 21836 7432 21888
rect 10600 21836 10652 21888
rect 10784 21947 10836 21956
rect 10784 21913 10793 21947
rect 10793 21913 10827 21947
rect 10827 21913 10836 21947
rect 11704 21947 11756 21956
rect 10784 21904 10836 21913
rect 11704 21913 11713 21947
rect 11713 21913 11747 21947
rect 11747 21913 11756 21947
rect 11704 21904 11756 21913
rect 14832 21947 14884 21956
rect 14832 21913 14841 21947
rect 14841 21913 14875 21947
rect 14875 21913 14884 21947
rect 14832 21904 14884 21913
rect 16028 21904 16080 21956
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 12348 21836 12400 21888
rect 16672 21904 16724 21956
rect 17776 21904 17828 21956
rect 18420 21904 18472 21956
rect 21088 21947 21140 21956
rect 19432 21836 19484 21888
rect 21088 21913 21097 21947
rect 21097 21913 21131 21947
rect 21131 21913 21140 21947
rect 21088 21904 21140 21913
rect 21180 21947 21232 21956
rect 21180 21913 21189 21947
rect 21189 21913 21223 21947
rect 21223 21913 21232 21947
rect 22652 21947 22704 21956
rect 21180 21904 21232 21913
rect 22652 21913 22661 21947
rect 22661 21913 22695 21947
rect 22695 21913 22704 21947
rect 22652 21904 22704 21913
rect 22744 21947 22796 21956
rect 22744 21913 22753 21947
rect 22753 21913 22787 21947
rect 22787 21913 22796 21947
rect 22744 21904 22796 21913
rect 23756 21879 23808 21888
rect 23756 21845 23765 21879
rect 23765 21845 23799 21879
rect 23799 21845 23808 21879
rect 23756 21836 23808 21845
rect 27528 21836 27580 21888
rect 34704 21836 34756 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 8392 21632 8444 21684
rect 10968 21632 11020 21684
rect 11060 21632 11112 21684
rect 8852 21564 8904 21616
rect 11704 21632 11756 21684
rect 17500 21675 17552 21684
rect 1584 21539 1636 21548
rect 1584 21505 1593 21539
rect 1593 21505 1627 21539
rect 1627 21505 1636 21539
rect 1584 21496 1636 21505
rect 7380 21496 7432 21548
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 10324 21496 10376 21548
rect 9864 21360 9916 21412
rect 1768 21335 1820 21344
rect 1768 21301 1777 21335
rect 1777 21301 1811 21335
rect 1811 21301 1820 21335
rect 1768 21292 1820 21301
rect 6920 21292 6972 21344
rect 8668 21292 8720 21344
rect 11152 21428 11204 21480
rect 13268 21564 13320 21616
rect 13820 21607 13872 21616
rect 13820 21573 13829 21607
rect 13829 21573 13863 21607
rect 13863 21573 13872 21607
rect 13820 21564 13872 21573
rect 15200 21564 15252 21616
rect 17500 21641 17509 21675
rect 17509 21641 17543 21675
rect 17543 21641 17552 21675
rect 17500 21632 17552 21641
rect 17868 21632 17920 21684
rect 19340 21564 19392 21616
rect 21088 21632 21140 21684
rect 22652 21675 22704 21684
rect 22652 21641 22661 21675
rect 22661 21641 22695 21675
rect 22695 21641 22704 21675
rect 22652 21632 22704 21641
rect 27528 21607 27580 21616
rect 16304 21496 16356 21548
rect 18604 21539 18656 21548
rect 12348 21428 12400 21480
rect 11060 21360 11112 21412
rect 12716 21428 12768 21480
rect 13820 21428 13872 21480
rect 15200 21471 15252 21480
rect 15200 21437 15209 21471
rect 15209 21437 15243 21471
rect 15243 21437 15252 21471
rect 15200 21428 15252 21437
rect 10784 21292 10836 21344
rect 14372 21360 14424 21412
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 19708 21496 19760 21548
rect 20904 21496 20956 21548
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 21272 21496 21324 21548
rect 23020 21496 23072 21548
rect 23756 21496 23808 21548
rect 23848 21496 23900 21548
rect 25504 21539 25556 21548
rect 25504 21505 25513 21539
rect 25513 21505 25547 21539
rect 25547 21505 25556 21539
rect 25504 21496 25556 21505
rect 17776 21360 17828 21412
rect 27068 21428 27120 21480
rect 27528 21573 27537 21607
rect 27537 21573 27571 21607
rect 27571 21573 27580 21607
rect 27528 21564 27580 21573
rect 27620 21607 27672 21616
rect 27620 21573 27629 21607
rect 27629 21573 27663 21607
rect 27663 21573 27672 21607
rect 27620 21564 27672 21573
rect 37372 21496 37424 21548
rect 30840 21428 30892 21480
rect 20720 21360 20772 21412
rect 15568 21292 15620 21344
rect 16028 21292 16080 21344
rect 16580 21292 16632 21344
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 19616 21292 19668 21344
rect 19708 21292 19760 21344
rect 20812 21292 20864 21344
rect 24032 21335 24084 21344
rect 24032 21301 24041 21335
rect 24041 21301 24075 21335
rect 24075 21301 24084 21335
rect 24032 21292 24084 21301
rect 24676 21335 24728 21344
rect 24676 21301 24685 21335
rect 24685 21301 24719 21335
rect 24719 21301 24728 21335
rect 24676 21292 24728 21301
rect 29460 21292 29512 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 8300 21088 8352 21140
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 8944 21088 8996 21140
rect 11152 21088 11204 21140
rect 5172 20952 5224 21004
rect 11060 21020 11112 21072
rect 16028 21020 16080 21072
rect 16120 21020 16172 21072
rect 17040 21020 17092 21072
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 7380 20927 7432 20936
rect 7380 20893 7389 20927
rect 7389 20893 7423 20927
rect 7423 20893 7432 20927
rect 7380 20884 7432 20893
rect 5264 20816 5316 20868
rect 12348 20995 12400 21004
rect 12348 20961 12357 20995
rect 12357 20961 12391 20995
rect 12391 20961 12400 20995
rect 12348 20952 12400 20961
rect 12624 20952 12676 21004
rect 13728 20952 13780 21004
rect 14556 20995 14608 21004
rect 14556 20961 14565 20995
rect 14565 20961 14599 20995
rect 14599 20961 14608 20995
rect 14556 20952 14608 20961
rect 15016 20952 15068 21004
rect 15844 20995 15896 21004
rect 15844 20961 15853 20995
rect 15853 20961 15887 20995
rect 15887 20961 15896 20995
rect 15844 20952 15896 20961
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 17592 21088 17644 21140
rect 21272 21088 21324 21140
rect 24584 21131 24636 21140
rect 24584 21097 24593 21131
rect 24593 21097 24627 21131
rect 24627 21097 24636 21131
rect 24584 21088 24636 21097
rect 25504 21088 25556 21140
rect 33968 21088 34020 21140
rect 23296 21020 23348 21072
rect 27712 21063 27764 21072
rect 27712 21029 27721 21063
rect 27721 21029 27755 21063
rect 27755 21029 27764 21063
rect 27712 21020 27764 21029
rect 20720 20995 20772 21004
rect 20720 20961 20729 20995
rect 20729 20961 20763 20995
rect 20763 20961 20772 20995
rect 20720 20952 20772 20961
rect 20996 20952 21048 21004
rect 24676 20952 24728 21004
rect 34796 20952 34848 21004
rect 8944 20884 8996 20936
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 10232 20884 10284 20936
rect 15384 20884 15436 20936
rect 8576 20816 8628 20868
rect 9680 20748 9732 20800
rect 10048 20748 10100 20800
rect 10508 20859 10560 20868
rect 10508 20825 10517 20859
rect 10517 20825 10551 20859
rect 10551 20825 10560 20859
rect 10508 20816 10560 20825
rect 10876 20816 10928 20868
rect 16764 20816 16816 20868
rect 17500 20859 17552 20868
rect 17500 20825 17509 20859
rect 17509 20825 17543 20859
rect 17543 20825 17552 20859
rect 17500 20816 17552 20825
rect 12256 20748 12308 20800
rect 19616 20859 19668 20868
rect 19616 20825 19625 20859
rect 19625 20825 19659 20859
rect 19659 20825 19668 20859
rect 19616 20816 19668 20825
rect 20168 20748 20220 20800
rect 20812 20748 20864 20800
rect 24124 20884 24176 20936
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 24032 20816 24084 20868
rect 27804 20816 27856 20868
rect 38200 20791 38252 20800
rect 38200 20757 38209 20791
rect 38209 20757 38243 20791
rect 38243 20757 38252 20791
rect 38200 20748 38252 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 7012 20519 7064 20528
rect 7012 20485 7021 20519
rect 7021 20485 7055 20519
rect 7055 20485 7064 20519
rect 7012 20476 7064 20485
rect 8024 20476 8076 20528
rect 8852 20544 8904 20596
rect 8944 20544 8996 20596
rect 8668 20519 8720 20528
rect 8668 20485 8677 20519
rect 8677 20485 8711 20519
rect 8711 20485 8720 20519
rect 8668 20476 8720 20485
rect 9680 20476 9732 20528
rect 10048 20476 10100 20528
rect 11244 20476 11296 20528
rect 12716 20544 12768 20596
rect 12992 20544 13044 20596
rect 16764 20544 16816 20596
rect 16672 20476 16724 20528
rect 12624 20408 12676 20460
rect 13176 20408 13228 20460
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 16304 20408 16356 20460
rect 16764 20408 16816 20460
rect 18604 20544 18656 20596
rect 19156 20544 19208 20596
rect 23848 20544 23900 20596
rect 24124 20587 24176 20596
rect 24124 20553 24133 20587
rect 24133 20553 24167 20587
rect 24167 20553 24176 20587
rect 24124 20544 24176 20553
rect 21088 20476 21140 20528
rect 19156 20451 19208 20460
rect 10232 20383 10284 20392
rect 7012 20272 7064 20324
rect 6184 20204 6236 20256
rect 10232 20349 10241 20383
rect 10241 20349 10275 20383
rect 10275 20349 10284 20383
rect 10232 20340 10284 20349
rect 11980 20340 12032 20392
rect 14372 20340 14424 20392
rect 15384 20340 15436 20392
rect 9128 20272 9180 20324
rect 13268 20204 13320 20256
rect 13544 20247 13596 20256
rect 13544 20213 13553 20247
rect 13553 20213 13587 20247
rect 13587 20213 13596 20247
rect 13544 20204 13596 20213
rect 15016 20272 15068 20324
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 20628 20408 20680 20460
rect 21640 20408 21692 20460
rect 24768 20408 24820 20460
rect 29184 20451 29236 20460
rect 29184 20417 29193 20451
rect 29193 20417 29227 20451
rect 29227 20417 29236 20451
rect 29184 20408 29236 20417
rect 33968 20451 34020 20460
rect 33968 20417 33977 20451
rect 33977 20417 34011 20451
rect 34011 20417 34020 20451
rect 33968 20408 34020 20417
rect 37832 20408 37884 20460
rect 20720 20340 20772 20392
rect 17684 20272 17736 20324
rect 20168 20272 20220 20324
rect 14464 20204 14516 20256
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 17776 20204 17828 20256
rect 20352 20204 20404 20256
rect 27528 20272 27580 20324
rect 21456 20204 21508 20256
rect 28724 20204 28776 20256
rect 33508 20204 33560 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 10048 20000 10100 20052
rect 12348 20000 12400 20052
rect 11796 19932 11848 19984
rect 12992 20000 13044 20052
rect 15660 20000 15712 20052
rect 16580 20043 16632 20052
rect 16580 20009 16589 20043
rect 16589 20009 16623 20043
rect 16623 20009 16632 20043
rect 16580 20000 16632 20009
rect 19432 20000 19484 20052
rect 12900 19932 12952 19984
rect 12532 19864 12584 19916
rect 13360 19864 13412 19916
rect 13728 19907 13780 19916
rect 13728 19873 13737 19907
rect 13737 19873 13771 19907
rect 13771 19873 13780 19907
rect 13728 19864 13780 19873
rect 14556 19864 14608 19916
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 16948 19864 17000 19916
rect 7564 19796 7616 19848
rect 8300 19796 8352 19848
rect 9220 19796 9272 19848
rect 10968 19796 11020 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 20352 20000 20404 20052
rect 20628 20000 20680 20052
rect 20812 20043 20864 20052
rect 20812 20009 20821 20043
rect 20821 20009 20855 20043
rect 20855 20009 20864 20043
rect 20812 20000 20864 20009
rect 21456 19839 21508 19848
rect 6736 19660 6788 19712
rect 6920 19771 6972 19780
rect 6920 19737 6929 19771
rect 6929 19737 6963 19771
rect 6963 19737 6972 19771
rect 6920 19728 6972 19737
rect 7104 19728 7156 19780
rect 7472 19771 7524 19780
rect 7472 19737 7481 19771
rect 7481 19737 7515 19771
rect 7515 19737 7524 19771
rect 7472 19728 7524 19737
rect 10416 19728 10468 19780
rect 11612 19771 11664 19780
rect 11612 19737 11621 19771
rect 11621 19737 11655 19771
rect 11655 19737 11664 19771
rect 11612 19728 11664 19737
rect 13544 19728 13596 19780
rect 15108 19771 15160 19780
rect 15108 19737 15117 19771
rect 15117 19737 15151 19771
rect 15151 19737 15160 19771
rect 15108 19728 15160 19737
rect 17224 19728 17276 19780
rect 17500 19771 17552 19780
rect 17500 19737 17509 19771
rect 17509 19737 17543 19771
rect 17543 19737 17552 19771
rect 17500 19728 17552 19737
rect 17592 19728 17644 19780
rect 21456 19805 21465 19839
rect 21465 19805 21499 19839
rect 21499 19805 21508 19839
rect 21456 19796 21508 19805
rect 26240 19932 26292 19984
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 13360 19660 13412 19712
rect 14280 19660 14332 19712
rect 14648 19660 14700 19712
rect 21824 19728 21876 19780
rect 27804 19839 27856 19848
rect 27804 19805 27813 19839
rect 27813 19805 27847 19839
rect 27847 19805 27856 19839
rect 27804 19796 27856 19805
rect 27252 19728 27304 19780
rect 29184 19796 29236 19848
rect 34704 19796 34756 19848
rect 28632 19728 28684 19780
rect 23756 19660 23808 19712
rect 26148 19660 26200 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 6828 19456 6880 19508
rect 7380 19456 7432 19508
rect 8024 19456 8076 19508
rect 9036 19456 9088 19508
rect 11612 19456 11664 19508
rect 11704 19456 11756 19508
rect 12900 19456 12952 19508
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 6920 19320 6972 19372
rect 7196 19363 7248 19372
rect 7196 19329 7205 19363
rect 7205 19329 7239 19363
rect 7239 19329 7248 19363
rect 7932 19363 7984 19372
rect 7196 19320 7248 19329
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 10692 19388 10744 19440
rect 10876 19388 10928 19440
rect 12348 19388 12400 19440
rect 14648 19431 14700 19440
rect 14648 19397 14657 19431
rect 14657 19397 14691 19431
rect 14691 19397 14700 19431
rect 14648 19388 14700 19397
rect 14924 19388 14976 19440
rect 10508 19363 10560 19372
rect 10508 19329 10517 19363
rect 10517 19329 10551 19363
rect 10551 19329 10560 19363
rect 10508 19320 10560 19329
rect 10784 19320 10836 19372
rect 8300 19252 8352 19304
rect 9220 19252 9272 19304
rect 8116 19184 8168 19236
rect 11612 19252 11664 19304
rect 12348 19252 12400 19304
rect 13268 19320 13320 19372
rect 15200 19431 15252 19440
rect 15200 19397 15209 19431
rect 15209 19397 15243 19431
rect 15243 19397 15252 19431
rect 15200 19388 15252 19397
rect 15568 19388 15620 19440
rect 23480 19456 23532 19508
rect 17592 19388 17644 19440
rect 17960 19431 18012 19440
rect 17960 19397 17969 19431
rect 17969 19397 18003 19431
rect 18003 19397 18012 19431
rect 17960 19388 18012 19397
rect 18052 19388 18104 19440
rect 19432 19388 19484 19440
rect 13268 19184 13320 19236
rect 17684 19320 17736 19372
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 19524 19252 19576 19304
rect 14556 19184 14608 19236
rect 4712 19116 4764 19168
rect 7932 19116 7984 19168
rect 9128 19116 9180 19168
rect 9588 19116 9640 19168
rect 13544 19116 13596 19168
rect 14740 19116 14792 19168
rect 28724 19363 28776 19372
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 30104 19363 30156 19372
rect 30104 19329 30113 19363
rect 30113 19329 30147 19363
rect 30147 19329 30156 19363
rect 30104 19320 30156 19329
rect 30196 19363 30248 19372
rect 30196 19329 30205 19363
rect 30205 19329 30239 19363
rect 30239 19329 30248 19363
rect 38108 19363 38160 19372
rect 30196 19320 30248 19329
rect 38108 19329 38117 19363
rect 38117 19329 38151 19363
rect 38151 19329 38160 19363
rect 38108 19320 38160 19329
rect 16672 19184 16724 19236
rect 17224 19184 17276 19236
rect 20904 19184 20956 19236
rect 17868 19116 17920 19168
rect 22560 19116 22612 19168
rect 28540 19159 28592 19168
rect 28540 19125 28549 19159
rect 28549 19125 28583 19159
rect 28583 19125 28592 19159
rect 28540 19116 28592 19125
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 6000 18912 6052 18964
rect 8484 18912 8536 18964
rect 10324 18912 10376 18964
rect 16856 18912 16908 18964
rect 16948 18912 17000 18964
rect 21088 18912 21140 18964
rect 7472 18844 7524 18896
rect 7288 18776 7340 18828
rect 9220 18819 9272 18828
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 5816 18708 5868 18760
rect 7380 18708 7432 18760
rect 7748 18751 7800 18760
rect 7748 18717 7757 18751
rect 7757 18717 7791 18751
rect 7791 18717 7800 18751
rect 7748 18708 7800 18717
rect 8300 18708 8352 18760
rect 8760 18708 8812 18760
rect 9220 18785 9229 18819
rect 9229 18785 9263 18819
rect 9263 18785 9272 18819
rect 9220 18776 9272 18785
rect 10140 18776 10192 18828
rect 13728 18844 13780 18896
rect 14556 18844 14608 18896
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 12348 18776 12400 18828
rect 12992 18776 13044 18828
rect 14648 18776 14700 18828
rect 15844 18776 15896 18828
rect 12164 18708 12216 18760
rect 10784 18683 10836 18692
rect 10784 18649 10793 18683
rect 10793 18649 10827 18683
rect 10827 18649 10836 18683
rect 10784 18640 10836 18649
rect 14464 18708 14516 18760
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 16120 18708 16172 18760
rect 17408 18776 17460 18828
rect 19524 18819 19576 18828
rect 19524 18785 19533 18819
rect 19533 18785 19567 18819
rect 19567 18785 19576 18819
rect 19524 18776 19576 18785
rect 26516 18844 26568 18896
rect 22468 18819 22520 18828
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 24676 18776 24728 18828
rect 17224 18708 17276 18760
rect 18512 18708 18564 18760
rect 20904 18708 20956 18760
rect 23756 18751 23808 18760
rect 23756 18717 23765 18751
rect 23765 18717 23799 18751
rect 23799 18717 23808 18751
rect 23756 18708 23808 18717
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 27528 18776 27580 18828
rect 35992 18776 36044 18828
rect 4344 18572 4396 18624
rect 6460 18572 6512 18624
rect 7104 18572 7156 18624
rect 9128 18572 9180 18624
rect 9220 18572 9272 18624
rect 11336 18572 11388 18624
rect 12716 18572 12768 18624
rect 15292 18572 15344 18624
rect 15568 18572 15620 18624
rect 16304 18572 16356 18624
rect 17040 18572 17092 18624
rect 20996 18640 21048 18692
rect 22560 18683 22612 18692
rect 22560 18649 22569 18683
rect 22569 18649 22603 18683
rect 22603 18649 22612 18683
rect 22560 18640 22612 18649
rect 23204 18640 23256 18692
rect 26700 18640 26752 18692
rect 20352 18572 20404 18624
rect 23756 18572 23808 18624
rect 24860 18615 24912 18624
rect 24860 18581 24869 18615
rect 24869 18581 24903 18615
rect 24903 18581 24912 18615
rect 24860 18572 24912 18581
rect 25504 18615 25556 18624
rect 25504 18581 25513 18615
rect 25513 18581 25547 18615
rect 25547 18581 25556 18615
rect 25504 18572 25556 18581
rect 26332 18572 26384 18624
rect 27712 18572 27764 18624
rect 28356 18572 28408 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 5816 18411 5868 18420
rect 5816 18377 5825 18411
rect 5825 18377 5859 18411
rect 5859 18377 5868 18411
rect 5816 18368 5868 18377
rect 10784 18368 10836 18420
rect 11060 18368 11112 18420
rect 11704 18368 11756 18420
rect 4344 18343 4396 18352
rect 4344 18309 4353 18343
rect 4353 18309 4387 18343
rect 4387 18309 4396 18343
rect 4344 18300 4396 18309
rect 7656 18300 7708 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 5724 18232 5776 18284
rect 6920 18232 6972 18284
rect 7288 18232 7340 18284
rect 4620 18164 4672 18216
rect 4896 18207 4948 18216
rect 4896 18173 4905 18207
rect 4905 18173 4939 18207
rect 4939 18173 4948 18207
rect 4896 18164 4948 18173
rect 7932 18232 7984 18284
rect 15292 18368 15344 18420
rect 9220 18232 9272 18284
rect 10876 18232 10928 18284
rect 10968 18275 11020 18284
rect 10968 18241 10977 18275
rect 10977 18241 11011 18275
rect 11011 18241 11020 18275
rect 11704 18275 11756 18284
rect 10968 18232 11020 18241
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 14556 18343 14608 18352
rect 14556 18309 14565 18343
rect 14565 18309 14599 18343
rect 14599 18309 14608 18343
rect 14556 18300 14608 18309
rect 16948 18300 17000 18352
rect 17408 18300 17460 18352
rect 22192 18343 22244 18352
rect 12164 18232 12216 18284
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 18420 18275 18472 18284
rect 12532 18232 12584 18241
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 18696 18232 18748 18284
rect 19616 18275 19668 18284
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 22192 18309 22201 18343
rect 22201 18309 22235 18343
rect 22235 18309 22244 18343
rect 22192 18300 22244 18309
rect 24860 18343 24912 18352
rect 24860 18309 24869 18343
rect 24869 18309 24903 18343
rect 24903 18309 24912 18343
rect 24860 18300 24912 18309
rect 26056 18343 26108 18352
rect 26056 18309 26065 18343
rect 26065 18309 26099 18343
rect 26099 18309 26108 18343
rect 26056 18300 26108 18309
rect 27252 18343 27304 18352
rect 27252 18309 27261 18343
rect 27261 18309 27295 18343
rect 27295 18309 27304 18343
rect 27252 18300 27304 18309
rect 21088 18232 21140 18284
rect 21456 18232 21508 18284
rect 23756 18275 23808 18284
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 28356 18275 28408 18284
rect 28356 18241 28365 18275
rect 28365 18241 28399 18275
rect 28399 18241 28408 18275
rect 28356 18232 28408 18241
rect 28540 18275 28592 18284
rect 28540 18241 28549 18275
rect 28549 18241 28583 18275
rect 28583 18241 28592 18275
rect 28540 18232 28592 18241
rect 13544 18207 13596 18216
rect 9864 18096 9916 18148
rect 6552 18028 6604 18080
rect 9680 18028 9732 18080
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 11428 18028 11480 18080
rect 12900 18096 12952 18148
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 16672 18164 16724 18216
rect 13360 18028 13412 18080
rect 14556 18096 14608 18148
rect 16212 18139 16264 18148
rect 16212 18105 16221 18139
rect 16221 18105 16255 18139
rect 16255 18105 16264 18139
rect 16212 18096 16264 18105
rect 16488 18096 16540 18148
rect 17316 18164 17368 18216
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 22100 18164 22152 18173
rect 23296 18164 23348 18216
rect 24860 18164 24912 18216
rect 26148 18164 26200 18216
rect 26608 18207 26660 18216
rect 26608 18173 26617 18207
rect 26617 18173 26651 18207
rect 26651 18173 26660 18207
rect 26608 18164 26660 18173
rect 27804 18139 27856 18148
rect 16764 18028 16816 18080
rect 18052 18028 18104 18080
rect 20444 18028 20496 18080
rect 23204 18028 23256 18080
rect 27804 18105 27813 18139
rect 27813 18105 27847 18139
rect 27847 18105 27856 18139
rect 27804 18096 27856 18105
rect 26240 18028 26292 18080
rect 29000 18071 29052 18080
rect 29000 18037 29009 18071
rect 29009 18037 29043 18071
rect 29043 18037 29052 18071
rect 29000 18028 29052 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 6736 17824 6788 17876
rect 9404 17824 9456 17876
rect 10876 17824 10928 17876
rect 11796 17824 11848 17876
rect 14372 17824 14424 17876
rect 15108 17824 15160 17876
rect 16212 17824 16264 17876
rect 19432 17824 19484 17876
rect 22192 17824 22244 17876
rect 26056 17824 26108 17876
rect 32128 17867 32180 17876
rect 32128 17833 32137 17867
rect 32137 17833 32171 17867
rect 32171 17833 32180 17867
rect 32128 17824 32180 17833
rect 4620 17688 4672 17740
rect 7472 17756 7524 17808
rect 8576 17756 8628 17808
rect 10416 17756 10468 17808
rect 10692 17756 10744 17808
rect 13268 17756 13320 17808
rect 15660 17799 15712 17808
rect 15660 17765 15669 17799
rect 15669 17765 15703 17799
rect 15703 17765 15712 17799
rect 15660 17756 15712 17765
rect 1860 17552 1912 17604
rect 6644 17688 6696 17740
rect 6828 17688 6880 17740
rect 7564 17688 7616 17740
rect 9956 17688 10008 17740
rect 10324 17731 10376 17740
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 20812 17756 20864 17808
rect 22100 17688 22152 17740
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 26240 17731 26292 17740
rect 26240 17697 26249 17731
rect 26249 17697 26283 17731
rect 26283 17697 26292 17731
rect 26240 17688 26292 17697
rect 29092 17688 29144 17740
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 6736 17620 6788 17672
rect 8668 17620 8720 17672
rect 11612 17620 11664 17672
rect 11980 17620 12032 17672
rect 12348 17663 12400 17672
rect 12348 17629 12357 17663
rect 12357 17629 12391 17663
rect 12391 17629 12400 17663
rect 12348 17620 12400 17629
rect 13820 17620 13872 17672
rect 14188 17620 14240 17672
rect 14648 17620 14700 17672
rect 17132 17620 17184 17672
rect 18512 17663 18564 17672
rect 18512 17629 18521 17663
rect 18521 17629 18555 17663
rect 18555 17629 18564 17663
rect 18512 17620 18564 17629
rect 19524 17663 19576 17672
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 19616 17620 19668 17672
rect 25780 17620 25832 17672
rect 27712 17663 27764 17672
rect 27712 17629 27721 17663
rect 27721 17629 27755 17663
rect 27755 17629 27764 17663
rect 27712 17620 27764 17629
rect 29184 17620 29236 17672
rect 6092 17552 6144 17604
rect 9772 17595 9824 17604
rect 9772 17561 9781 17595
rect 9781 17561 9815 17595
rect 9815 17561 9824 17595
rect 9772 17552 9824 17561
rect 10968 17552 11020 17604
rect 13268 17552 13320 17604
rect 15108 17595 15160 17604
rect 15108 17561 15117 17595
rect 15117 17561 15151 17595
rect 15151 17561 15160 17595
rect 15108 17552 15160 17561
rect 17500 17595 17552 17604
rect 5908 17484 5960 17536
rect 8392 17484 8444 17536
rect 10692 17484 10744 17536
rect 12532 17484 12584 17536
rect 14832 17484 14884 17536
rect 17500 17561 17509 17595
rect 17509 17561 17543 17595
rect 17543 17561 17552 17595
rect 17500 17552 17552 17561
rect 17592 17552 17644 17604
rect 18236 17552 18288 17604
rect 19156 17552 19208 17604
rect 23204 17552 23256 17604
rect 26332 17595 26384 17604
rect 26332 17561 26341 17595
rect 26341 17561 26375 17595
rect 26375 17561 26384 17595
rect 26332 17552 26384 17561
rect 27160 17552 27212 17604
rect 37280 17620 37332 17672
rect 16396 17484 16448 17536
rect 17408 17484 17460 17536
rect 19984 17484 20036 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 27896 17484 27948 17536
rect 29276 17484 29328 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 3700 17144 3752 17196
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 8576 17280 8628 17332
rect 7196 17212 7248 17264
rect 8024 17212 8076 17264
rect 8484 17144 8536 17196
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 9404 17212 9456 17264
rect 10508 17212 10560 17264
rect 10692 17212 10744 17264
rect 15108 17280 15160 17332
rect 11428 17212 11480 17264
rect 16304 17212 16356 17264
rect 11980 17187 12032 17196
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 6736 17076 6788 17128
rect 7564 17076 7616 17128
rect 10140 17076 10192 17128
rect 6828 17008 6880 17060
rect 10048 17008 10100 17060
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 13268 17187 13320 17196
rect 11244 17076 11296 17128
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 17224 17187 17276 17196
rect 17224 17153 17233 17187
rect 17233 17153 17267 17187
rect 17267 17153 17276 17187
rect 17224 17144 17276 17153
rect 13728 17076 13780 17128
rect 14556 17119 14608 17128
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 15660 17119 15712 17128
rect 15660 17085 15669 17119
rect 15669 17085 15703 17119
rect 15703 17085 15712 17119
rect 15660 17076 15712 17085
rect 19156 17280 19208 17332
rect 20260 17280 20312 17332
rect 22744 17280 22796 17332
rect 25044 17280 25096 17332
rect 18052 17255 18104 17264
rect 18052 17221 18061 17255
rect 18061 17221 18095 17255
rect 18095 17221 18104 17255
rect 18052 17212 18104 17221
rect 19248 17255 19300 17264
rect 19248 17221 19257 17255
rect 19257 17221 19291 17255
rect 19291 17221 19300 17255
rect 19248 17212 19300 17221
rect 20444 17255 20496 17264
rect 20444 17221 20453 17255
rect 20453 17221 20487 17255
rect 20487 17221 20496 17255
rect 20444 17212 20496 17221
rect 23388 17255 23440 17264
rect 23388 17221 23397 17255
rect 23397 17221 23431 17255
rect 23431 17221 23440 17255
rect 23388 17212 23440 17221
rect 25504 17212 25556 17264
rect 25964 17255 26016 17264
rect 25964 17221 25973 17255
rect 25973 17221 26007 17255
rect 26007 17221 26016 17255
rect 25964 17212 26016 17221
rect 26056 17255 26108 17264
rect 26056 17221 26065 17255
rect 26065 17221 26099 17255
rect 26099 17221 26108 17255
rect 27896 17255 27948 17264
rect 26056 17212 26108 17221
rect 27896 17221 27905 17255
rect 27905 17221 27939 17255
rect 27939 17221 27948 17255
rect 27896 17212 27948 17221
rect 29092 17212 29144 17264
rect 18972 17076 19024 17128
rect 19800 17076 19852 17128
rect 21272 17076 21324 17128
rect 24216 17076 24268 17128
rect 24584 17144 24636 17196
rect 29276 17187 29328 17196
rect 29276 17153 29285 17187
rect 29285 17153 29319 17187
rect 29319 17153 29328 17187
rect 29276 17144 29328 17153
rect 38292 17187 38344 17196
rect 38292 17153 38301 17187
rect 38301 17153 38335 17187
rect 38335 17153 38344 17187
rect 38292 17144 38344 17153
rect 24860 17076 24912 17128
rect 26608 17119 26660 17128
rect 26608 17085 26617 17119
rect 26617 17085 26651 17119
rect 26651 17085 26660 17119
rect 26608 17076 26660 17085
rect 27068 17076 27120 17128
rect 3332 16940 3384 16992
rect 4712 16940 4764 16992
rect 5448 16940 5500 16992
rect 9956 16940 10008 16992
rect 13728 16940 13780 16992
rect 15108 17008 15160 17060
rect 19432 17008 19484 17060
rect 20168 17008 20220 17060
rect 29828 17076 29880 17128
rect 30196 17076 30248 17128
rect 29000 17008 29052 17060
rect 15200 16940 15252 16992
rect 16580 16940 16632 16992
rect 17592 16940 17644 16992
rect 19892 16940 19944 16992
rect 22192 16940 22244 16992
rect 38108 16983 38160 16992
rect 38108 16949 38117 16983
rect 38117 16949 38151 16983
rect 38151 16949 38160 16983
rect 38108 16940 38160 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5816 16736 5868 16788
rect 7932 16736 7984 16788
rect 2688 16532 2740 16584
rect 4804 16532 4856 16584
rect 6368 16668 6420 16720
rect 5724 16600 5776 16652
rect 6552 16600 6604 16652
rect 7564 16600 7616 16652
rect 8116 16600 8168 16652
rect 8208 16532 8260 16584
rect 13268 16736 13320 16788
rect 8484 16668 8536 16720
rect 8576 16600 8628 16652
rect 9404 16600 9456 16652
rect 10324 16668 10376 16720
rect 11336 16668 11388 16720
rect 13912 16736 13964 16788
rect 17592 16736 17644 16788
rect 19248 16736 19300 16788
rect 19800 16779 19852 16788
rect 19800 16745 19809 16779
rect 19809 16745 19843 16779
rect 19843 16745 19852 16779
rect 19800 16736 19852 16745
rect 19892 16736 19944 16788
rect 22284 16736 22336 16788
rect 26056 16736 26108 16788
rect 10600 16532 10652 16584
rect 11060 16600 11112 16652
rect 11796 16643 11848 16652
rect 11796 16609 11805 16643
rect 11805 16609 11839 16643
rect 11839 16609 11848 16643
rect 11796 16600 11848 16609
rect 14372 16668 14424 16720
rect 11244 16532 11296 16584
rect 14464 16600 14516 16652
rect 16028 16668 16080 16720
rect 16672 16600 16724 16652
rect 17132 16532 17184 16584
rect 18512 16668 18564 16720
rect 18972 16668 19024 16720
rect 21732 16668 21784 16720
rect 17592 16532 17644 16584
rect 9404 16464 9456 16516
rect 2780 16396 2832 16448
rect 2872 16396 2924 16448
rect 3424 16396 3476 16448
rect 5080 16396 5132 16448
rect 6276 16396 6328 16448
rect 8300 16396 8352 16448
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 9128 16396 9180 16448
rect 9864 16464 9916 16516
rect 12716 16464 12768 16516
rect 15568 16464 15620 16516
rect 16488 16464 16540 16516
rect 17960 16464 18012 16516
rect 10876 16439 10928 16448
rect 10876 16405 10885 16439
rect 10885 16405 10919 16439
rect 10919 16405 10928 16439
rect 10876 16396 10928 16405
rect 11704 16396 11756 16448
rect 13268 16396 13320 16448
rect 14832 16396 14884 16448
rect 17040 16396 17092 16448
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 20076 16600 20128 16652
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 20812 16643 20864 16652
rect 20812 16609 20821 16643
rect 20821 16609 20855 16643
rect 20855 16609 20864 16643
rect 20812 16600 20864 16609
rect 20904 16600 20956 16652
rect 22652 16532 22704 16584
rect 27160 16575 27212 16584
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 38108 16600 38160 16652
rect 20628 16507 20680 16516
rect 20628 16473 20637 16507
rect 20637 16473 20671 16507
rect 20671 16473 20680 16507
rect 21732 16507 21784 16516
rect 20628 16464 20680 16473
rect 21732 16473 21741 16507
rect 21741 16473 21775 16507
rect 21775 16473 21784 16507
rect 21732 16464 21784 16473
rect 22192 16464 22244 16516
rect 22376 16507 22428 16516
rect 22376 16473 22385 16507
rect 22385 16473 22419 16507
rect 22419 16473 22428 16507
rect 22376 16464 22428 16473
rect 22468 16464 22520 16516
rect 22100 16396 22152 16448
rect 22836 16439 22888 16448
rect 22836 16405 22845 16439
rect 22845 16405 22879 16439
rect 22879 16405 22888 16439
rect 22836 16396 22888 16405
rect 24492 16396 24544 16448
rect 27252 16439 27304 16448
rect 27252 16405 27261 16439
rect 27261 16405 27295 16439
rect 27295 16405 27304 16439
rect 27252 16396 27304 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 7380 16192 7432 16244
rect 8392 16192 8444 16244
rect 8484 16192 8536 16244
rect 4068 16124 4120 16176
rect 5448 16167 5500 16176
rect 5448 16133 5457 16167
rect 5457 16133 5491 16167
rect 5491 16133 5500 16167
rect 5448 16124 5500 16133
rect 6276 16124 6328 16176
rect 9036 16124 9088 16176
rect 9128 16124 9180 16176
rect 10048 16124 10100 16176
rect 12072 16124 12124 16176
rect 15292 16192 15344 16244
rect 15752 16192 15804 16244
rect 17500 16192 17552 16244
rect 22100 16192 22152 16244
rect 23296 16192 23348 16244
rect 23388 16192 23440 16244
rect 27252 16192 27304 16244
rect 15936 16124 15988 16176
rect 19248 16124 19300 16176
rect 20352 16167 20404 16176
rect 20352 16133 20361 16167
rect 20361 16133 20395 16167
rect 20395 16133 20404 16167
rect 20352 16124 20404 16133
rect 20444 16124 20496 16176
rect 20628 16124 20680 16176
rect 22836 16167 22888 16176
rect 22836 16133 22845 16167
rect 22845 16133 22879 16167
rect 22879 16133 22888 16167
rect 22836 16124 22888 16133
rect 22928 16167 22980 16176
rect 22928 16133 22937 16167
rect 22937 16133 22971 16167
rect 22971 16133 22980 16167
rect 24492 16167 24544 16176
rect 22928 16124 22980 16133
rect 24492 16133 24501 16167
rect 24501 16133 24535 16167
rect 24535 16133 24544 16167
rect 24492 16124 24544 16133
rect 26056 16167 26108 16176
rect 26056 16133 26065 16167
rect 26065 16133 26099 16167
rect 26099 16133 26108 16167
rect 26056 16124 26108 16133
rect 27804 16124 27856 16176
rect 3976 16099 4028 16108
rect 3976 16065 3985 16099
rect 3985 16065 4019 16099
rect 4019 16065 4028 16099
rect 3976 16056 4028 16065
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 6920 16056 6972 16065
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8208 16099 8260 16108
rect 8208 16065 8217 16099
rect 8217 16065 8251 16099
rect 8251 16065 8260 16099
rect 8208 16056 8260 16065
rect 3700 15988 3752 16040
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6092 15988 6144 16040
rect 7104 15988 7156 16040
rect 9128 15988 9180 16040
rect 10692 16056 10744 16108
rect 9680 15988 9732 16040
rect 11060 15988 11112 16040
rect 12440 16056 12492 16108
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 16212 16056 16264 16108
rect 17316 16056 17368 16108
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 18236 16056 18288 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 22652 16056 22704 16108
rect 38292 16099 38344 16108
rect 13176 15988 13228 16040
rect 14188 16031 14240 16040
rect 14188 15997 14197 16031
rect 14197 15997 14231 16031
rect 14231 15997 14240 16031
rect 14188 15988 14240 15997
rect 2228 15920 2280 15972
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 3056 15852 3108 15904
rect 4896 15852 4948 15904
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 8576 15852 8628 15904
rect 8944 15895 8996 15904
rect 8944 15861 8953 15895
rect 8953 15861 8987 15895
rect 8987 15861 8996 15895
rect 8944 15852 8996 15861
rect 9772 15920 9824 15972
rect 16764 15920 16816 15972
rect 17868 15988 17920 16040
rect 18052 15988 18104 16040
rect 17776 15920 17828 15972
rect 21272 15988 21324 16040
rect 21364 15988 21416 16040
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 23112 15988 23164 15997
rect 24400 16031 24452 16040
rect 24400 15997 24409 16031
rect 24409 15997 24443 16031
rect 24443 15997 24452 16031
rect 24400 15988 24452 15997
rect 18972 15920 19024 15972
rect 23388 15920 23440 15972
rect 12164 15852 12216 15904
rect 12808 15852 12860 15904
rect 13636 15852 13688 15904
rect 14188 15852 14240 15904
rect 17592 15852 17644 15904
rect 17868 15852 17920 15904
rect 19432 15852 19484 15904
rect 22376 15852 22428 15904
rect 24124 15852 24176 15904
rect 38292 16065 38301 16099
rect 38301 16065 38335 16099
rect 38335 16065 38344 16099
rect 38292 16056 38344 16065
rect 26148 15988 26200 16040
rect 29644 15920 29696 15972
rect 25964 15852 26016 15904
rect 29000 15852 29052 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 4988 15648 5040 15700
rect 7012 15648 7064 15700
rect 9864 15648 9916 15700
rect 11060 15648 11112 15700
rect 3976 15580 4028 15632
rect 7288 15580 7340 15632
rect 7564 15580 7616 15632
rect 9128 15580 9180 15632
rect 9496 15580 9548 15632
rect 10692 15580 10744 15632
rect 10876 15580 10928 15632
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 2688 15444 2740 15496
rect 4620 15512 4672 15564
rect 6460 15555 6512 15564
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 4804 15444 4856 15496
rect 5080 15419 5132 15428
rect 5080 15385 5089 15419
rect 5089 15385 5123 15419
rect 5123 15385 5132 15419
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 7104 15444 7156 15496
rect 8576 15444 8628 15496
rect 5080 15376 5132 15385
rect 7380 15376 7432 15428
rect 7840 15419 7892 15428
rect 7840 15385 7849 15419
rect 7849 15385 7883 15419
rect 7883 15385 7892 15419
rect 7840 15376 7892 15385
rect 9772 15419 9824 15428
rect 3240 15308 3292 15360
rect 4344 15351 4396 15360
rect 4344 15317 4353 15351
rect 4353 15317 4387 15351
rect 4387 15317 4396 15351
rect 4344 15308 4396 15317
rect 7012 15308 7064 15360
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 9772 15385 9781 15419
rect 9781 15385 9815 15419
rect 9815 15385 9824 15419
rect 9772 15376 9824 15385
rect 9956 15376 10008 15428
rect 11888 15512 11940 15564
rect 12348 15580 12400 15632
rect 15660 15648 15712 15700
rect 16764 15691 16816 15700
rect 16764 15657 16773 15691
rect 16773 15657 16807 15691
rect 16807 15657 16816 15691
rect 16764 15648 16816 15657
rect 18788 15648 18840 15700
rect 22928 15648 22980 15700
rect 23020 15648 23072 15700
rect 24400 15648 24452 15700
rect 11612 15444 11664 15496
rect 11428 15376 11480 15428
rect 12164 15419 12216 15428
rect 12164 15385 12173 15419
rect 12173 15385 12207 15419
rect 12207 15385 12216 15419
rect 13728 15580 13780 15632
rect 15568 15580 15620 15632
rect 22376 15580 22428 15632
rect 23112 15580 23164 15632
rect 13268 15512 13320 15564
rect 15384 15555 15436 15564
rect 15384 15521 15393 15555
rect 15393 15521 15427 15555
rect 15427 15521 15436 15555
rect 15384 15512 15436 15521
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16856 15512 16908 15564
rect 18144 15512 18196 15564
rect 20904 15512 20956 15564
rect 22744 15555 22796 15564
rect 22744 15521 22753 15555
rect 22753 15521 22787 15555
rect 22787 15521 22796 15555
rect 22744 15512 22796 15521
rect 23664 15512 23716 15564
rect 29828 15555 29880 15564
rect 14280 15444 14332 15496
rect 20444 15444 20496 15496
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 12164 15376 12216 15385
rect 17868 15419 17920 15428
rect 17868 15385 17877 15419
rect 17877 15385 17911 15419
rect 17911 15385 17920 15419
rect 17868 15376 17920 15385
rect 19984 15376 20036 15428
rect 23388 15487 23440 15496
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 23848 15487 23900 15496
rect 23388 15444 23440 15453
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 36360 15512 36412 15564
rect 37740 15555 37792 15564
rect 37740 15521 37749 15555
rect 37749 15521 37783 15555
rect 37783 15521 37792 15555
rect 37740 15512 37792 15521
rect 24768 15444 24820 15496
rect 24860 15444 24912 15496
rect 29000 15487 29052 15496
rect 29000 15453 29009 15487
rect 29009 15453 29043 15487
rect 29043 15453 29052 15487
rect 29000 15444 29052 15453
rect 37188 15444 37240 15496
rect 8484 15308 8536 15317
rect 10048 15308 10100 15360
rect 10324 15308 10376 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 20076 15308 20128 15360
rect 29920 15419 29972 15428
rect 29920 15385 29929 15419
rect 29929 15385 29963 15419
rect 29963 15385 29972 15419
rect 29920 15376 29972 15385
rect 23940 15351 23992 15360
rect 23940 15317 23949 15351
rect 23949 15317 23983 15351
rect 23983 15317 23992 15351
rect 23940 15308 23992 15317
rect 24032 15308 24084 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2412 14968 2464 15020
rect 4252 15036 4304 15088
rect 3792 14968 3844 15020
rect 6276 15036 6328 15088
rect 5816 15011 5868 15020
rect 3608 14900 3660 14952
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 4988 14832 5040 14884
rect 7288 15036 7340 15088
rect 8024 15036 8076 15088
rect 7840 14968 7892 15020
rect 9496 15104 9548 15156
rect 8300 15036 8352 15088
rect 8944 14968 8996 15020
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 11244 14968 11296 15020
rect 12440 15036 12492 15088
rect 12992 15036 13044 15088
rect 13360 15079 13412 15088
rect 13360 15045 13369 15079
rect 13369 15045 13403 15079
rect 13403 15045 13412 15079
rect 13360 15036 13412 15045
rect 13912 15079 13964 15088
rect 13912 15045 13921 15079
rect 13921 15045 13955 15079
rect 13955 15045 13964 15079
rect 13912 15036 13964 15045
rect 15660 15104 15712 15156
rect 17408 15079 17460 15088
rect 17408 15045 17417 15079
rect 17417 15045 17451 15079
rect 17451 15045 17460 15079
rect 17408 15036 17460 15045
rect 18604 15079 18656 15088
rect 18604 15045 18613 15079
rect 18613 15045 18647 15079
rect 18647 15045 18656 15079
rect 18604 15036 18656 15045
rect 19524 15104 19576 15156
rect 20168 15104 20220 15156
rect 20260 15104 20312 15156
rect 7380 14900 7432 14952
rect 8392 14832 8444 14884
rect 11796 14900 11848 14952
rect 13360 14900 13412 14952
rect 16396 14968 16448 15020
rect 19248 14968 19300 15020
rect 19800 14968 19852 15020
rect 20444 14968 20496 15020
rect 23572 15104 23624 15156
rect 21180 15036 21232 15088
rect 22468 15036 22520 15088
rect 26240 15104 26292 15156
rect 27620 15104 27672 15156
rect 24032 15036 24084 15088
rect 24768 15036 24820 15088
rect 28264 15011 28316 15020
rect 16488 14900 16540 14952
rect 16672 14900 16724 14952
rect 17592 14943 17644 14952
rect 17592 14909 17601 14943
rect 17601 14909 17635 14943
rect 17635 14909 17644 14943
rect 17592 14900 17644 14909
rect 17684 14900 17736 14952
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 21916 14900 21968 14952
rect 23020 14900 23072 14952
rect 23296 14900 23348 14952
rect 2596 14764 2648 14816
rect 2964 14764 3016 14816
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5632 14764 5684 14816
rect 6920 14764 6972 14816
rect 7104 14764 7156 14816
rect 8208 14764 8260 14816
rect 9404 14764 9456 14816
rect 12992 14832 13044 14884
rect 20168 14832 20220 14884
rect 12716 14764 12768 14816
rect 12808 14764 12860 14816
rect 14004 14764 14056 14816
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 16856 14764 16908 14816
rect 17316 14764 17368 14816
rect 17684 14764 17736 14816
rect 19800 14764 19852 14816
rect 21088 14764 21140 14816
rect 21272 14832 21324 14884
rect 22376 14832 22428 14884
rect 24676 14900 24728 14952
rect 28264 14977 28273 15011
rect 28273 14977 28307 15011
rect 28307 14977 28316 15011
rect 28264 14968 28316 14977
rect 38016 15011 38068 15020
rect 38016 14977 38025 15011
rect 38025 14977 38059 15011
rect 38059 14977 38068 15011
rect 38016 14968 38068 14977
rect 28356 14900 28408 14952
rect 30012 14900 30064 14952
rect 22744 14764 22796 14816
rect 27252 14764 27304 14816
rect 30196 14764 30248 14816
rect 37924 14764 37976 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4528 14560 4580 14612
rect 8484 14560 8536 14612
rect 6920 14492 6972 14544
rect 8392 14492 8444 14544
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 4620 14424 4672 14476
rect 9220 14424 9272 14476
rect 12716 14560 12768 14612
rect 14188 14560 14240 14612
rect 2504 14356 2556 14408
rect 6276 14356 6328 14408
rect 7288 14356 7340 14408
rect 8392 14399 8444 14408
rect 2872 14331 2924 14340
rect 2872 14297 2881 14331
rect 2881 14297 2915 14331
rect 2915 14297 2924 14331
rect 2872 14288 2924 14297
rect 3516 14288 3568 14340
rect 4712 14288 4764 14340
rect 5448 14331 5500 14340
rect 5448 14297 5457 14331
rect 5457 14297 5491 14331
rect 5491 14297 5500 14331
rect 5448 14288 5500 14297
rect 7656 14288 7708 14340
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 8852 14356 8904 14408
rect 11612 14492 11664 14544
rect 13728 14492 13780 14544
rect 17408 14560 17460 14612
rect 17776 14560 17828 14612
rect 20720 14560 20772 14612
rect 26056 14560 26108 14612
rect 26240 14603 26292 14612
rect 26240 14569 26249 14603
rect 26249 14569 26283 14603
rect 26283 14569 26292 14603
rect 26240 14560 26292 14569
rect 26608 14560 26660 14612
rect 27712 14560 27764 14612
rect 38016 14560 38068 14612
rect 16304 14492 16356 14544
rect 22100 14492 22152 14544
rect 22192 14492 22244 14544
rect 10232 14424 10284 14476
rect 12072 14424 12124 14476
rect 13176 14424 13228 14476
rect 14556 14424 14608 14476
rect 16488 14424 16540 14476
rect 16764 14424 16816 14476
rect 17776 14467 17828 14476
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 20352 14424 20404 14476
rect 21916 14424 21968 14476
rect 23480 14467 23532 14476
rect 23480 14433 23489 14467
rect 23489 14433 23523 14467
rect 23523 14433 23532 14467
rect 23480 14424 23532 14433
rect 8576 14288 8628 14340
rect 17316 14356 17368 14408
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 29368 14492 29420 14544
rect 30012 14467 30064 14476
rect 25228 14399 25280 14408
rect 25228 14365 25237 14399
rect 25237 14365 25271 14399
rect 25271 14365 25280 14399
rect 25228 14356 25280 14365
rect 25596 14356 25648 14408
rect 27252 14399 27304 14408
rect 27252 14365 27261 14399
rect 27261 14365 27295 14399
rect 27295 14365 27304 14399
rect 27252 14356 27304 14365
rect 27712 14399 27764 14408
rect 27712 14365 27721 14399
rect 27721 14365 27755 14399
rect 27755 14365 27764 14399
rect 27712 14356 27764 14365
rect 28356 14399 28408 14408
rect 28356 14365 28365 14399
rect 28365 14365 28399 14399
rect 28399 14365 28408 14399
rect 28356 14356 28408 14365
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 8024 14220 8076 14272
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 10692 14220 10744 14272
rect 10876 14331 10928 14340
rect 10876 14297 10885 14331
rect 10885 14297 10919 14331
rect 10919 14297 10928 14331
rect 10876 14288 10928 14297
rect 11244 14288 11296 14340
rect 12348 14288 12400 14340
rect 13728 14331 13780 14340
rect 11152 14220 11204 14272
rect 13728 14297 13737 14331
rect 13737 14297 13771 14331
rect 13771 14297 13780 14331
rect 13728 14288 13780 14297
rect 14832 14288 14884 14340
rect 15660 14331 15712 14340
rect 15660 14297 15669 14331
rect 15669 14297 15703 14331
rect 15703 14297 15712 14331
rect 15660 14288 15712 14297
rect 16396 14331 16448 14340
rect 16396 14297 16405 14331
rect 16405 14297 16439 14331
rect 16439 14297 16448 14331
rect 16396 14288 16448 14297
rect 16488 14288 16540 14340
rect 19248 14288 19300 14340
rect 19524 14331 19576 14340
rect 19524 14297 19533 14331
rect 19533 14297 19567 14331
rect 19567 14297 19576 14331
rect 19524 14288 19576 14297
rect 22836 14331 22888 14340
rect 13084 14220 13136 14272
rect 13452 14220 13504 14272
rect 15752 14220 15804 14272
rect 18972 14220 19024 14272
rect 19432 14220 19484 14272
rect 22836 14297 22845 14331
rect 22845 14297 22879 14331
rect 22879 14297 22888 14331
rect 22836 14288 22888 14297
rect 19984 14220 20036 14272
rect 22008 14220 22060 14272
rect 27344 14288 27396 14340
rect 30012 14433 30021 14467
rect 30021 14433 30055 14467
rect 30055 14433 30064 14467
rect 30012 14424 30064 14433
rect 30196 14467 30248 14476
rect 30196 14433 30205 14467
rect 30205 14433 30239 14467
rect 30239 14433 30248 14467
rect 30196 14424 30248 14433
rect 38200 14288 38252 14340
rect 25320 14263 25372 14272
rect 25320 14229 25329 14263
rect 25329 14229 25363 14263
rect 25363 14229 25372 14263
rect 25320 14220 25372 14229
rect 27712 14220 27764 14272
rect 28172 14220 28224 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4804 14016 4856 14068
rect 8300 14016 8352 14068
rect 3056 13948 3108 14000
rect 3332 13991 3384 14000
rect 3332 13957 3341 13991
rect 3341 13957 3375 13991
rect 3375 13957 3384 13991
rect 3332 13948 3384 13957
rect 5264 13948 5316 14000
rect 7288 13991 7340 14000
rect 7288 13957 7297 13991
rect 7297 13957 7331 13991
rect 7331 13957 7340 13991
rect 7288 13948 7340 13957
rect 7656 13948 7708 14000
rect 12072 14016 12124 14068
rect 2688 13880 2740 13932
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4712 13880 4764 13932
rect 4896 13880 4948 13932
rect 5448 13880 5500 13932
rect 5540 13880 5592 13932
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 7840 13880 7892 13889
rect 8300 13880 8352 13932
rect 10140 13948 10192 14000
rect 15108 14016 15160 14068
rect 15660 14016 15712 14068
rect 12532 13991 12584 14000
rect 12532 13957 12541 13991
rect 12541 13957 12575 13991
rect 12575 13957 12584 13991
rect 12532 13948 12584 13957
rect 13452 13948 13504 14000
rect 14188 13991 14240 14000
rect 14188 13957 14197 13991
rect 14197 13957 14231 13991
rect 14231 13957 14240 13991
rect 14188 13948 14240 13957
rect 14648 13948 14700 14000
rect 15752 13991 15804 14000
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 3884 13812 3936 13864
rect 5080 13812 5132 13864
rect 7012 13812 7064 13864
rect 8852 13812 8904 13864
rect 9956 13880 10008 13932
rect 11060 13855 11112 13864
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 3976 13676 4028 13728
rect 4896 13676 4948 13728
rect 5172 13676 5224 13728
rect 5356 13676 5408 13728
rect 6460 13744 6512 13796
rect 6000 13676 6052 13728
rect 7012 13676 7064 13728
rect 8576 13676 8628 13728
rect 9036 13676 9088 13728
rect 11060 13821 11069 13855
rect 11069 13821 11103 13855
rect 11103 13821 11112 13855
rect 11060 13812 11112 13821
rect 12164 13880 12216 13932
rect 13912 13880 13964 13932
rect 12992 13744 13044 13796
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 15200 13880 15252 13932
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 15752 13948 15804 13957
rect 16304 13991 16356 14000
rect 16304 13957 16313 13991
rect 16313 13957 16347 13991
rect 16347 13957 16356 13991
rect 16304 13948 16356 13957
rect 17040 13991 17092 14000
rect 17040 13957 17049 13991
rect 17049 13957 17083 13991
rect 17083 13957 17092 13991
rect 17040 13948 17092 13957
rect 19156 14016 19208 14068
rect 20260 14016 20312 14068
rect 29920 14016 29972 14068
rect 17776 13948 17828 14000
rect 19248 13948 19300 14000
rect 21088 13948 21140 14000
rect 22100 13948 22152 14000
rect 23112 13948 23164 14000
rect 25320 13948 25372 14000
rect 27344 13991 27396 14000
rect 27344 13957 27353 13991
rect 27353 13957 27387 13991
rect 27387 13957 27396 13991
rect 27344 13948 27396 13957
rect 27712 13948 27764 14000
rect 18144 13923 18196 13932
rect 15384 13812 15436 13864
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13880 18196 13889
rect 15844 13812 15896 13864
rect 16672 13744 16724 13796
rect 19248 13812 19300 13864
rect 19340 13812 19392 13864
rect 20628 13812 20680 13864
rect 21364 13855 21416 13864
rect 21364 13821 21373 13855
rect 21373 13821 21407 13855
rect 21407 13821 21416 13855
rect 21364 13812 21416 13821
rect 22836 13812 22888 13864
rect 20352 13744 20404 13796
rect 20720 13744 20772 13796
rect 23388 13812 23440 13864
rect 24308 13855 24360 13864
rect 24308 13821 24317 13855
rect 24317 13821 24351 13855
rect 24351 13821 24360 13855
rect 24308 13812 24360 13821
rect 24400 13812 24452 13864
rect 27896 13923 27948 13932
rect 27896 13889 27905 13923
rect 27905 13889 27939 13923
rect 27939 13889 27948 13923
rect 27896 13880 27948 13889
rect 37280 13880 37332 13932
rect 27252 13855 27304 13864
rect 24584 13744 24636 13796
rect 10140 13676 10192 13728
rect 11336 13676 11388 13728
rect 13728 13676 13780 13728
rect 18696 13676 18748 13728
rect 20168 13676 20220 13728
rect 21916 13676 21968 13728
rect 22100 13719 22152 13728
rect 22100 13685 22109 13719
rect 22109 13685 22143 13719
rect 22143 13685 22152 13719
rect 22100 13676 22152 13685
rect 23112 13676 23164 13728
rect 24308 13676 24360 13728
rect 27252 13821 27261 13855
rect 27261 13821 27295 13855
rect 27295 13821 27304 13855
rect 27252 13812 27304 13821
rect 29368 13855 29420 13864
rect 29368 13821 29377 13855
rect 29377 13821 29411 13855
rect 29411 13821 29420 13855
rect 29368 13812 29420 13821
rect 29644 13855 29696 13864
rect 29644 13821 29653 13855
rect 29653 13821 29687 13855
rect 29687 13821 29696 13855
rect 29644 13812 29696 13821
rect 37188 13812 37240 13864
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 3792 13472 3844 13524
rect 6000 13472 6052 13524
rect 6184 13472 6236 13524
rect 7288 13472 7340 13524
rect 8760 13472 8812 13524
rect 9128 13472 9180 13524
rect 12716 13472 12768 13524
rect 12808 13472 12860 13524
rect 14372 13472 14424 13524
rect 15384 13472 15436 13524
rect 16120 13472 16172 13524
rect 16304 13472 16356 13524
rect 16672 13472 16724 13524
rect 11244 13404 11296 13456
rect 6920 13336 6972 13388
rect 7288 13379 7340 13388
rect 7288 13345 7297 13379
rect 7297 13345 7331 13379
rect 7331 13345 7340 13379
rect 7288 13336 7340 13345
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 15936 13404 15988 13456
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 1952 13243 2004 13252
rect 1952 13209 1961 13243
rect 1961 13209 1995 13243
rect 1995 13209 2004 13243
rect 5540 13268 5592 13320
rect 5632 13268 5684 13320
rect 6184 13268 6236 13320
rect 1952 13200 2004 13209
rect 5172 13132 5224 13184
rect 5816 13200 5868 13252
rect 6828 13243 6880 13252
rect 6828 13209 6837 13243
rect 6837 13209 6871 13243
rect 6871 13209 6880 13243
rect 6828 13200 6880 13209
rect 7012 13200 7064 13252
rect 8300 13200 8352 13252
rect 11060 13268 11112 13320
rect 17316 13336 17368 13388
rect 19156 13404 19208 13456
rect 21456 13472 21508 13524
rect 25044 13472 25096 13524
rect 9588 13200 9640 13252
rect 9772 13200 9824 13252
rect 11152 13200 11204 13252
rect 11520 13243 11572 13252
rect 11520 13209 11529 13243
rect 11529 13209 11563 13243
rect 11563 13209 11572 13243
rect 11520 13200 11572 13209
rect 12532 13200 12584 13252
rect 14372 13243 14424 13252
rect 14372 13209 14381 13243
rect 14381 13209 14415 13243
rect 14415 13209 14424 13243
rect 14372 13200 14424 13209
rect 14464 13243 14516 13252
rect 14464 13209 14473 13243
rect 14473 13209 14507 13243
rect 14507 13209 14516 13243
rect 14464 13200 14516 13209
rect 15200 13200 15252 13252
rect 8116 13132 8168 13184
rect 8392 13132 8444 13184
rect 9220 13132 9272 13184
rect 12348 13132 12400 13184
rect 12808 13132 12860 13184
rect 14004 13132 14056 13184
rect 15844 13200 15896 13252
rect 16580 13200 16632 13252
rect 17408 13200 17460 13252
rect 20812 13336 20864 13388
rect 16488 13132 16540 13184
rect 17040 13132 17092 13184
rect 17868 13243 17920 13252
rect 17868 13209 17877 13243
rect 17877 13209 17911 13243
rect 17911 13209 17920 13243
rect 17868 13200 17920 13209
rect 18328 13200 18380 13252
rect 19432 13200 19484 13252
rect 19800 13243 19852 13252
rect 19800 13209 19809 13243
rect 19809 13209 19843 13243
rect 19843 13209 19852 13243
rect 19800 13200 19852 13209
rect 20168 13200 20220 13252
rect 20720 13243 20772 13252
rect 20720 13209 20729 13243
rect 20729 13209 20763 13243
rect 20763 13209 20772 13243
rect 27988 13404 28040 13456
rect 21364 13268 21416 13320
rect 21916 13268 21968 13320
rect 25872 13336 25924 13388
rect 25964 13336 26016 13388
rect 22652 13268 22704 13320
rect 22836 13268 22888 13320
rect 23388 13268 23440 13320
rect 23756 13311 23808 13320
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 20720 13200 20772 13209
rect 24308 13200 24360 13252
rect 25688 13243 25740 13252
rect 18512 13132 18564 13184
rect 18972 13132 19024 13184
rect 21272 13175 21324 13184
rect 21272 13141 21281 13175
rect 21281 13141 21315 13175
rect 21315 13141 21324 13175
rect 21272 13132 21324 13141
rect 22008 13132 22060 13184
rect 22100 13132 22152 13184
rect 25688 13209 25697 13243
rect 25697 13209 25731 13243
rect 25731 13209 25740 13243
rect 25688 13200 25740 13209
rect 26332 13243 26384 13252
rect 26332 13209 26341 13243
rect 26341 13209 26375 13243
rect 26375 13209 26384 13243
rect 26332 13200 26384 13209
rect 27160 13200 27212 13252
rect 28080 13243 28132 13252
rect 28080 13209 28089 13243
rect 28089 13209 28123 13243
rect 28123 13209 28132 13243
rect 28080 13200 28132 13209
rect 28172 13243 28224 13252
rect 28172 13209 28181 13243
rect 28181 13209 28215 13243
rect 28215 13209 28224 13243
rect 28172 13200 28224 13209
rect 29460 13132 29512 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3976 12928 4028 12980
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 2780 12835 2832 12844
rect 2780 12801 2789 12835
rect 2789 12801 2823 12835
rect 2823 12801 2832 12835
rect 5632 12860 5684 12912
rect 6276 12860 6328 12912
rect 6828 12903 6880 12912
rect 6828 12869 6837 12903
rect 6837 12869 6871 12903
rect 6871 12869 6880 12903
rect 6828 12860 6880 12869
rect 7380 12903 7432 12912
rect 7380 12869 7389 12903
rect 7389 12869 7423 12903
rect 7423 12869 7432 12903
rect 7380 12860 7432 12869
rect 7472 12860 7524 12912
rect 9220 12928 9272 12980
rect 9404 12928 9456 12980
rect 9588 12928 9640 12980
rect 2780 12792 2832 12801
rect 3792 12792 3844 12844
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 4988 12792 5040 12844
rect 5540 12792 5592 12844
rect 6552 12792 6604 12844
rect 11704 12928 11756 12980
rect 11888 12928 11940 12980
rect 12440 12928 12492 12980
rect 11060 12860 11112 12912
rect 11244 12792 11296 12844
rect 11520 12792 11572 12844
rect 12072 12860 12124 12912
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 2872 12631 2924 12640
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 2872 12588 2924 12597
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 4712 12588 4764 12640
rect 4896 12588 4948 12640
rect 6092 12656 6144 12708
rect 6460 12656 6512 12708
rect 9220 12724 9272 12776
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 10048 12724 10100 12776
rect 10416 12724 10468 12776
rect 12624 12767 12676 12776
rect 12624 12733 12633 12767
rect 12633 12733 12667 12767
rect 12667 12733 12676 12767
rect 12624 12724 12676 12733
rect 15660 12928 15712 12980
rect 16396 12928 16448 12980
rect 14740 12860 14792 12912
rect 24216 12928 24268 12980
rect 24768 12928 24820 12980
rect 25320 12928 25372 12980
rect 25688 12928 25740 12980
rect 22376 12903 22428 12912
rect 22376 12869 22385 12903
rect 22385 12869 22419 12903
rect 22419 12869 22428 12903
rect 22376 12860 22428 12869
rect 26792 12860 26844 12912
rect 29368 12928 29420 12980
rect 36728 12860 36780 12912
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 20444 12835 20496 12844
rect 16120 12724 16172 12776
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 17960 12767 18012 12776
rect 17960 12733 17969 12767
rect 17969 12733 18003 12767
rect 18003 12733 18012 12767
rect 17960 12724 18012 12733
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 18696 12724 18748 12776
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 20720 12792 20772 12844
rect 21456 12792 21508 12844
rect 23388 12792 23440 12844
rect 20352 12724 20404 12776
rect 22652 12724 22704 12776
rect 24308 12792 24360 12844
rect 11704 12656 11756 12708
rect 10232 12588 10284 12640
rect 11060 12588 11112 12640
rect 11244 12588 11296 12640
rect 12072 12588 12124 12640
rect 13728 12588 13780 12640
rect 22928 12699 22980 12708
rect 22928 12665 22937 12699
rect 22937 12665 22971 12699
rect 22971 12665 22980 12699
rect 22928 12656 22980 12665
rect 36912 12792 36964 12844
rect 27620 12724 27672 12776
rect 28816 12767 28868 12776
rect 28816 12733 28825 12767
rect 28825 12733 28859 12767
rect 28859 12733 28868 12767
rect 28816 12724 28868 12733
rect 29000 12767 29052 12776
rect 29000 12733 29009 12767
rect 29009 12733 29043 12767
rect 29043 12733 29052 12767
rect 29000 12724 29052 12733
rect 19432 12588 19484 12640
rect 20444 12588 20496 12640
rect 20812 12588 20864 12640
rect 21732 12588 21784 12640
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 24308 12588 24360 12640
rect 27528 12588 27580 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1952 12384 2004 12436
rect 6092 12384 6144 12436
rect 6552 12384 6604 12436
rect 7380 12384 7432 12436
rect 8484 12384 8536 12436
rect 8852 12384 8904 12436
rect 10416 12384 10468 12436
rect 11336 12384 11388 12436
rect 2872 12248 2924 12300
rect 4988 12248 5040 12300
rect 8484 12248 8536 12300
rect 9404 12248 9456 12300
rect 9772 12248 9824 12300
rect 9864 12248 9916 12300
rect 10324 12248 10376 12300
rect 11612 12248 11664 12300
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 2136 12180 2188 12232
rect 5908 12180 5960 12232
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 8116 12180 8168 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 11888 12180 11940 12232
rect 6920 12112 6972 12164
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 8484 12087 8536 12096
rect 7840 12044 7892 12053
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 9864 12112 9916 12164
rect 10232 12112 10284 12164
rect 11796 12112 11848 12164
rect 12348 12112 12400 12164
rect 11060 12044 11112 12096
rect 11336 12044 11388 12096
rect 11980 12044 12032 12096
rect 13912 12112 13964 12164
rect 14188 12384 14240 12436
rect 16304 12384 16356 12436
rect 14096 12316 14148 12368
rect 14740 12316 14792 12368
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16672 12248 16724 12300
rect 16396 12112 16448 12164
rect 15200 12044 15252 12096
rect 23756 12384 23808 12436
rect 27344 12384 27396 12436
rect 29000 12384 29052 12436
rect 19432 12316 19484 12368
rect 21088 12316 21140 12368
rect 21272 12316 21324 12368
rect 22008 12316 22060 12368
rect 18604 12112 18656 12164
rect 18328 12044 18380 12096
rect 18880 12044 18932 12096
rect 19248 12044 19300 12096
rect 19708 12112 19760 12164
rect 20812 12112 20864 12164
rect 20536 12044 20588 12096
rect 20720 12044 20772 12096
rect 22376 12248 22428 12300
rect 23020 12248 23072 12300
rect 22928 12223 22980 12232
rect 22928 12189 22937 12223
rect 22937 12189 22971 12223
rect 22971 12189 22980 12223
rect 22928 12180 22980 12189
rect 23204 12180 23256 12232
rect 23296 12180 23348 12232
rect 27620 12291 27672 12300
rect 27620 12257 27629 12291
rect 27629 12257 27663 12291
rect 27663 12257 27672 12291
rect 27620 12248 27672 12257
rect 30840 12291 30892 12300
rect 30840 12257 30849 12291
rect 30849 12257 30883 12291
rect 30883 12257 30892 12291
rect 30840 12248 30892 12257
rect 24952 12180 25004 12232
rect 26884 12180 26936 12232
rect 28264 12223 28316 12232
rect 28264 12189 28273 12223
rect 28273 12189 28307 12223
rect 28307 12189 28316 12223
rect 28264 12180 28316 12189
rect 29828 12155 29880 12164
rect 29828 12121 29837 12155
rect 29837 12121 29871 12155
rect 29871 12121 29880 12155
rect 29828 12112 29880 12121
rect 21272 12087 21324 12096
rect 21272 12053 21281 12087
rect 21281 12053 21315 12087
rect 21315 12053 21324 12087
rect 21272 12044 21324 12053
rect 21640 12044 21692 12096
rect 23020 12044 23072 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 2780 11840 2832 11892
rect 2504 11772 2556 11824
rect 11336 11840 11388 11892
rect 16304 11883 16356 11892
rect 6828 11772 6880 11824
rect 8116 11772 8168 11824
rect 9036 11772 9088 11824
rect 11244 11772 11296 11824
rect 11888 11772 11940 11824
rect 1768 11747 1820 11756
rect 1768 11713 1777 11747
rect 1777 11713 1811 11747
rect 1811 11713 1820 11747
rect 1768 11704 1820 11713
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 1584 11568 1636 11620
rect 5632 11704 5684 11756
rect 7012 11704 7064 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 16304 11849 16313 11883
rect 16313 11849 16347 11883
rect 16347 11849 16356 11883
rect 16304 11840 16356 11849
rect 12348 11772 12400 11824
rect 12624 11772 12676 11824
rect 12808 11772 12860 11824
rect 13820 11772 13872 11824
rect 14280 11772 14332 11824
rect 21272 11840 21324 11892
rect 21456 11840 21508 11892
rect 22100 11840 22152 11892
rect 19524 11772 19576 11824
rect 14372 11704 14424 11756
rect 14556 11747 14608 11756
rect 14556 11713 14565 11747
rect 14565 11713 14599 11747
rect 14599 11713 14608 11747
rect 14556 11704 14608 11713
rect 6000 11636 6052 11688
rect 5632 11568 5684 11620
rect 7196 11636 7248 11688
rect 8300 11636 8352 11688
rect 11060 11636 11112 11688
rect 9220 11568 9272 11620
rect 11704 11636 11756 11688
rect 13084 11636 13136 11688
rect 13820 11636 13872 11688
rect 11888 11568 11940 11620
rect 12072 11568 12124 11620
rect 14188 11636 14240 11688
rect 14556 11568 14608 11620
rect 7656 11500 7708 11552
rect 9036 11500 9088 11552
rect 9496 11500 9548 11552
rect 16672 11704 16724 11756
rect 18052 11704 18104 11756
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 17040 11679 17092 11688
rect 17040 11645 17049 11679
rect 17049 11645 17083 11679
rect 17083 11645 17092 11679
rect 17040 11636 17092 11645
rect 18512 11636 18564 11688
rect 19064 11636 19116 11688
rect 20904 11636 20956 11688
rect 21088 11679 21140 11688
rect 21088 11645 21097 11679
rect 21097 11645 21131 11679
rect 21131 11645 21140 11679
rect 21088 11636 21140 11645
rect 22284 11636 22336 11688
rect 23020 11815 23072 11824
rect 23020 11781 23029 11815
rect 23029 11781 23063 11815
rect 23063 11781 23072 11815
rect 23020 11772 23072 11781
rect 23388 11840 23440 11892
rect 25412 11840 25464 11892
rect 26792 11840 26844 11892
rect 28264 11840 28316 11892
rect 36912 11840 36964 11892
rect 27252 11815 27304 11824
rect 27252 11781 27261 11815
rect 27261 11781 27295 11815
rect 27295 11781 27304 11815
rect 27252 11772 27304 11781
rect 27344 11815 27396 11824
rect 27344 11781 27353 11815
rect 27353 11781 27387 11815
rect 27387 11781 27396 11815
rect 27344 11772 27396 11781
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 25136 11704 25188 11756
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 33232 11704 33284 11756
rect 23112 11636 23164 11688
rect 26148 11636 26200 11688
rect 27436 11636 27488 11688
rect 27620 11636 27672 11688
rect 16120 11500 16172 11552
rect 21272 11500 21324 11552
rect 22376 11500 22428 11552
rect 24676 11568 24728 11620
rect 26332 11568 26384 11620
rect 23480 11500 23532 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3424 11296 3476 11348
rect 5080 11296 5132 11348
rect 6828 11296 6880 11348
rect 6920 11296 6972 11348
rect 7564 11296 7616 11348
rect 8300 11296 8352 11348
rect 9312 11296 9364 11348
rect 12440 11296 12492 11348
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 16856 11339 16908 11348
rect 16856 11305 16886 11339
rect 16886 11305 16908 11339
rect 16856 11296 16908 11305
rect 17500 11296 17552 11348
rect 18328 11339 18380 11348
rect 18328 11305 18337 11339
rect 18337 11305 18371 11339
rect 18371 11305 18380 11339
rect 18328 11296 18380 11305
rect 21272 11296 21324 11348
rect 21364 11296 21416 11348
rect 21548 11296 21600 11348
rect 22008 11296 22060 11348
rect 22100 11296 22152 11348
rect 8760 11228 8812 11280
rect 11888 11228 11940 11280
rect 12992 11228 13044 11280
rect 18052 11228 18104 11280
rect 19248 11228 19300 11280
rect 2688 11160 2740 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 9220 11160 9272 11212
rect 9404 11160 9456 11212
rect 11244 11160 11296 11212
rect 11612 11160 11664 11212
rect 13176 11160 13228 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 15936 11160 15988 11212
rect 4988 11092 5040 11144
rect 6092 11092 6144 11144
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 5540 11024 5592 11076
rect 7012 11024 7064 11076
rect 7196 11024 7248 11076
rect 2780 10956 2832 11008
rect 5264 10956 5316 11008
rect 6460 10956 6512 11008
rect 8668 10956 8720 11008
rect 9036 10956 9088 11008
rect 9496 11092 9548 11144
rect 9588 11092 9640 11144
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 21088 11092 21140 11144
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 24676 11296 24728 11348
rect 25596 11296 25648 11348
rect 27344 11296 27396 11348
rect 33232 11339 33284 11348
rect 33232 11305 33241 11339
rect 33241 11305 33275 11339
rect 33275 11305 33284 11339
rect 33232 11296 33284 11305
rect 25412 11092 25464 11144
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 29276 11092 29328 11144
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 10324 11024 10376 11076
rect 10876 11067 10928 11076
rect 10876 11033 10885 11067
rect 10885 11033 10919 11067
rect 10919 11033 10928 11067
rect 10876 11024 10928 11033
rect 11336 11024 11388 11076
rect 12164 11024 12216 11076
rect 17316 11024 17368 11076
rect 19064 11024 19116 11076
rect 10968 10956 11020 11008
rect 14740 10956 14792 11008
rect 17040 10956 17092 11008
rect 22284 11067 22336 11076
rect 22284 11033 22293 11067
rect 22293 11033 22327 11067
rect 22327 11033 22336 11067
rect 22284 11024 22336 11033
rect 22744 11024 22796 11076
rect 23756 10999 23808 11008
rect 23756 10965 23765 10999
rect 23765 10965 23799 10999
rect 23799 10965 23808 10999
rect 23756 10956 23808 10965
rect 23848 10956 23900 11008
rect 38016 10956 38068 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4620 10752 4672 10804
rect 5816 10752 5868 10804
rect 6552 10752 6604 10804
rect 6736 10752 6788 10804
rect 6920 10752 6972 10804
rect 8024 10752 8076 10804
rect 12808 10752 12860 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 2780 10616 2832 10668
rect 3148 10616 3200 10668
rect 4620 10616 4672 10668
rect 5632 10616 5684 10668
rect 6276 10616 6328 10668
rect 6460 10616 6512 10668
rect 6920 10616 6972 10668
rect 1952 10548 2004 10600
rect 2504 10548 2556 10600
rect 6736 10548 6788 10600
rect 7380 10616 7432 10668
rect 9404 10616 9456 10668
rect 10232 10616 10284 10668
rect 10508 10616 10560 10668
rect 10968 10616 11020 10668
rect 11612 10548 11664 10600
rect 12900 10616 12952 10668
rect 13268 10752 13320 10804
rect 13820 10752 13872 10804
rect 17776 10752 17828 10804
rect 19340 10752 19392 10804
rect 13452 10684 13504 10736
rect 14280 10684 14332 10736
rect 16488 10684 16540 10736
rect 19156 10684 19208 10736
rect 21272 10752 21324 10804
rect 22652 10752 22704 10804
rect 26700 10752 26752 10804
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 14004 10548 14056 10600
rect 9128 10480 9180 10532
rect 12624 10480 12676 10532
rect 2044 10412 2096 10464
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 6920 10412 6972 10464
rect 7196 10412 7248 10464
rect 7564 10412 7616 10464
rect 8208 10412 8260 10464
rect 8300 10412 8352 10464
rect 9404 10412 9456 10464
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 10876 10455 10928 10464
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 11612 10412 11664 10464
rect 12716 10412 12768 10464
rect 21456 10684 21508 10736
rect 21916 10684 21968 10736
rect 22008 10659 22060 10668
rect 15660 10548 15712 10600
rect 17132 10548 17184 10600
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 37832 10616 37884 10668
rect 19248 10591 19300 10600
rect 19248 10557 19257 10591
rect 19257 10557 19291 10591
rect 19291 10557 19300 10591
rect 19248 10548 19300 10557
rect 20076 10548 20128 10600
rect 21180 10548 21232 10600
rect 21824 10480 21876 10532
rect 22928 10548 22980 10600
rect 23572 10548 23624 10600
rect 28080 10548 28132 10600
rect 28540 10548 28592 10600
rect 23388 10480 23440 10532
rect 28448 10523 28500 10532
rect 16488 10412 16540 10464
rect 17132 10412 17184 10464
rect 17592 10412 17644 10464
rect 28448 10489 28457 10523
rect 28457 10489 28491 10523
rect 28491 10489 28500 10523
rect 28448 10480 28500 10489
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 10048 10208 10100 10260
rect 8300 10072 8352 10124
rect 1952 10004 2004 10056
rect 2688 10047 2740 10056
rect 2688 10013 2697 10047
rect 2697 10013 2731 10047
rect 2731 10013 2740 10047
rect 2688 10004 2740 10013
rect 2964 10004 3016 10056
rect 3792 10004 3844 10056
rect 4068 10004 4120 10056
rect 4896 10004 4948 10056
rect 6276 10004 6328 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 3792 9868 3844 9920
rect 4988 9868 5040 9920
rect 5264 9868 5316 9920
rect 7196 9936 7248 9988
rect 7380 9936 7432 9988
rect 7564 9936 7616 9988
rect 23756 10208 23808 10260
rect 37832 10251 37884 10260
rect 37832 10217 37841 10251
rect 37841 10217 37875 10251
rect 37875 10217 37884 10251
rect 37832 10208 37884 10217
rect 11244 10140 11296 10192
rect 13268 10140 13320 10192
rect 15200 10140 15252 10192
rect 15660 10072 15712 10124
rect 18144 10140 18196 10192
rect 19432 10140 19484 10192
rect 21272 10140 21324 10192
rect 23204 10140 23256 10192
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 13728 10004 13780 10056
rect 9956 9936 10008 9988
rect 7932 9868 7984 9920
rect 8116 9868 8168 9920
rect 12624 9936 12676 9988
rect 14740 9936 14792 9988
rect 15108 9936 15160 9988
rect 18696 10004 18748 10056
rect 19432 10004 19484 10056
rect 23112 10072 23164 10124
rect 28448 10140 28500 10192
rect 23388 10072 23440 10124
rect 22008 10004 22060 10056
rect 16672 9936 16724 9988
rect 21916 9936 21968 9988
rect 23756 9936 23808 9988
rect 24400 10004 24452 10056
rect 25228 10047 25280 10056
rect 25228 10013 25237 10047
rect 25237 10013 25271 10047
rect 25271 10013 25280 10047
rect 25228 10004 25280 10013
rect 38016 10047 38068 10056
rect 38016 10013 38025 10047
rect 38025 10013 38059 10047
rect 38059 10013 38068 10047
rect 38016 10004 38068 10013
rect 12532 9868 12584 9920
rect 13544 9868 13596 9920
rect 15292 9868 15344 9920
rect 15384 9868 15436 9920
rect 21180 9868 21232 9920
rect 23664 9868 23716 9920
rect 24860 9868 24912 9920
rect 27436 9911 27488 9920
rect 27436 9877 27445 9911
rect 27445 9877 27479 9911
rect 27479 9877 27488 9911
rect 27436 9868 27488 9877
rect 29184 9936 29236 9988
rect 29828 9979 29880 9988
rect 29828 9945 29837 9979
rect 29837 9945 29871 9979
rect 29871 9945 29880 9979
rect 29828 9936 29880 9945
rect 29920 9979 29972 9988
rect 29920 9945 29929 9979
rect 29929 9945 29963 9979
rect 29963 9945 29972 9979
rect 29920 9936 29972 9945
rect 30012 9868 30064 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2688 9664 2740 9716
rect 1952 9596 2004 9648
rect 2780 9528 2832 9580
rect 1860 9460 1912 9512
rect 3056 9596 3108 9648
rect 4988 9596 5040 9648
rect 6276 9664 6328 9716
rect 9220 9664 9272 9716
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3332 9460 3384 9512
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 4988 9460 5040 9512
rect 6828 9528 6880 9580
rect 8668 9460 8720 9512
rect 9680 9664 9732 9716
rect 11336 9664 11388 9716
rect 12348 9664 12400 9716
rect 10232 9596 10284 9648
rect 17500 9664 17552 9716
rect 20168 9664 20220 9716
rect 20628 9664 20680 9716
rect 22652 9664 22704 9716
rect 25228 9664 25280 9716
rect 29920 9707 29972 9716
rect 29920 9673 29929 9707
rect 29929 9673 29963 9707
rect 29963 9673 29972 9707
rect 29920 9664 29972 9673
rect 30012 9664 30064 9716
rect 34520 9664 34572 9716
rect 13912 9596 13964 9648
rect 11060 9528 11112 9580
rect 12992 9528 13044 9580
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 6920 9392 6972 9444
rect 8852 9392 8904 9444
rect 9772 9460 9824 9512
rect 15844 9596 15896 9648
rect 19984 9596 20036 9648
rect 24768 9639 24820 9648
rect 24768 9605 24777 9639
rect 24777 9605 24811 9639
rect 24811 9605 24820 9639
rect 24768 9596 24820 9605
rect 24860 9639 24912 9648
rect 24860 9605 24869 9639
rect 24869 9605 24903 9639
rect 24903 9605 24912 9639
rect 27436 9639 27488 9648
rect 24860 9596 24912 9605
rect 27436 9605 27445 9639
rect 27445 9605 27479 9639
rect 27479 9605 27488 9639
rect 27436 9596 27488 9605
rect 28356 9596 28408 9648
rect 28816 9596 28868 9648
rect 15016 9528 15068 9580
rect 16304 9528 16356 9580
rect 16672 9460 16724 9512
rect 17132 9503 17184 9512
rect 16120 9392 16172 9444
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 17500 9460 17552 9512
rect 8024 9324 8076 9376
rect 9312 9324 9364 9376
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 11336 9324 11388 9376
rect 17224 9324 17276 9376
rect 17592 9324 17644 9376
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 18696 9324 18748 9376
rect 18972 9324 19024 9376
rect 19432 9460 19484 9512
rect 19156 9392 19208 9444
rect 21640 9460 21692 9512
rect 23388 9528 23440 9580
rect 24216 9528 24268 9580
rect 25412 9528 25464 9580
rect 25872 9571 25924 9580
rect 25872 9537 25881 9571
rect 25881 9537 25915 9571
rect 25915 9537 25924 9571
rect 25872 9528 25924 9537
rect 29644 9528 29696 9580
rect 32404 9528 32456 9580
rect 24768 9460 24820 9512
rect 27988 9503 28040 9512
rect 27988 9469 27997 9503
rect 27997 9469 28031 9503
rect 28031 9469 28040 9503
rect 27988 9460 28040 9469
rect 20904 9392 20956 9444
rect 21364 9324 21416 9376
rect 22560 9367 22612 9376
rect 22560 9333 22569 9367
rect 22569 9333 22603 9367
rect 22603 9333 22612 9367
rect 22560 9324 22612 9333
rect 23112 9324 23164 9376
rect 24952 9392 25004 9444
rect 29276 9392 29328 9444
rect 24492 9324 24544 9376
rect 29920 9324 29972 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4620 9120 4672 9172
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 3240 9052 3292 9104
rect 9404 9120 9456 9172
rect 8024 9052 8076 9104
rect 11152 9120 11204 9172
rect 14188 9120 14240 9172
rect 14280 9120 14332 9172
rect 13452 9052 13504 9104
rect 15476 9120 15528 9172
rect 15568 9120 15620 9172
rect 16580 9120 16632 9172
rect 16856 9163 16908 9172
rect 16856 9129 16865 9163
rect 16865 9129 16899 9163
rect 16899 9129 16908 9163
rect 16856 9120 16908 9129
rect 17868 9120 17920 9172
rect 18420 9052 18472 9104
rect 18972 9052 19024 9104
rect 3148 8984 3200 9036
rect 8392 8984 8444 9036
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3884 8916 3936 8968
rect 4712 8916 4764 8968
rect 6460 8916 6512 8968
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 8576 8916 8628 8968
rect 10416 8984 10468 9036
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 12900 8984 12952 9036
rect 16120 8984 16172 9036
rect 16396 8984 16448 9036
rect 19708 9052 19760 9104
rect 21180 9120 21232 9172
rect 24676 9120 24728 9172
rect 24768 9120 24820 9172
rect 32128 9120 32180 9172
rect 19340 8984 19392 9036
rect 21824 8984 21876 9036
rect 22008 8984 22060 9036
rect 23756 9052 23808 9104
rect 25780 9052 25832 9104
rect 25872 9052 25924 9104
rect 26148 9052 26200 9104
rect 26424 8984 26476 9036
rect 27988 9052 28040 9104
rect 33048 9052 33100 9104
rect 2044 8780 2096 8832
rect 3056 8780 3108 8832
rect 4988 8780 5040 8832
rect 8760 8848 8812 8900
rect 16672 8916 16724 8968
rect 18420 8959 18472 8968
rect 7748 8780 7800 8832
rect 8024 8780 8076 8832
rect 9680 8780 9732 8832
rect 10048 8848 10100 8900
rect 12164 8891 12216 8900
rect 12164 8857 12173 8891
rect 12173 8857 12207 8891
rect 12207 8857 12216 8891
rect 12164 8848 12216 8857
rect 12256 8848 12308 8900
rect 15476 8848 15528 8900
rect 17684 8848 17736 8900
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 21456 8916 21508 8968
rect 20168 8848 20220 8900
rect 21824 8891 21876 8900
rect 13728 8780 13780 8832
rect 21088 8780 21140 8832
rect 21824 8857 21833 8891
rect 21833 8857 21867 8891
rect 21867 8857 21876 8891
rect 21824 8848 21876 8857
rect 24492 8916 24544 8968
rect 24676 8916 24728 8968
rect 25412 8916 25464 8968
rect 34520 8916 34572 8968
rect 36084 8916 36136 8968
rect 22468 8848 22520 8900
rect 26148 8891 26200 8900
rect 26148 8857 26157 8891
rect 26157 8857 26191 8891
rect 26191 8857 26200 8891
rect 26148 8848 26200 8857
rect 26240 8891 26292 8900
rect 26240 8857 26249 8891
rect 26249 8857 26283 8891
rect 26283 8857 26292 8891
rect 26240 8848 26292 8857
rect 25228 8780 25280 8832
rect 36268 8780 36320 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3608 8576 3660 8628
rect 6000 8619 6052 8628
rect 3148 8508 3200 8560
rect 2688 8440 2740 8492
rect 4620 8508 4672 8560
rect 6000 8585 6009 8619
rect 6009 8585 6043 8619
rect 6043 8585 6052 8619
rect 6000 8576 6052 8585
rect 9680 8576 9732 8628
rect 10508 8576 10560 8628
rect 14372 8576 14424 8628
rect 15016 8576 15068 8628
rect 16672 8576 16724 8628
rect 11612 8508 11664 8560
rect 11888 8508 11940 8560
rect 13452 8551 13504 8560
rect 13452 8517 13461 8551
rect 13461 8517 13495 8551
rect 13495 8517 13504 8551
rect 13452 8508 13504 8517
rect 13544 8508 13596 8560
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 10232 8440 10284 8492
rect 12348 8440 12400 8492
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 16120 8440 16172 8492
rect 19432 8576 19484 8628
rect 19524 8576 19576 8628
rect 23204 8576 23256 8628
rect 28356 8619 28408 8628
rect 28356 8585 28365 8619
rect 28365 8585 28399 8619
rect 28399 8585 28408 8619
rect 28356 8576 28408 8585
rect 28540 8576 28592 8628
rect 36084 8619 36136 8628
rect 36084 8585 36093 8619
rect 36093 8585 36127 8619
rect 36127 8585 36136 8619
rect 36084 8576 36136 8585
rect 21640 8508 21692 8560
rect 23664 8551 23716 8560
rect 23664 8517 23673 8551
rect 23673 8517 23707 8551
rect 23707 8517 23716 8551
rect 23664 8508 23716 8517
rect 25228 8551 25280 8560
rect 25228 8517 25237 8551
rect 25237 8517 25271 8551
rect 25271 8517 25280 8551
rect 25228 8508 25280 8517
rect 25320 8508 25372 8560
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 2320 8304 2372 8356
rect 6828 8372 6880 8424
rect 13544 8372 13596 8424
rect 16948 8372 17000 8424
rect 17592 8372 17644 8424
rect 8576 8304 8628 8356
rect 12164 8304 12216 8356
rect 4620 8236 4672 8288
rect 8760 8236 8812 8288
rect 9128 8236 9180 8288
rect 11244 8236 11296 8288
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 18604 8304 18656 8356
rect 21088 8372 21140 8424
rect 23112 8440 23164 8492
rect 26056 8440 26108 8492
rect 28356 8440 28408 8492
rect 29092 8440 29144 8492
rect 35808 8440 35860 8492
rect 36268 8483 36320 8492
rect 36268 8449 36277 8483
rect 36277 8449 36311 8483
rect 36311 8449 36320 8483
rect 36268 8440 36320 8449
rect 21364 8372 21416 8424
rect 23020 8372 23072 8424
rect 24032 8415 24084 8424
rect 24032 8381 24041 8415
rect 24041 8381 24075 8415
rect 24075 8381 24084 8415
rect 24032 8372 24084 8381
rect 24860 8372 24912 8424
rect 25964 8372 26016 8424
rect 26608 8372 26660 8424
rect 18972 8279 19024 8288
rect 18972 8245 18981 8279
rect 18981 8245 19015 8279
rect 19015 8245 19024 8279
rect 18972 8236 19024 8245
rect 23480 8304 23532 8356
rect 28448 8304 28500 8356
rect 28356 8236 28408 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2412 8032 2464 8084
rect 3976 8032 4028 8084
rect 6000 8032 6052 8084
rect 6368 8075 6420 8084
rect 6368 8041 6377 8075
rect 6377 8041 6411 8075
rect 6411 8041 6420 8075
rect 6368 8032 6420 8041
rect 6092 7964 6144 8016
rect 10140 8032 10192 8084
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 5632 7896 5684 7948
rect 6736 7896 6788 7948
rect 15108 8032 15160 8084
rect 12808 7964 12860 8016
rect 17132 8032 17184 8084
rect 17684 8032 17736 8084
rect 18144 7964 18196 8016
rect 18696 7964 18748 8016
rect 21180 8032 21232 8084
rect 24400 8032 24452 8084
rect 26332 8032 26384 8084
rect 27620 8032 27672 8084
rect 13176 7896 13228 7948
rect 16120 7896 16172 7948
rect 18972 7896 19024 7948
rect 19524 7939 19576 7948
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 20812 7896 20864 7948
rect 24768 7964 24820 8016
rect 22744 7896 22796 7948
rect 24216 7896 24268 7948
rect 25780 7896 25832 7948
rect 26148 7896 26200 7948
rect 28540 7939 28592 7948
rect 28540 7905 28549 7939
rect 28549 7905 28583 7939
rect 28583 7905 28592 7939
rect 28540 7896 28592 7905
rect 29276 7896 29328 7948
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2780 7828 2832 7880
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 12900 7828 12952 7880
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 5908 7760 5960 7812
rect 6184 7760 6236 7812
rect 11244 7803 11296 7812
rect 11244 7769 11253 7803
rect 11253 7769 11287 7803
rect 11287 7769 11296 7803
rect 11244 7760 11296 7769
rect 11888 7760 11940 7812
rect 12532 7760 12584 7812
rect 14740 7803 14792 7812
rect 14740 7769 14749 7803
rect 14749 7769 14783 7803
rect 14783 7769 14792 7803
rect 14740 7760 14792 7769
rect 15108 7760 15160 7812
rect 18788 7760 18840 7812
rect 22836 7828 22888 7880
rect 19892 7760 19944 7812
rect 21088 7760 21140 7812
rect 24216 7760 24268 7812
rect 24952 7760 25004 7812
rect 26148 7760 26200 7812
rect 1676 7692 1728 7744
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 3884 7692 3936 7744
rect 7012 7692 7064 7744
rect 9312 7692 9364 7744
rect 12072 7692 12124 7744
rect 18052 7692 18104 7744
rect 18972 7692 19024 7744
rect 21180 7692 21232 7744
rect 22744 7692 22796 7744
rect 26332 7692 26384 7744
rect 27620 7760 27672 7812
rect 27896 7692 27948 7744
rect 31576 7692 31628 7744
rect 38200 7735 38252 7744
rect 38200 7701 38209 7735
rect 38209 7701 38243 7735
rect 38243 7701 38252 7735
rect 38200 7692 38252 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 5356 7488 5408 7540
rect 5632 7420 5684 7472
rect 6644 7463 6696 7472
rect 6644 7429 6653 7463
rect 6653 7429 6687 7463
rect 6687 7429 6696 7463
rect 6644 7420 6696 7429
rect 6920 7420 6972 7472
rect 8300 7420 8352 7472
rect 9772 7488 9824 7540
rect 10508 7488 10560 7540
rect 10232 7463 10284 7472
rect 10232 7429 10241 7463
rect 10241 7429 10275 7463
rect 10275 7429 10284 7463
rect 10232 7420 10284 7429
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 1952 7352 2004 7404
rect 3792 7395 3844 7404
rect 3792 7361 3801 7395
rect 3801 7361 3835 7395
rect 3835 7361 3844 7395
rect 3792 7352 3844 7361
rect 3884 7352 3936 7404
rect 5540 7352 5592 7404
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 2228 7284 2280 7336
rect 6184 7284 6236 7336
rect 7012 7284 7064 7336
rect 10140 7352 10192 7404
rect 15016 7488 15068 7540
rect 10876 7420 10928 7472
rect 11888 7420 11940 7472
rect 13268 7463 13320 7472
rect 13268 7429 13277 7463
rect 13277 7429 13311 7463
rect 13311 7429 13320 7463
rect 13268 7420 13320 7429
rect 20444 7488 20496 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 21272 7488 21324 7540
rect 19800 7420 19852 7472
rect 20996 7420 21048 7472
rect 24032 7420 24084 7472
rect 24216 7463 24268 7472
rect 24216 7429 24225 7463
rect 24225 7429 24259 7463
rect 24259 7429 24268 7463
rect 24216 7420 24268 7429
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 26240 7488 26292 7540
rect 11152 7352 11204 7404
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 23756 7352 23808 7404
rect 26792 7420 26844 7472
rect 27160 7395 27212 7404
rect 9772 7327 9824 7336
rect 2136 7216 2188 7268
rect 9772 7293 9781 7327
rect 9781 7293 9815 7327
rect 9815 7293 9824 7327
rect 9772 7284 9824 7293
rect 10048 7284 10100 7336
rect 16856 7327 16908 7336
rect 9864 7216 9916 7268
rect 6092 7148 6144 7200
rect 7104 7148 7156 7200
rect 11428 7148 11480 7200
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 18604 7284 18656 7336
rect 19340 7284 19392 7336
rect 19800 7284 19852 7336
rect 22008 7284 22060 7336
rect 23480 7284 23532 7336
rect 24032 7284 24084 7336
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 26240 7284 26292 7336
rect 27252 7284 27304 7336
rect 31668 7284 31720 7336
rect 15108 7148 15160 7200
rect 16764 7148 16816 7200
rect 18788 7148 18840 7200
rect 20720 7148 20772 7200
rect 20904 7148 20956 7200
rect 21916 7216 21968 7268
rect 23940 7216 23992 7268
rect 24124 7216 24176 7268
rect 25044 7216 25096 7268
rect 26148 7216 26200 7268
rect 22100 7148 22152 7200
rect 34520 7148 34572 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 9312 6944 9364 6996
rect 18696 6944 18748 6996
rect 20352 6944 20404 6996
rect 20444 6944 20496 6996
rect 27252 6944 27304 6996
rect 3976 6808 4028 6860
rect 4252 6808 4304 6860
rect 2228 6740 2280 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3240 6672 3292 6724
rect 4620 6672 4672 6724
rect 5356 6672 5408 6724
rect 6736 6808 6788 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 8116 6808 8168 6860
rect 9680 6808 9732 6860
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12072 6808 12124 6860
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 12256 6740 12308 6792
rect 14740 6808 14792 6860
rect 15108 6783 15160 6792
rect 7012 6672 7064 6724
rect 7656 6672 7708 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 2504 6604 2556 6656
rect 4712 6604 4764 6656
rect 5632 6604 5684 6656
rect 7288 6604 7340 6656
rect 7380 6604 7432 6656
rect 9588 6672 9640 6724
rect 9956 6672 10008 6724
rect 12440 6672 12492 6724
rect 14740 6672 14792 6724
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 11428 6604 11480 6656
rect 12348 6604 12400 6656
rect 13728 6604 13780 6656
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 16672 6672 16724 6724
rect 21088 6876 21140 6928
rect 19432 6808 19484 6860
rect 21180 6808 21232 6860
rect 23480 6876 23532 6928
rect 25320 6876 25372 6928
rect 27804 6851 27856 6860
rect 26148 6740 26200 6792
rect 27804 6817 27813 6851
rect 27813 6817 27847 6851
rect 27847 6817 27856 6851
rect 27804 6808 27856 6817
rect 28448 6783 28500 6792
rect 28448 6749 28457 6783
rect 28457 6749 28491 6783
rect 28491 6749 28500 6783
rect 28448 6740 28500 6749
rect 29092 6740 29144 6792
rect 19892 6672 19944 6724
rect 22192 6715 22244 6724
rect 17684 6604 17736 6656
rect 17960 6604 18012 6656
rect 20904 6604 20956 6656
rect 21456 6647 21508 6656
rect 21456 6613 21465 6647
rect 21465 6613 21499 6647
rect 21499 6613 21508 6647
rect 21456 6604 21508 6613
rect 22192 6681 22201 6715
rect 22201 6681 22235 6715
rect 22235 6681 22244 6715
rect 22192 6672 22244 6681
rect 24676 6672 24728 6724
rect 24768 6672 24820 6724
rect 22100 6604 22152 6656
rect 22284 6604 22336 6656
rect 25964 6672 26016 6724
rect 26608 6647 26660 6656
rect 26608 6613 26617 6647
rect 26617 6613 26651 6647
rect 26651 6613 26660 6647
rect 26608 6604 26660 6613
rect 27804 6604 27856 6656
rect 34336 6808 34388 6860
rect 34520 6740 34572 6792
rect 30656 6604 30708 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 3424 6400 3476 6452
rect 5356 6400 5408 6452
rect 6920 6400 6972 6452
rect 9036 6400 9088 6452
rect 4528 6375 4580 6384
rect 4528 6341 4537 6375
rect 4537 6341 4571 6375
rect 4571 6341 4580 6375
rect 4528 6332 4580 6341
rect 5172 6332 5224 6384
rect 1676 6264 1728 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 3608 6264 3660 6316
rect 3976 6264 4028 6316
rect 4252 6307 4304 6316
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 7012 6332 7064 6384
rect 12256 6400 12308 6452
rect 12440 6400 12492 6452
rect 15936 6400 15988 6452
rect 8208 6264 8260 6316
rect 9128 6264 9180 6316
rect 14096 6332 14148 6384
rect 16856 6400 16908 6452
rect 19340 6400 19392 6452
rect 20076 6400 20128 6452
rect 21548 6400 21600 6452
rect 10784 6264 10836 6316
rect 12256 6307 12308 6316
rect 12256 6273 12265 6307
rect 12265 6273 12299 6307
rect 12299 6273 12308 6307
rect 12256 6264 12308 6273
rect 13636 6264 13688 6316
rect 15292 6264 15344 6316
rect 15844 6264 15896 6316
rect 16120 6264 16172 6316
rect 17224 6332 17276 6384
rect 26608 6400 26660 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 27896 6443 27948 6452
rect 27896 6409 27905 6443
rect 27905 6409 27939 6443
rect 27939 6409 27948 6443
rect 27896 6400 27948 6409
rect 29184 6443 29236 6452
rect 29184 6409 29193 6443
rect 29193 6409 29227 6443
rect 29227 6409 29236 6443
rect 29184 6400 29236 6409
rect 29828 6443 29880 6452
rect 29828 6409 29837 6443
rect 29837 6409 29871 6443
rect 29871 6409 29880 6443
rect 29828 6400 29880 6409
rect 23020 6375 23072 6384
rect 23020 6341 23029 6375
rect 23029 6341 23063 6375
rect 23063 6341 23072 6375
rect 23020 6332 23072 6341
rect 28908 6332 28960 6384
rect 30380 6332 30432 6384
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 18236 6264 18288 6316
rect 20996 6264 21048 6316
rect 22468 6264 22520 6316
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 24860 6264 24912 6316
rect 25044 6264 25096 6316
rect 2228 6196 2280 6248
rect 6552 6196 6604 6248
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 2780 6128 2832 6180
rect 8300 6128 8352 6180
rect 2872 6060 2924 6112
rect 5172 6060 5224 6112
rect 6644 6060 6696 6112
rect 8208 6060 8260 6112
rect 10692 6196 10744 6248
rect 16764 6196 16816 6248
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 17224 6196 17276 6248
rect 19248 6196 19300 6248
rect 19340 6196 19392 6248
rect 23572 6196 23624 6248
rect 25872 6307 25924 6316
rect 25872 6273 25881 6307
rect 25881 6273 25915 6307
rect 25915 6273 25924 6307
rect 26424 6307 26476 6316
rect 25872 6264 25924 6273
rect 26424 6273 26433 6307
rect 26433 6273 26467 6307
rect 26467 6273 26476 6307
rect 26424 6264 26476 6273
rect 26148 6196 26200 6248
rect 12164 6128 12216 6180
rect 18328 6128 18380 6180
rect 20720 6128 20772 6180
rect 21180 6128 21232 6180
rect 22100 6128 22152 6180
rect 22192 6128 22244 6180
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 14648 6060 14700 6112
rect 16672 6060 16724 6112
rect 22008 6060 22060 6112
rect 23020 6128 23072 6180
rect 24860 6128 24912 6180
rect 25780 6128 25832 6180
rect 26424 6128 26476 6180
rect 27252 6264 27304 6316
rect 26700 6196 26752 6248
rect 29460 6264 29512 6316
rect 29092 6128 29144 6180
rect 36728 6128 36780 6180
rect 24768 6060 24820 6112
rect 26516 6103 26568 6112
rect 26516 6069 26525 6103
rect 26525 6069 26559 6103
rect 26559 6069 26568 6103
rect 26516 6060 26568 6069
rect 32496 6060 32548 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3148 5856 3200 5908
rect 6276 5856 6328 5908
rect 3884 5720 3936 5772
rect 8576 5856 8628 5908
rect 8852 5856 8904 5908
rect 8208 5788 8260 5840
rect 10784 5856 10836 5908
rect 7012 5720 7064 5772
rect 7288 5720 7340 5772
rect 2504 5652 2556 5704
rect 3976 5695 4028 5704
rect 20 5516 72 5568
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 5724 5652 5776 5704
rect 6000 5652 6052 5704
rect 8392 5720 8444 5772
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 11060 5788 11112 5840
rect 10416 5720 10468 5772
rect 10968 5720 11020 5772
rect 4252 5584 4304 5636
rect 4804 5584 4856 5636
rect 6644 5584 6696 5636
rect 6736 5516 6788 5568
rect 8484 5584 8536 5636
rect 12808 5652 12860 5704
rect 9496 5584 9548 5636
rect 11980 5584 12032 5636
rect 7840 5516 7892 5568
rect 11796 5516 11848 5568
rect 13636 5856 13688 5908
rect 22744 5856 22796 5908
rect 24676 5856 24728 5908
rect 29000 5856 29052 5908
rect 13544 5788 13596 5840
rect 16764 5788 16816 5840
rect 15844 5720 15896 5772
rect 15936 5720 15988 5772
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 16488 5652 16540 5704
rect 17040 5720 17092 5772
rect 21088 5788 21140 5840
rect 19340 5720 19392 5772
rect 20720 5720 20772 5772
rect 32312 5788 32364 5840
rect 24308 5720 24360 5772
rect 24860 5720 24912 5772
rect 24952 5720 25004 5772
rect 26332 5720 26384 5772
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 15292 5584 15344 5636
rect 15384 5627 15436 5636
rect 15384 5593 15393 5627
rect 15393 5593 15427 5627
rect 15427 5593 15436 5627
rect 22008 5695 22060 5704
rect 22008 5661 22017 5695
rect 22017 5661 22051 5695
rect 22051 5661 22060 5695
rect 22008 5652 22060 5661
rect 15384 5584 15436 5593
rect 14372 5516 14424 5568
rect 23848 5652 23900 5704
rect 25412 5652 25464 5704
rect 25688 5652 25740 5704
rect 27528 5720 27580 5772
rect 26792 5652 26844 5704
rect 28264 5720 28316 5772
rect 29276 5720 29328 5772
rect 27804 5695 27856 5704
rect 27804 5661 27813 5695
rect 27813 5661 27847 5695
rect 27847 5661 27856 5695
rect 27804 5652 27856 5661
rect 27988 5652 28040 5704
rect 28908 5652 28960 5704
rect 29092 5652 29144 5704
rect 29644 5652 29696 5704
rect 29920 5695 29972 5704
rect 29920 5661 29929 5695
rect 29929 5661 29963 5695
rect 29963 5661 29972 5695
rect 29920 5652 29972 5661
rect 30380 5695 30432 5704
rect 30380 5661 30389 5695
rect 30389 5661 30423 5695
rect 30423 5661 30432 5695
rect 30380 5652 30432 5661
rect 31024 5695 31076 5704
rect 31024 5661 31033 5695
rect 31033 5661 31067 5695
rect 31067 5661 31076 5695
rect 31024 5652 31076 5661
rect 31852 5695 31904 5704
rect 31852 5661 31861 5695
rect 31861 5661 31895 5695
rect 31895 5661 31904 5695
rect 31852 5652 31904 5661
rect 38016 5695 38068 5704
rect 21088 5516 21140 5568
rect 21548 5559 21600 5568
rect 21548 5525 21557 5559
rect 21557 5525 21591 5559
rect 21591 5525 21600 5559
rect 21548 5516 21600 5525
rect 22008 5516 22060 5568
rect 23664 5516 23716 5568
rect 24768 5627 24820 5636
rect 24768 5593 24777 5627
rect 24777 5593 24811 5627
rect 24811 5593 24820 5627
rect 24768 5584 24820 5593
rect 27344 5584 27396 5636
rect 28540 5584 28592 5636
rect 38016 5661 38025 5695
rect 38025 5661 38059 5695
rect 38059 5661 38068 5695
rect 38016 5652 38068 5661
rect 30564 5516 30616 5568
rect 34612 5516 34664 5568
rect 38016 5516 38068 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 2596 5176 2648 5228
rect 7012 5244 7064 5296
rect 4252 5219 4304 5228
rect 664 4972 716 5024
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 4068 5108 4120 5160
rect 5632 5040 5684 5092
rect 5540 4972 5592 5024
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 6092 5040 6144 5092
rect 11152 5312 11204 5364
rect 8668 5244 8720 5296
rect 10324 5244 10376 5296
rect 14648 5312 14700 5364
rect 13176 5244 13228 5296
rect 22652 5312 22704 5364
rect 23204 5312 23256 5364
rect 26608 5312 26660 5364
rect 15752 5244 15804 5296
rect 19064 5244 19116 5296
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 11520 5176 11572 5228
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 19340 5244 19392 5296
rect 19432 5287 19484 5296
rect 19432 5253 19441 5287
rect 19441 5253 19475 5287
rect 19475 5253 19484 5287
rect 19432 5244 19484 5253
rect 22284 5244 22336 5296
rect 25044 5244 25096 5296
rect 31576 5355 31628 5364
rect 31576 5321 31585 5355
rect 31585 5321 31619 5355
rect 31619 5321 31628 5355
rect 31576 5312 31628 5321
rect 28264 5244 28316 5296
rect 28540 5287 28592 5296
rect 28540 5253 28549 5287
rect 28549 5253 28583 5287
rect 28583 5253 28592 5287
rect 28540 5244 28592 5253
rect 28816 5244 28868 5296
rect 30472 5244 30524 5296
rect 32588 5244 32640 5296
rect 12624 5108 12676 5160
rect 6552 4972 6604 5024
rect 13268 4972 13320 5024
rect 13636 4972 13688 5024
rect 14372 5108 14424 5160
rect 15108 5108 15160 5160
rect 17868 5108 17920 5160
rect 21272 5176 21324 5228
rect 22008 5219 22060 5228
rect 22008 5185 22017 5219
rect 22017 5185 22051 5219
rect 22051 5185 22060 5219
rect 22008 5176 22060 5185
rect 24492 5176 24544 5228
rect 25504 5176 25556 5228
rect 26424 5176 26476 5228
rect 29552 5219 29604 5228
rect 29552 5185 29561 5219
rect 29561 5185 29595 5219
rect 29595 5185 29604 5219
rect 29552 5176 29604 5185
rect 29644 5176 29696 5228
rect 31208 5176 31260 5228
rect 14004 5083 14056 5092
rect 14004 5049 14013 5083
rect 14013 5049 14047 5083
rect 14047 5049 14056 5083
rect 14004 5040 14056 5049
rect 16304 4972 16356 5024
rect 21088 5108 21140 5160
rect 21180 5108 21232 5160
rect 26148 5108 26200 5160
rect 28448 5151 28500 5160
rect 28448 5117 28457 5151
rect 28457 5117 28491 5151
rect 28491 5117 28500 5151
rect 28448 5108 28500 5117
rect 31668 5176 31720 5228
rect 18788 5040 18840 5092
rect 23480 5040 23532 5092
rect 18604 4972 18656 5024
rect 23572 4972 23624 5024
rect 23756 5015 23808 5024
rect 23756 4981 23765 5015
rect 23765 4981 23799 5015
rect 23799 4981 23808 5015
rect 23756 4972 23808 4981
rect 24032 4972 24084 5024
rect 29000 5083 29052 5092
rect 29000 5049 29009 5083
rect 29009 5049 29043 5083
rect 29043 5049 29052 5083
rect 29000 5040 29052 5049
rect 31024 5040 31076 5092
rect 25320 5015 25372 5024
rect 25320 4981 25329 5015
rect 25329 4981 25363 5015
rect 25363 4981 25372 5015
rect 25320 4972 25372 4981
rect 28816 4972 28868 5024
rect 29828 4972 29880 5024
rect 29920 4972 29972 5024
rect 33784 4972 33836 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4252 4768 4304 4820
rect 7932 4811 7984 4820
rect 3608 4700 3660 4752
rect 3884 4700 3936 4752
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8300 4768 8352 4820
rect 11704 4768 11756 4820
rect 21180 4811 21232 4820
rect 9496 4700 9548 4752
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 3516 4496 3568 4548
rect 7012 4632 7064 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 10048 4632 10100 4684
rect 11704 4632 11756 4684
rect 12256 4632 12308 4684
rect 8392 4564 8444 4616
rect 9220 4564 9272 4616
rect 13820 4700 13872 4752
rect 21180 4777 21189 4811
rect 21189 4777 21223 4811
rect 21223 4777 21232 4811
rect 21180 4768 21232 4777
rect 31852 4768 31904 4820
rect 23572 4700 23624 4752
rect 27528 4700 27580 4752
rect 33600 4743 33652 4752
rect 33600 4709 33609 4743
rect 33609 4709 33643 4743
rect 33643 4709 33652 4743
rect 33600 4700 33652 4709
rect 16304 4632 16356 4684
rect 16580 4632 16632 4684
rect 17316 4632 17368 4684
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14556 4564 14608 4616
rect 18604 4632 18656 4684
rect 19156 4632 19208 4684
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 19340 4564 19392 4616
rect 21548 4564 21600 4616
rect 25412 4564 25464 4616
rect 25688 4564 25740 4616
rect 26148 4564 26200 4616
rect 26884 4564 26936 4616
rect 27804 4564 27856 4616
rect 27988 4607 28040 4616
rect 27988 4573 27997 4607
rect 27997 4573 28031 4607
rect 28031 4573 28040 4607
rect 27988 4564 28040 4573
rect 28540 4564 28592 4616
rect 28908 4564 28960 4616
rect 29276 4564 29328 4616
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 3976 4496 4028 4548
rect 4528 4496 4580 4548
rect 5264 4496 5316 4548
rect 6000 4496 6052 4548
rect 6368 4496 6420 4548
rect 10048 4539 10100 4548
rect 5908 4428 5960 4480
rect 6184 4428 6236 4480
rect 10048 4505 10057 4539
rect 10057 4505 10091 4539
rect 10091 4505 10100 4539
rect 10048 4496 10100 4505
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 12348 4496 12400 4548
rect 14832 4428 14884 4480
rect 17132 4496 17184 4548
rect 18788 4496 18840 4548
rect 18972 4496 19024 4548
rect 19984 4496 20036 4548
rect 20996 4496 21048 4548
rect 22008 4496 22060 4548
rect 18052 4428 18104 4480
rect 19340 4428 19392 4480
rect 21088 4428 21140 4480
rect 22100 4428 22152 4480
rect 24032 4496 24084 4548
rect 24676 4539 24728 4548
rect 24676 4505 24685 4539
rect 24685 4505 24719 4539
rect 24719 4505 24728 4539
rect 24676 4496 24728 4505
rect 23848 4471 23900 4480
rect 23848 4437 23857 4471
rect 23857 4437 23891 4471
rect 23891 4437 23900 4471
rect 23848 4428 23900 4437
rect 26516 4496 26568 4548
rect 26148 4471 26200 4480
rect 26148 4437 26157 4471
rect 26157 4437 26191 4471
rect 26191 4437 26200 4471
rect 26148 4428 26200 4437
rect 26240 4428 26292 4480
rect 27528 4496 27580 4548
rect 26792 4471 26844 4480
rect 26792 4437 26801 4471
rect 26801 4437 26835 4471
rect 26835 4437 26844 4471
rect 26792 4428 26844 4437
rect 26884 4428 26936 4480
rect 28080 4471 28132 4480
rect 28080 4437 28089 4471
rect 28089 4437 28123 4471
rect 28123 4437 28132 4471
rect 28080 4428 28132 4437
rect 28264 4496 28316 4548
rect 30748 4564 30800 4616
rect 31208 4564 31260 4616
rect 31668 4607 31720 4616
rect 31668 4573 31677 4607
rect 31677 4573 31711 4607
rect 31711 4573 31720 4607
rect 31668 4564 31720 4573
rect 32496 4607 32548 4616
rect 32496 4573 32505 4607
rect 32505 4573 32539 4607
rect 32539 4573 32548 4607
rect 32496 4564 32548 4573
rect 33784 4607 33836 4616
rect 33784 4573 33793 4607
rect 33793 4573 33827 4607
rect 33827 4573 33836 4607
rect 33784 4564 33836 4573
rect 38016 4607 38068 4616
rect 38016 4573 38025 4607
rect 38025 4573 38059 4607
rect 38059 4573 38068 4607
rect 38016 4564 38068 4573
rect 31116 4539 31168 4548
rect 31116 4505 31125 4539
rect 31125 4505 31159 4539
rect 31159 4505 31168 4539
rect 31116 4496 31168 4505
rect 29920 4428 29972 4480
rect 30472 4471 30524 4480
rect 30472 4437 30481 4471
rect 30481 4437 30515 4471
rect 30515 4437 30524 4471
rect 30472 4428 30524 4437
rect 30656 4428 30708 4480
rect 38200 4471 38252 4480
rect 38200 4437 38209 4471
rect 38209 4437 38243 4471
rect 38243 4437 38252 4471
rect 38200 4428 38252 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4804 4224 4856 4276
rect 9220 4224 9272 4276
rect 4252 4156 4304 4208
rect 4528 4199 4580 4208
rect 4528 4165 4537 4199
rect 4537 4165 4571 4199
rect 4571 4165 4580 4199
rect 4528 4156 4580 4165
rect 5816 4156 5868 4208
rect 5908 4156 5960 4208
rect 7104 4156 7156 4208
rect 26148 4224 26200 4276
rect 26240 4224 26292 4276
rect 29000 4224 29052 4276
rect 29460 4224 29512 4276
rect 9772 4156 9824 4208
rect 10968 4156 11020 4208
rect 13268 4156 13320 4208
rect 14924 4156 14976 4208
rect 16396 4156 16448 4208
rect 17132 4199 17184 4208
rect 17132 4165 17141 4199
rect 17141 4165 17175 4199
rect 17175 4165 17184 4199
rect 17132 4156 17184 4165
rect 19340 4156 19392 4208
rect 19432 4199 19484 4208
rect 19432 4165 19441 4199
rect 19441 4165 19475 4199
rect 19475 4165 19484 4199
rect 19432 4156 19484 4165
rect 20168 4156 20220 4208
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 3424 4020 3476 4072
rect 4068 4020 4120 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8208 4020 8260 4072
rect 10140 4020 10192 4072
rect 11336 4020 11388 4072
rect 11980 4063 12032 4072
rect 3700 3884 3752 3936
rect 3884 3884 3936 3936
rect 4896 3884 4948 3936
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 11060 3952 11112 4004
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 12624 4020 12676 4072
rect 13544 4020 13596 4072
rect 13728 4063 13780 4072
rect 13728 4029 13737 4063
rect 13737 4029 13771 4063
rect 13771 4029 13780 4063
rect 13728 4020 13780 4029
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 16856 4063 16908 4072
rect 16856 4029 16865 4063
rect 16865 4029 16899 4063
rect 16899 4029 16908 4063
rect 16856 4020 16908 4029
rect 18972 4020 19024 4072
rect 19064 4020 19116 4072
rect 22100 4156 22152 4208
rect 21364 4088 21416 4140
rect 23020 4020 23072 4072
rect 8300 3884 8352 3893
rect 10048 3884 10100 3936
rect 13084 3884 13136 3936
rect 18604 3927 18656 3936
rect 18604 3893 18613 3927
rect 18613 3893 18647 3927
rect 18647 3893 18656 3927
rect 18604 3884 18656 3893
rect 20444 3884 20496 3936
rect 20536 3884 20588 3936
rect 22652 3952 22704 4004
rect 26792 4156 26844 4208
rect 24952 4088 25004 4140
rect 25044 4131 25096 4140
rect 25044 4097 25053 4131
rect 25053 4097 25087 4131
rect 25087 4097 25096 4131
rect 25044 4088 25096 4097
rect 25596 4088 25648 4140
rect 27436 4156 27488 4208
rect 28540 4156 28592 4208
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 27804 4131 27856 4140
rect 27804 4097 27813 4131
rect 27813 4097 27847 4131
rect 27847 4097 27856 4131
rect 27804 4088 27856 4097
rect 27988 4088 28040 4140
rect 28908 4088 28960 4140
rect 29092 4131 29144 4140
rect 29092 4097 29101 4131
rect 29101 4097 29135 4131
rect 29135 4097 29144 4131
rect 29092 4088 29144 4097
rect 23388 4063 23440 4072
rect 23388 4029 23397 4063
rect 23397 4029 23431 4063
rect 23431 4029 23440 4063
rect 23388 4020 23440 4029
rect 23940 4063 23992 4072
rect 23940 4029 23949 4063
rect 23949 4029 23983 4063
rect 23983 4029 23992 4063
rect 23940 4020 23992 4029
rect 28356 4020 28408 4072
rect 31668 4156 31720 4208
rect 29276 4088 29328 4140
rect 29644 4020 29696 4072
rect 30564 4088 30616 4140
rect 30748 4088 30800 4140
rect 31576 4088 31628 4140
rect 32404 4088 32456 4140
rect 31116 4020 31168 4072
rect 38292 4131 38344 4140
rect 24860 3952 24912 4004
rect 25320 3952 25372 4004
rect 29276 3952 29328 4004
rect 33048 4020 33100 4072
rect 38292 4097 38301 4131
rect 38301 4097 38335 4131
rect 38335 4097 38344 4131
rect 38292 4088 38344 4097
rect 21364 3884 21416 3936
rect 22376 3884 22428 3936
rect 22560 3884 22612 3936
rect 23940 3884 23992 3936
rect 25228 3884 25280 3936
rect 26516 3927 26568 3936
rect 26516 3893 26525 3927
rect 26525 3893 26559 3927
rect 26559 3893 26568 3927
rect 26516 3884 26568 3893
rect 26792 3884 26844 3936
rect 27620 3884 27672 3936
rect 28356 3884 28408 3936
rect 28540 3927 28592 3936
rect 28540 3893 28549 3927
rect 28549 3893 28583 3927
rect 28583 3893 28592 3927
rect 28540 3884 28592 3893
rect 29368 3884 29420 3936
rect 30564 3884 30616 3936
rect 31300 3884 31352 3936
rect 35808 3952 35860 4004
rect 33048 3927 33100 3936
rect 33048 3893 33057 3927
rect 33057 3893 33091 3927
rect 33091 3893 33100 3927
rect 33048 3884 33100 3893
rect 35716 3884 35768 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3148 3680 3200 3732
rect 2044 3544 2096 3596
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 4988 3680 5040 3732
rect 6828 3680 6880 3732
rect 7104 3680 7156 3732
rect 9404 3680 9456 3732
rect 8484 3612 8536 3664
rect 11888 3680 11940 3732
rect 11060 3612 11112 3664
rect 12808 3680 12860 3732
rect 12900 3680 12952 3732
rect 13728 3612 13780 3664
rect 6552 3544 6604 3596
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 10784 3544 10836 3596
rect 14556 3544 14608 3596
rect 17776 3612 17828 3664
rect 16580 3544 16632 3596
rect 16672 3544 16724 3596
rect 4804 3408 4856 3460
rect 4896 3451 4948 3460
rect 4896 3417 4905 3451
rect 4905 3417 4939 3451
rect 4939 3417 4948 3451
rect 4896 3408 4948 3417
rect 6828 3408 6880 3460
rect 7012 3408 7064 3460
rect 7196 3408 7248 3460
rect 5264 3340 5316 3392
rect 5540 3340 5592 3392
rect 8484 3340 8536 3392
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 9128 3383 9180 3392
rect 8576 3340 8628 3349
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 14740 3476 14792 3528
rect 17776 3476 17828 3528
rect 9404 3408 9456 3460
rect 10140 3408 10192 3460
rect 12164 3408 12216 3460
rect 12532 3408 12584 3460
rect 13544 3408 13596 3460
rect 16120 3451 16172 3460
rect 10876 3340 10928 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 16120 3417 16129 3451
rect 16129 3417 16163 3451
rect 16163 3417 16172 3451
rect 16120 3408 16172 3417
rect 17960 3408 18012 3460
rect 20996 3680 21048 3732
rect 19156 3544 19208 3596
rect 28540 3680 28592 3732
rect 28724 3680 28776 3732
rect 29644 3680 29696 3732
rect 29828 3723 29880 3732
rect 29828 3689 29837 3723
rect 29837 3689 29871 3723
rect 29871 3689 29880 3723
rect 29828 3680 29880 3689
rect 30380 3680 30432 3732
rect 36728 3723 36780 3732
rect 36728 3689 36737 3723
rect 36737 3689 36771 3723
rect 36771 3689 36780 3723
rect 36728 3680 36780 3689
rect 21272 3612 21324 3664
rect 24952 3612 25004 3664
rect 25688 3612 25740 3664
rect 29276 3612 29328 3664
rect 30656 3612 30708 3664
rect 23848 3544 23900 3596
rect 23940 3544 23992 3596
rect 28540 3544 28592 3596
rect 28908 3544 28960 3596
rect 21180 3476 21232 3528
rect 19432 3408 19484 3460
rect 19984 3408 20036 3460
rect 13728 3340 13780 3349
rect 18144 3340 18196 3392
rect 24492 3476 24544 3528
rect 23296 3408 23348 3460
rect 24308 3340 24360 3392
rect 24768 3451 24820 3460
rect 24768 3417 24777 3451
rect 24777 3417 24811 3451
rect 24811 3417 24820 3451
rect 24768 3408 24820 3417
rect 26148 3476 26200 3528
rect 26332 3519 26384 3528
rect 26332 3485 26341 3519
rect 26341 3485 26375 3519
rect 26375 3485 26384 3519
rect 26332 3476 26384 3485
rect 26424 3476 26476 3528
rect 26884 3476 26936 3528
rect 28264 3476 28316 3528
rect 28448 3476 28500 3528
rect 28724 3476 28776 3528
rect 29092 3476 29144 3528
rect 32772 3544 32824 3596
rect 31208 3476 31260 3528
rect 31392 3476 31444 3528
rect 32496 3519 32548 3528
rect 32496 3485 32505 3519
rect 32505 3485 32539 3519
rect 32539 3485 32548 3519
rect 32496 3476 32548 3485
rect 32588 3476 32640 3528
rect 34704 3476 34756 3528
rect 35716 3519 35768 3528
rect 35716 3485 35725 3519
rect 35725 3485 35759 3519
rect 35759 3485 35768 3519
rect 35716 3476 35768 3485
rect 37372 3476 37424 3528
rect 37924 3476 37976 3528
rect 25964 3408 26016 3460
rect 25596 3340 25648 3392
rect 26148 3383 26200 3392
rect 26148 3349 26157 3383
rect 26157 3349 26191 3383
rect 26191 3349 26200 3383
rect 26148 3340 26200 3349
rect 26424 3340 26476 3392
rect 28172 3340 28224 3392
rect 28816 3340 28868 3392
rect 30748 3340 30800 3392
rect 31116 3383 31168 3392
rect 31116 3349 31125 3383
rect 31125 3349 31159 3383
rect 31159 3349 31168 3383
rect 31116 3340 31168 3349
rect 31208 3340 31260 3392
rect 34428 3408 34480 3460
rect 33600 3383 33652 3392
rect 33600 3349 33609 3383
rect 33609 3349 33643 3383
rect 33643 3349 33652 3383
rect 33600 3340 33652 3349
rect 33692 3340 33744 3392
rect 36636 3340 36688 3392
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5540 3136 5592 3188
rect 5816 3136 5868 3188
rect 3976 3068 4028 3120
rect 6828 3068 6880 3120
rect 8116 3068 8168 3120
rect 8576 3111 8628 3120
rect 8576 3077 8585 3111
rect 8585 3077 8619 3111
rect 8619 3077 8628 3111
rect 8576 3068 8628 3077
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 1676 2932 1728 2984
rect 4068 2932 4120 2984
rect 5264 2932 5316 2984
rect 3792 2907 3844 2916
rect 3792 2873 3801 2907
rect 3801 2873 3835 2907
rect 3835 2873 3844 2907
rect 3792 2864 3844 2873
rect 3608 2796 3660 2848
rect 6920 2932 6972 2984
rect 9312 3000 9364 3052
rect 9588 3068 9640 3120
rect 9956 3068 10008 3120
rect 10968 3068 11020 3120
rect 11888 3068 11940 3120
rect 12624 3111 12676 3120
rect 12624 3077 12633 3111
rect 12633 3077 12667 3111
rect 12667 3077 12676 3111
rect 12624 3068 12676 3077
rect 11612 3000 11664 3052
rect 13728 3000 13780 3052
rect 5632 2796 5684 2848
rect 10692 2932 10744 2984
rect 10876 2932 10928 2984
rect 12348 2975 12400 2984
rect 11612 2864 11664 2916
rect 9496 2796 9548 2848
rect 12348 2941 12357 2975
rect 12357 2941 12391 2975
rect 12391 2941 12400 2975
rect 12348 2932 12400 2941
rect 12624 2932 12676 2984
rect 14464 3068 14516 3120
rect 16488 3068 16540 3120
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 16028 2932 16080 2984
rect 16304 2975 16356 2984
rect 16304 2941 16313 2975
rect 16313 2941 16347 2975
rect 16347 2941 16356 2975
rect 16304 2932 16356 2941
rect 13360 2796 13412 2848
rect 14924 2796 14976 2848
rect 17776 3136 17828 3188
rect 19892 3136 19944 3188
rect 26424 3136 26476 3188
rect 21916 3068 21968 3120
rect 25320 3068 25372 3120
rect 25596 3111 25648 3120
rect 25596 3077 25605 3111
rect 25605 3077 25639 3111
rect 25639 3077 25648 3111
rect 25596 3068 25648 3077
rect 25688 3111 25740 3120
rect 25688 3077 25697 3111
rect 25697 3077 25731 3111
rect 25731 3077 25740 3111
rect 26608 3111 26660 3120
rect 25688 3068 25740 3077
rect 26608 3077 26617 3111
rect 26617 3077 26651 3111
rect 26651 3077 26660 3111
rect 26608 3068 26660 3077
rect 33048 3136 33100 3188
rect 34336 3179 34388 3188
rect 34336 3145 34345 3179
rect 34345 3145 34379 3179
rect 34379 3145 34388 3179
rect 34336 3136 34388 3145
rect 35624 3179 35676 3188
rect 35624 3145 35633 3179
rect 35633 3145 35667 3179
rect 35667 3145 35676 3179
rect 35624 3136 35676 3145
rect 27436 3068 27488 3120
rect 16856 3000 16908 3052
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 19156 3000 19208 3052
rect 23848 3043 23900 3052
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 24584 3000 24636 3052
rect 28540 3043 28592 3052
rect 28540 3009 28549 3043
rect 28549 3009 28583 3043
rect 28583 3009 28592 3043
rect 28540 3000 28592 3009
rect 33692 3068 33744 3120
rect 19064 2932 19116 2984
rect 20996 2932 21048 2984
rect 22376 2975 22428 2984
rect 21364 2864 21416 2916
rect 18420 2796 18472 2848
rect 21916 2864 21968 2916
rect 22376 2941 22385 2975
rect 22385 2941 22419 2975
rect 22419 2941 22428 2975
rect 22376 2932 22428 2941
rect 22652 2975 22704 2984
rect 22652 2941 22661 2975
rect 22661 2941 22695 2975
rect 22695 2941 22704 2975
rect 22652 2932 22704 2941
rect 25872 2932 25924 2984
rect 27252 2975 27304 2984
rect 27252 2941 27261 2975
rect 27261 2941 27295 2975
rect 27295 2941 27304 2975
rect 27252 2932 27304 2941
rect 29736 2975 29788 2984
rect 23940 2907 23992 2916
rect 23940 2873 23949 2907
rect 23949 2873 23983 2907
rect 23983 2873 23992 2907
rect 23940 2864 23992 2873
rect 24308 2864 24360 2916
rect 25044 2864 25096 2916
rect 27620 2864 27672 2916
rect 27896 2864 27948 2916
rect 29736 2941 29745 2975
rect 29745 2941 29779 2975
rect 29779 2941 29788 2975
rect 29736 2932 29788 2941
rect 30840 3000 30892 3052
rect 31208 2932 31260 2984
rect 31668 3000 31720 3052
rect 32772 3000 32824 3052
rect 29092 2864 29144 2916
rect 30748 2864 30800 2916
rect 28172 2796 28224 2848
rect 28724 2796 28776 2848
rect 33140 2932 33192 2984
rect 34428 3000 34480 3052
rect 35532 3043 35584 3052
rect 35532 3009 35541 3043
rect 35541 3009 35575 3043
rect 35575 3009 35584 3043
rect 35532 3000 35584 3009
rect 35440 2932 35492 2984
rect 36636 3000 36688 3052
rect 33232 2864 33284 2916
rect 31668 2839 31720 2848
rect 31668 2805 31677 2839
rect 31677 2805 31711 2839
rect 31711 2805 31720 2839
rect 31668 2796 31720 2805
rect 32404 2839 32456 2848
rect 32404 2805 32413 2839
rect 32413 2805 32447 2839
rect 32447 2805 32456 2839
rect 32404 2796 32456 2805
rect 32864 2796 32916 2848
rect 34520 2796 34572 2848
rect 36176 2839 36228 2848
rect 36176 2805 36185 2839
rect 36185 2805 36219 2839
rect 36219 2805 36228 2839
rect 36176 2796 36228 2805
rect 38660 2796 38712 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3424 2635 3476 2644
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 5632 2592 5684 2644
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 3792 2456 3844 2508
rect 4068 2456 4120 2508
rect 6552 2456 6604 2508
rect 13636 2592 13688 2644
rect 15476 2592 15528 2644
rect 19432 2592 19484 2644
rect 19524 2592 19576 2644
rect 21180 2635 21232 2644
rect 21180 2601 21189 2635
rect 21189 2601 21223 2635
rect 21223 2601 21232 2635
rect 21180 2592 21232 2601
rect 11888 2524 11940 2576
rect 18420 2524 18472 2576
rect 9772 2456 9824 2508
rect 12348 2456 12400 2508
rect 14556 2499 14608 2508
rect 14556 2465 14565 2499
rect 14565 2465 14599 2499
rect 14599 2465 14608 2499
rect 14556 2456 14608 2465
rect 16028 2456 16080 2508
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 19156 2456 19208 2508
rect 23480 2592 23532 2644
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 24860 2592 24912 2644
rect 26332 2592 26384 2644
rect 22652 2499 22704 2508
rect 22652 2465 22661 2499
rect 22661 2465 22695 2499
rect 22695 2465 22704 2499
rect 22652 2456 22704 2465
rect 4068 2320 4120 2372
rect 5908 2320 5960 2372
rect 5816 2252 5868 2304
rect 8944 2320 8996 2372
rect 9956 2320 10008 2372
rect 12164 2320 12216 2372
rect 10600 2252 10652 2304
rect 13728 2320 13780 2372
rect 17316 2320 17368 2372
rect 22192 2388 22244 2440
rect 23296 2388 23348 2440
rect 24768 2431 24820 2440
rect 24768 2397 24777 2431
rect 24777 2397 24811 2431
rect 24811 2397 24820 2431
rect 24768 2388 24820 2397
rect 27896 2456 27948 2508
rect 28632 2456 28684 2508
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 26148 2388 26200 2440
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 27712 2388 27764 2440
rect 29000 2388 29052 2440
rect 22468 2363 22520 2372
rect 16120 2252 16172 2304
rect 16304 2295 16356 2304
rect 16304 2261 16313 2295
rect 16313 2261 16347 2295
rect 16347 2261 16356 2295
rect 16304 2252 16356 2261
rect 19524 2252 19576 2304
rect 22468 2329 22477 2363
rect 22477 2329 22511 2363
rect 22511 2329 22520 2363
rect 22468 2320 22520 2329
rect 32128 2592 32180 2644
rect 37188 2524 37240 2576
rect 34612 2456 34664 2508
rect 32312 2431 32364 2440
rect 32312 2397 32321 2431
rect 32321 2397 32355 2431
rect 32355 2397 32364 2431
rect 32312 2388 32364 2397
rect 33508 2388 33560 2440
rect 34796 2388 34848 2440
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 35900 2388 35952 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 33048 2320 33100 2372
rect 25780 2252 25832 2304
rect 26148 2252 26200 2304
rect 29552 2252 29604 2304
rect 30288 2252 30340 2304
rect 32220 2252 32272 2304
rect 33508 2252 33560 2304
rect 34152 2252 34204 2304
rect 36728 2252 36780 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 2780 2048 2832 2100
rect 4712 2048 4764 2100
rect 22468 2048 22520 2100
rect 26792 2048 26844 2100
rect 17316 1980 17368 2032
rect 13636 1912 13688 1964
rect 23664 1912 23716 1964
rect 24768 1980 24820 2032
rect 30840 1980 30892 2032
rect 31116 1912 31168 1964
rect 17960 1844 18012 1896
rect 29092 1844 29144 1896
rect 9956 1776 10008 1828
rect 18880 1776 18932 1828
rect 20996 1776 21048 1828
rect 11796 1708 11848 1760
rect 18420 1708 18472 1760
rect 16304 1640 16356 1692
rect 27804 1708 27856 1760
rect 19984 1640 20036 1692
rect 27344 1640 27396 1692
rect 36176 1640 36228 1692
rect 23204 1572 23256 1624
rect 27436 1572 27488 1624
rect 21272 1504 21324 1556
rect 23296 1504 23348 1556
rect 12164 1436 12216 1488
rect 25228 1436 25280 1488
rect 21180 1368 21232 1420
rect 25136 1368 25188 1420
rect 20444 1300 20496 1352
rect 31392 1300 31444 1352
rect 10968 1232 11020 1284
rect 34520 1232 34572 1284
rect 13268 1164 13320 1216
rect 29276 1164 29328 1216
rect 16396 1096 16448 1148
rect 32404 1096 32456 1148
rect 11980 1028 12032 1080
rect 27160 1028 27212 1080
rect 4068 960 4120 1012
rect 31668 960 31720 1012
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2594 39200 2650 39800
rect 3146 39536 3202 39545
rect 3146 39471 3202 39480
rect 676 35698 704 39200
rect 1582 38856 1638 38865
rect 1582 38791 1638 38800
rect 1596 37330 1624 38791
rect 1766 37496 1822 37505
rect 1766 37431 1822 37440
rect 1584 37324 1636 37330
rect 1584 37266 1636 37272
rect 1780 36922 1808 37431
rect 1860 37256 1912 37262
rect 1860 37198 1912 37204
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1768 36168 1820 36174
rect 1766 36136 1768 36145
rect 1820 36136 1822 36145
rect 1766 36071 1822 36080
rect 1872 35894 1900 37198
rect 1964 36786 1992 39200
rect 2608 37244 2636 39200
rect 2780 37256 2832 37262
rect 2608 37216 2780 37244
rect 2780 37198 2832 37204
rect 3160 36786 3188 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 5814 39200 5870 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 16118 39200 16174 39800
rect 16224 39222 16528 39250
rect 3896 37330 3924 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3884 37324 3936 37330
rect 3884 37266 3936 37272
rect 5184 37262 5212 39200
rect 5828 37330 5856 39200
rect 5816 37324 5868 37330
rect 5816 37266 5868 37272
rect 7116 37262 7144 39200
rect 8404 37330 8432 39200
rect 8392 37324 8444 37330
rect 8392 37266 8444 37272
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 6828 37256 6880 37262
rect 6828 37198 6880 37204
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 4264 36922 4292 37198
rect 5264 37120 5316 37126
rect 5264 37062 5316 37068
rect 4252 36916 4304 36922
rect 4252 36858 4304 36864
rect 1952 36780 2004 36786
rect 1952 36722 2004 36728
rect 3148 36780 3200 36786
rect 3148 36722 3200 36728
rect 4620 36712 4672 36718
rect 4620 36654 4672 36660
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2688 36032 2740 36038
rect 2688 35974 2740 35980
rect 1872 35866 1992 35894
rect 664 35692 716 35698
rect 664 35634 716 35640
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1596 30122 1624 34546
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34105 1808 34342
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 1768 32768 1820 32774
rect 1766 32736 1768 32745
rect 1820 32736 1822 32745
rect 1766 32671 1822 32680
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1766 30696 1822 30705
rect 1766 30631 1822 30640
rect 1780 30598 1808 30631
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1584 30116 1636 30122
rect 1584 30058 1636 30064
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1780 29345 1808 29582
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1768 29028 1820 29034
rect 1768 28970 1820 28976
rect 1780 28665 1808 28970
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 27305 1808 27406
rect 1766 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1780 25945 1808 26318
rect 1766 25936 1822 25945
rect 1766 25871 1822 25880
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1596 24410 1624 24754
rect 1768 24608 1820 24614
rect 1766 24576 1768 24585
rect 1820 24576 1822 24585
rect 1766 24511 1822 24520
rect 1584 24404 1636 24410
rect 1584 24346 1636 24352
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1766 23831 1822 23840
rect 1964 23118 1992 35866
rect 2596 32428 2648 32434
rect 2596 32370 2648 32376
rect 2320 29164 2372 29170
rect 2320 29106 2372 29112
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1688 22545 1716 22578
rect 1674 22536 1730 22545
rect 1674 22471 1730 22480
rect 1768 22432 1820 22438
rect 1768 22374 1820 22380
rect 1780 22234 1808 22374
rect 1768 22228 1820 22234
rect 1768 22170 1820 22176
rect 1964 22030 1992 23054
rect 2332 22778 2360 29106
rect 2608 26858 2636 32370
rect 2700 30734 2728 35974
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 33658 4660 36654
rect 4620 33652 4672 33658
rect 4620 33594 4672 33600
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3424 32292 3476 32298
rect 3424 32234 3476 32240
rect 2688 30728 2740 30734
rect 2688 30670 2740 30676
rect 2596 26852 2648 26858
rect 2596 26794 2648 26800
rect 3436 25430 3464 32234
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 5276 29714 5304 37062
rect 6736 36644 6788 36650
rect 6736 36586 6788 36592
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5264 29708 5316 29714
rect 5264 29650 5316 29656
rect 5552 29594 5580 32846
rect 5736 31346 5764 35430
rect 5828 31822 5856 36518
rect 6644 33516 6696 33522
rect 6644 33458 6696 33464
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 6000 30252 6052 30258
rect 6000 30194 6052 30200
rect 5552 29566 5764 29594
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 2688 25424 2740 25430
rect 2688 25366 2740 25372
rect 3424 25424 3476 25430
rect 3424 25366 3476 25372
rect 2700 24206 2728 25366
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2320 22772 2372 22778
rect 2320 22714 2372 22720
rect 4080 22710 4108 27270
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 5540 26512 5592 26518
rect 5540 26454 5592 26460
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 5552 23730 5580 26454
rect 5644 24818 5672 29446
rect 5736 26382 5764 29566
rect 6012 27130 6040 30194
rect 6000 27124 6052 27130
rect 6000 27066 6052 27072
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2516 22545 2544 22578
rect 2502 22536 2558 22545
rect 2502 22471 2504 22480
rect 2556 22471 2558 22480
rect 2504 22442 2556 22448
rect 2516 22411 2544 22442
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1596 21554 1624 21830
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1780 21185 1808 21286
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 1766 21176 1822 21185
rect 4214 21179 4522 21188
rect 1766 21111 1822 21120
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1780 19145 1808 19314
rect 4712 19168 4764 19174
rect 1766 19136 1822 19145
rect 4712 19110 4764 19116
rect 1766 19071 1822 19080
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4724 18766 4752 19110
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18358 4384 18566
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17785 1808 18226
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 1766 17776 1822 17785
rect 4632 17746 4660 18158
rect 1766 17711 1822 17720
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1872 17202 1900 17546
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 3700 17196 3752 17202
rect 3700 17138 3752 17144
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 1584 17128 1636 17134
rect 1582 17096 1584 17105
rect 1636 17096 1638 17105
rect 1582 17031 1638 17040
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2700 16250 2728 16526
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 1582 16144 1638 16153
rect 1582 16079 1584 16088
rect 1636 16079 1638 16088
rect 1584 16050 1636 16056
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 15337 2176 15438
rect 2134 15328 2190 15337
rect 2134 15263 2190 15272
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1780 14278 1808 14311
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1768 13728 1820 13734
rect 1766 13696 1768 13705
rect 1820 13696 1822 13705
rect 1766 13631 1822 13640
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 11626 1624 12786
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12345 1808 12582
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1584 11620 1636 11626
rect 1584 11562 1636 11568
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1596 10985 1624 11086
rect 1582 10976 1638 10985
rect 1582 10911 1638 10920
rect 1582 10840 1638 10849
rect 1582 10775 1638 10784
rect 1596 10674 1624 10775
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1780 10305 1808 11698
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1872 9518 1900 13194
rect 1964 12442 1992 13194
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10266 1992 10542
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1964 9654 1992 9998
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 2056 8974 2084 10406
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6905 1624 7278
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 20 5568 72 5574
rect 20 5510 72 5516
rect 32 800 60 5510
rect 1596 5234 1624 6598
rect 1688 6322 1716 7686
rect 1872 7410 1900 8191
rect 2056 7886 2084 8774
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 664 5024 716 5030
rect 664 4966 716 4972
rect 676 800 704 4966
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1688 4078 1716 4558
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1688 3534 1716 4014
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 2990 1716 3470
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2514 1716 2926
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1964 800 1992 7346
rect 2148 7274 2176 12174
rect 2240 7342 2268 15914
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2412 15020 2464 15026
rect 2412 14962 2464 14968
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6254 2268 6734
rect 2332 6322 2360 8298
rect 2424 8090 2452 14962
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 11830 2544 14350
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2516 10266 2544 10542
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2516 5710 2544 6598
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2608 5234 2636 14758
rect 2700 13938 2728 15438
rect 2792 14482 2820 16390
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2884 14346 2912 16390
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2686 13016 2742 13025
rect 2686 12951 2742 12960
rect 2700 11218 2728 12951
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2792 11898 2820 12786
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2884 12306 2912 12582
rect 2976 12434 3004 14758
rect 3068 14006 3096 15846
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 2976 12406 3096 12434
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10674 2820 10950
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2700 9722 2728 9998
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 8401 2728 8434
rect 2686 8392 2742 8401
rect 2686 8327 2742 8336
rect 2792 8344 2820 9522
rect 2872 8968 2924 8974
rect 2870 8936 2872 8945
rect 2924 8936 2926 8945
rect 2870 8871 2926 8880
rect 2792 8316 2912 8344
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 7585 2820 7822
rect 2778 7576 2834 7585
rect 2884 7546 2912 8316
rect 2778 7511 2834 7520
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2792 4185 2820 6122
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 2042 3632 2098 3641
rect 2042 3567 2044 3576
rect 2096 3567 2098 3576
rect 2044 3538 2096 3544
rect 2056 3369 2084 3538
rect 2884 3505 2912 6054
rect 2976 5545 3004 9998
rect 3068 9654 3096 12406
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10266 3188 10610
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3252 9602 3280 15302
rect 3344 14006 3372 16934
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3436 11914 3464 16390
rect 3712 16046 3740 17138
rect 4172 17105 4200 17138
rect 4158 17096 4214 17105
rect 4158 17031 4214 17040
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3528 13870 3556 14282
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 12050 3556 12582
rect 3620 12186 3648 14894
rect 3712 12434 3740 15982
rect 3988 15638 4016 16050
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3804 13530 3832 14962
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3804 12850 3832 13466
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3712 12406 3832 12434
rect 3620 12158 3740 12186
rect 3528 12022 3648 12050
rect 3436 11886 3556 11914
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3436 11354 3464 11698
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3148 9580 3200 9586
rect 3252 9574 3464 9602
rect 3148 9522 3200 9528
rect 3160 9042 3188 9522
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9110 3280 9318
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 6798 3096 8774
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3160 7750 3188 8502
rect 3344 7970 3372 9454
rect 3252 7942 3372 7970
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3252 6882 3280 7942
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3160 6854 3280 6882
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3160 5914 3188 6854
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2962 5536 3018 5545
rect 2962 5471 3018 5480
rect 3160 3738 3188 5850
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2042 3360 2098 3369
rect 2042 3295 2098 3304
rect 2778 2136 2834 2145
rect 2778 2071 2780 2080
rect 2832 2071 2834 2080
rect 2780 2042 2832 2048
rect 3252 800 3280 6666
rect 3344 921 3372 7822
rect 3436 6458 3464 9574
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3528 4554 3556 11886
rect 3620 8634 3648 12022
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3606 6352 3662 6361
rect 3606 6287 3608 6296
rect 3660 6287 3662 6296
rect 3608 6258 3660 6264
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3436 2650 3464 4014
rect 3620 2854 3648 4694
rect 3712 3942 3740 12158
rect 3804 10062 3832 12406
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 7410 3832 9862
rect 3896 8974 3924 13806
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 12986 4016 13670
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 4080 11762 4108 16118
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 16050
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4264 15094 4292 15438
rect 4344 15360 4396 15366
rect 4342 15328 4344 15337
rect 4396 15328 4398 15337
rect 4342 15263 4398 15272
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14657 4660 14758
rect 4618 14648 4674 14657
rect 4528 14612 4580 14618
rect 4618 14583 4674 14592
rect 4528 14554 4580 14560
rect 4540 13938 4568 14554
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4158 11112 4214 11121
rect 4158 11047 4214 11056
rect 4172 10452 4200 11047
rect 4632 10810 4660 14418
rect 4724 14346 4752 16934
rect 4804 16584 4856 16590
rect 4908 16561 4936 18158
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4804 16526 4856 16532
rect 4894 16552 4950 16561
rect 4816 15502 4844 16526
rect 4894 16487 4950 16496
rect 4908 15910 4936 16487
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 5000 15706 5028 17138
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4804 15496 4856 15502
rect 4856 15456 4936 15484
rect 4804 15438 4856 15444
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4724 12850 4752 13874
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4724 12753 4752 12786
rect 4710 12744 4766 12753
rect 4710 12679 4766 12688
rect 4712 12640 4764 12646
rect 4710 12608 4712 12617
rect 4764 12608 4766 12617
rect 4710 12543 4766 12552
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 3988 10424 4200 10452
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3988 8090 4016 10424
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7410 3924 7686
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3988 6866 4016 7822
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3882 6760 3938 6769
rect 3882 6695 3938 6704
rect 3896 5778 3924 6695
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3988 5710 4016 6258
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4080 5250 4108 9998
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 10610
rect 4710 10432 4766 10441
rect 4710 10367 4766 10376
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4724 9058 4752 10367
rect 4632 9030 4752 9058
rect 4632 8566 4660 9030
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8230
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4264 6322 4292 6802
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4526 6624 4582 6633
rect 4526 6559 4582 6568
rect 4540 6390 4568 6559
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 3896 5222 4108 5250
rect 4264 5234 4292 5578
rect 4252 5228 4304 5234
rect 3896 4758 3924 5222
rect 4252 5170 4304 5176
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 4080 4570 4108 5102
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3988 4554 4108 4570
rect 3976 4548 4108 4554
rect 4028 4542 4108 4548
rect 3976 4490 4028 4496
rect 4080 4078 4108 4542
rect 4264 4214 4292 4762
rect 4526 4720 4582 4729
rect 4526 4655 4582 4664
rect 4540 4554 4568 4655
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4526 4312 4582 4321
rect 4526 4247 4582 4256
rect 4540 4214 4568 4247
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4068 4072 4120 4078
rect 3790 4040 3846 4049
rect 4068 4014 4120 4020
rect 3790 3975 3846 3984
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3804 2922 3832 3975
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3804 2514 3832 2858
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3330 912 3386 921
rect 3330 847 3386 856
rect 3896 800 3924 3878
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3988 1737 4016 3062
rect 4080 2990 4108 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4080 2514 4108 2926
rect 4632 2774 4660 6666
rect 4724 6662 4752 8910
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4816 5642 4844 14010
rect 4908 13938 4936 15456
rect 5092 15434 5120 16390
rect 5080 15428 5132 15434
rect 5080 15370 5132 15376
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4908 12730 4936 13670
rect 5000 12850 5028 14826
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4908 12702 5028 12730
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 10169 4936 12582
rect 5000 12306 5028 12702
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5092 11354 5120 13806
rect 5184 13734 5212 20946
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5276 16561 5304 20810
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6012 18970 6040 19314
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5828 18426 5856 18702
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5262 16552 5318 16561
rect 5262 16487 5318 16496
rect 5460 16182 5488 16934
rect 5736 16658 5764 18226
rect 6104 17610 6132 31078
rect 6656 30326 6684 33458
rect 6644 30320 6696 30326
rect 6644 30262 6696 30268
rect 6748 29646 6776 36586
rect 6840 32910 6868 37198
rect 9048 36786 9076 39200
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 9416 36854 9444 37198
rect 10336 37126 10364 39200
rect 11624 37262 11652 39200
rect 11612 37256 11664 37262
rect 12268 37244 12296 39200
rect 13556 37262 13584 39200
rect 12440 37256 12492 37262
rect 12268 37216 12440 37244
rect 11612 37198 11664 37204
rect 12440 37198 12492 37204
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 11060 37188 11112 37194
rect 11060 37130 11112 37136
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 9404 36848 9456 36854
rect 9404 36790 9456 36796
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 8024 36576 8076 36582
rect 8024 36518 8076 36524
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 8036 30734 8064 36518
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 8208 30592 8260 30598
rect 8208 30534 8260 30540
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 7012 29504 7064 29510
rect 7012 29446 7064 29452
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5828 16794 5856 17138
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10985 5028 11086
rect 4986 10976 5042 10985
rect 4986 10911 5042 10920
rect 4894 10160 4950 10169
rect 4894 10095 4950 10104
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4816 3466 4844 4218
rect 4908 3942 4936 9998
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5000 9654 5028 9862
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4988 9512 5040 9518
rect 4986 9480 4988 9489
rect 5040 9480 5042 9489
rect 4986 9415 5042 9424
rect 4986 9208 5042 9217
rect 4986 9143 4988 9152
rect 5040 9143 5042 9152
rect 4988 9114 5040 9120
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 5000 3738 5028 8774
rect 5184 6390 5212 13126
rect 5276 11937 5304 13942
rect 5368 13734 5396 15982
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5460 14113 5488 14282
rect 5446 14104 5502 14113
rect 5446 14039 5502 14048
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5460 12730 5488 13874
rect 5552 13326 5580 13874
rect 5644 13569 5672 14758
rect 5630 13560 5686 13569
rect 5630 13495 5686 13504
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5552 12850 5580 13262
rect 5644 12918 5672 13262
rect 5632 12912 5684 12918
rect 5632 12854 5684 12860
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5630 12744 5686 12753
rect 5460 12702 5580 12730
rect 5552 12220 5580 12702
rect 5630 12679 5686 12688
rect 5354 12200 5410 12209
rect 5354 12135 5410 12144
rect 5460 12192 5580 12220
rect 5262 11928 5318 11937
rect 5262 11863 5318 11872
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 9926 5304 10950
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5262 9752 5318 9761
rect 5262 9687 5318 9696
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4894 3496 4950 3505
rect 4804 3460 4856 3466
rect 4894 3431 4896 3440
rect 4804 3402 4856 3408
rect 4948 3431 4950 3440
rect 4896 3402 4948 3408
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4632 2746 4752 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 3974 1728 4030 1737
rect 3974 1663 4030 1672
rect 4080 1018 4108 2314
rect 4724 2106 4752 2746
rect 4712 2100 4764 2106
rect 4712 2042 4764 2048
rect 4068 1012 4120 1018
rect 4068 954 4120 960
rect 5184 800 5212 6054
rect 5276 4554 5304 9687
rect 5368 7546 5396 12135
rect 5460 10985 5488 12192
rect 5644 11762 5672 12679
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5446 10976 5502 10985
rect 5446 10911 5502 10920
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5552 7410 5580 11018
rect 5644 10674 5672 11562
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5644 7478 5672 7890
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5368 6458 5396 6666
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5552 5030 5580 7346
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 5098 5672 6598
rect 5736 5710 5764 16594
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 14249 5856 14962
rect 5814 14240 5870 14249
rect 5814 14175 5870 14184
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5828 10810 5856 13194
rect 5920 12238 5948 17478
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 6000 13728 6052 13734
rect 6104 13705 6132 15982
rect 6000 13670 6052 13676
rect 6090 13696 6146 13705
rect 6012 13530 6040 13670
rect 6090 13631 6146 13640
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6104 13297 6132 13631
rect 6196 13530 6224 20198
rect 6932 19786 6960 21286
rect 7024 20534 7052 29446
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 7012 20528 7064 20534
rect 7012 20470 7064 20476
rect 7024 20330 7052 20470
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 7116 19786 7144 26930
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7208 21962 7236 22578
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7300 22030 7328 22374
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6368 16720 6420 16726
rect 6368 16662 6420 16668
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 16182 6316 16390
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6288 14414 6316 15030
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6184 13320 6236 13326
rect 6090 13288 6146 13297
rect 6184 13262 6236 13268
rect 6090 13223 6146 13232
rect 6196 12866 6224 13262
rect 6288 12918 6316 14350
rect 6012 12838 6224 12866
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6012 11778 6040 12838
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6104 12442 6132 12650
rect 6182 12608 6238 12617
rect 6182 12543 6238 12552
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5920 11750 6040 11778
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5920 10690 5948 11750
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5828 10662 5948 10690
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5538 4856 5594 4865
rect 5538 4791 5594 4800
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5552 3618 5580 4791
rect 5828 4214 5856 10662
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 7818 5948 10406
rect 6012 8634 6040 11630
rect 6104 11150 6132 12174
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 6012 8090 6040 8570
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 6104 7206 6132 7958
rect 6196 7818 6224 12543
rect 6288 10674 6316 12854
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9722 6316 9998
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6380 8090 6408 16662
rect 6472 15570 6500 18566
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6564 17678 6592 18022
rect 6748 17882 6776 19654
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6642 17776 6698 17785
rect 6840 17746 6868 19450
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 6932 18290 6960 19314
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6642 17711 6644 17720
rect 6696 17711 6698 17720
rect 6828 17740 6880 17746
rect 6644 17682 6696 17688
rect 6828 17682 6880 17688
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6748 17134 6776 17614
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6550 16688 6606 16697
rect 6550 16623 6552 16632
rect 6604 16623 6606 16632
rect 6552 16594 6604 16600
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6472 12714 6500 13738
rect 6550 13696 6606 13705
rect 6550 13631 6606 13640
rect 6564 12850 6592 13631
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6472 12209 6500 12650
rect 6552 12436 6604 12442
rect 6748 12434 6776 17070
rect 6828 17060 6880 17066
rect 6828 17002 6880 17008
rect 6840 13258 6868 17002
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6932 15337 6960 16050
rect 7116 16046 7144 18566
rect 7208 17270 7236 19314
rect 7300 18834 7328 21830
rect 7392 21554 7420 21830
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7392 19514 7420 20878
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8036 20058 8064 20470
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 7484 18902 7512 19722
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7380 18760 7432 18766
rect 7576 18714 7604 19790
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 7944 19174 7972 19314
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7380 18702 7432 18708
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7196 17264 7248 17270
rect 7196 17206 7248 17212
rect 7300 17082 7328 18226
rect 7208 17054 7328 17082
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 7024 15706 7052 15846
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7116 15502 7144 15982
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7012 15360 7064 15366
rect 6918 15328 6974 15337
rect 7012 15302 7064 15308
rect 6918 15263 6974 15272
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6932 14550 6960 14758
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 7024 13870 7052 15302
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6552 12378 6604 12384
rect 6656 12406 6776 12434
rect 6458 12200 6514 12209
rect 6458 12135 6514 12144
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10674 6500 10950
rect 6564 10810 6592 12378
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5166 6040 5646
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6012 4554 6040 5102
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4729 6132 5034
rect 6090 4720 6146 4729
rect 6090 4655 6146 4664
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6196 4486 6224 7278
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6288 5817 6316 5850
rect 6274 5808 6330 5817
rect 6274 5743 6330 5752
rect 6380 4554 6408 8026
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 5920 4214 5948 4422
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 5276 3590 5580 3618
rect 5276 3398 5304 3590
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5264 2984 5316 2990
rect 5262 2952 5264 2961
rect 5316 2952 5318 2961
rect 5262 2887 5318 2896
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2650 5672 2790
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5828 2310 5856 3130
rect 5906 2408 5962 2417
rect 5906 2343 5908 2352
rect 5960 2343 5962 2352
rect 5908 2314 5960 2320
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6472 800 6500 8910
rect 6656 7478 6684 12406
rect 6840 11830 6868 12854
rect 6932 12170 6960 13330
rect 7024 13258 7052 13670
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 7024 11762 7052 13194
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6920 11348 6972 11354
rect 6972 11308 7052 11336
rect 6920 11290 6972 11296
rect 6840 11234 6868 11290
rect 6840 11206 6960 11234
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6734 10840 6790 10849
rect 6734 10775 6736 10784
rect 6788 10775 6790 10784
rect 6736 10746 6788 10752
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 10441 6776 10542
rect 6734 10432 6790 10441
rect 6734 10367 6790 10376
rect 6840 10062 6868 11086
rect 6932 10810 6960 11206
rect 7024 11082 7052 11308
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6932 10470 6960 10610
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6840 9586 6868 9998
rect 6918 9752 6974 9761
rect 6918 9687 6974 9696
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6932 9450 6960 9687
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6826 8936 6882 8945
rect 6748 7954 6776 8910
rect 6826 8871 6882 8880
rect 6840 8430 6868 8871
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6564 6254 6592 7346
rect 6748 6866 6776 7890
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6552 6248 6604 6254
rect 6840 6225 6868 8366
rect 6932 7478 6960 9386
rect 7024 7750 7052 11018
rect 7116 7970 7144 14758
rect 7208 12434 7236 17054
rect 7392 16289 7420 18702
rect 7484 18686 7604 18714
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7484 17814 7512 18686
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 7562 17776 7618 17785
rect 7378 16280 7434 16289
rect 7378 16215 7380 16224
rect 7432 16215 7434 16224
rect 7380 16186 7432 16192
rect 7392 16155 7420 16186
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7300 15094 7328 15574
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7300 14414 7328 15030
rect 7392 14958 7420 15370
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7288 14000 7340 14006
rect 7286 13968 7288 13977
rect 7340 13968 7342 13977
rect 7286 13903 7342 13912
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7300 13394 7328 13466
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7392 12918 7420 14894
rect 7484 13682 7512 17750
rect 7562 17711 7564 17720
rect 7616 17711 7618 17720
rect 7564 17682 7616 17688
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16658 7604 17070
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7576 15638 7604 16050
rect 7564 15632 7616 15638
rect 7564 15574 7616 15580
rect 7668 14498 7696 18294
rect 7576 14470 7696 14498
rect 7576 13818 7604 14470
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7668 14006 7696 14282
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7576 13790 7696 13818
rect 7484 13654 7604 13682
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7380 12436 7432 12442
rect 7208 12406 7328 12434
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 11082 7236 11630
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 9994 7236 10406
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7116 7942 7236 7970
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 6730 7052 7278
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7116 6866 7144 7142
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6552 6190 6604 6196
rect 6826 6216 6882 6225
rect 6564 5030 6592 6190
rect 6826 6151 6882 6160
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5642 6684 6054
rect 6734 5944 6790 5953
rect 6734 5879 6790 5888
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6748 5574 6776 5879
rect 6826 5672 6882 5681
rect 6826 5607 6882 5616
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6564 3602 6592 4014
rect 6840 3738 6868 5607
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6564 3058 6592 3538
rect 6828 3460 6880 3466
rect 6932 3448 6960 6394
rect 7024 6390 7052 6666
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7024 5778 7052 6326
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7024 5302 7052 5714
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 7024 4690 7052 5238
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7116 4214 7144 6190
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7012 3460 7064 3466
rect 6932 3420 7012 3448
rect 6828 3402 6880 3408
rect 7012 3402 7064 3408
rect 6840 3346 6868 3402
rect 6840 3318 6960 3346
rect 6828 3120 6880 3126
rect 6826 3088 6828 3097
rect 6880 3088 6882 3097
rect 6552 3052 6604 3058
rect 6826 3023 6882 3032
rect 6552 2994 6604 3000
rect 6564 2514 6592 2994
rect 6932 2990 6960 3318
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 7116 800 7144 3674
rect 7208 3466 7236 7942
rect 7300 6662 7328 12406
rect 7380 12378 7432 12384
rect 7392 11762 7420 12378
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 10674 7420 11698
rect 7484 10849 7512 12854
rect 7576 11354 7604 13654
rect 7668 11642 7696 13790
rect 7760 12434 7788 18702
rect 7944 18290 7972 19110
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 8036 18170 8064 19450
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7944 18142 8064 18170
rect 7944 16794 7972 18142
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7838 15464 7894 15473
rect 7838 15399 7840 15408
rect 7892 15399 7894 15408
rect 7840 15370 7892 15376
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7852 13938 7880 14962
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7944 13433 7972 16730
rect 8036 15094 8064 17206
rect 8128 16658 8156 19178
rect 8220 18057 8248 30534
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8312 19854 8340 21082
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8312 18766 8340 19246
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8404 18612 8432 21626
rect 8496 21146 8524 24210
rect 9048 24206 9076 24754
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8588 23118 8616 23462
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8588 19334 8616 20810
rect 8680 20534 8708 21286
rect 8864 20602 8892 21558
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 8956 20942 8984 21082
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8588 19306 8892 19334
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8312 18584 8432 18612
rect 8206 18048 8262 18057
rect 8206 17983 8262 17992
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8208 16584 8260 16590
rect 8206 16552 8208 16561
rect 8260 16552 8262 16561
rect 8312 16538 8340 18584
rect 8392 17536 8444 17542
rect 8496 17513 8524 18906
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8392 17478 8444 17484
rect 8482 17504 8538 17513
rect 8404 16810 8432 17478
rect 8482 17439 8538 17448
rect 8482 17368 8538 17377
rect 8588 17338 8616 17750
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8482 17303 8538 17312
rect 8576 17332 8628 17338
rect 8496 17202 8524 17303
rect 8576 17274 8628 17280
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8404 16782 8524 16810
rect 8496 16726 8524 16782
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8312 16510 8432 16538
rect 8206 16487 8262 16496
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8220 15337 8248 16050
rect 8206 15328 8262 15337
rect 8206 15263 8262 15272
rect 8312 15094 8340 16390
rect 8404 16250 8432 16510
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 16250 8524 16390
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8588 16130 8616 16594
rect 8404 16102 8616 16130
rect 8024 15088 8076 15094
rect 8300 15088 8352 15094
rect 8076 15048 8156 15076
rect 8024 15030 8076 15036
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7930 13424 7986 13433
rect 7930 13359 7986 13368
rect 7760 12406 7972 12434
rect 7838 12200 7894 12209
rect 7838 12135 7894 12144
rect 7852 12102 7880 12135
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7668 11614 7788 11642
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7562 11248 7618 11257
rect 7562 11183 7618 11192
rect 7470 10840 7526 10849
rect 7470 10775 7526 10784
rect 7576 10690 7604 11183
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7484 10662 7604 10690
rect 7380 9988 7432 9994
rect 7484 9976 7512 10662
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 9994 7604 10406
rect 7432 9948 7512 9976
rect 7380 9930 7432 9936
rect 7288 6656 7340 6662
rect 7380 6656 7432 6662
rect 7288 6598 7340 6604
rect 7378 6624 7380 6633
rect 7432 6624 7434 6633
rect 7378 6559 7434 6568
rect 7286 5808 7342 5817
rect 7286 5743 7288 5752
rect 7340 5743 7342 5752
rect 7288 5714 7340 5720
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7484 2961 7512 9948
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7668 6730 7696 11494
rect 7760 8838 7788 11614
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7852 5574 7880 12038
rect 7944 9926 7972 12406
rect 8036 11529 8064 14214
rect 8128 13190 8156 15048
rect 8300 15030 8352 15036
rect 8404 14890 8432 16102
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8588 15745 8616 15846
rect 8574 15736 8630 15745
rect 8574 15671 8630 15680
rect 8482 15600 8538 15609
rect 8482 15535 8538 15544
rect 8496 15366 8524 15535
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8482 14920 8538 14929
rect 8392 14884 8444 14890
rect 8482 14855 8538 14864
rect 8392 14826 8444 14832
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8298 14784 8354 14793
rect 8220 14521 8248 14758
rect 8298 14719 8354 14728
rect 8206 14512 8262 14521
rect 8206 14447 8262 14456
rect 8312 14074 8340 14719
rect 8390 14648 8446 14657
rect 8496 14618 8524 14855
rect 8390 14583 8446 14592
rect 8484 14612 8536 14618
rect 8404 14550 8432 14583
rect 8484 14554 8536 14560
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 13258 8340 13874
rect 8404 13841 8432 14350
rect 8588 14346 8616 15438
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8484 14272 8536 14278
rect 8482 14240 8484 14249
rect 8536 14240 8538 14249
rect 8482 14175 8538 14184
rect 8390 13832 8446 13841
rect 8390 13767 8446 13776
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8128 12238 8156 13126
rect 8404 12481 8432 13126
rect 8390 12472 8446 12481
rect 8390 12407 8446 12416
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8496 12306 8524 12378
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8114 11928 8170 11937
rect 8114 11863 8170 11872
rect 8128 11830 8156 11863
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8022 11520 8078 11529
rect 8022 11455 8078 11464
rect 8312 11354 8340 11630
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8036 10282 8064 10746
rect 8208 10464 8260 10470
rect 8206 10432 8208 10441
rect 8300 10464 8352 10470
rect 8260 10432 8262 10441
rect 8404 10452 8432 12174
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8352 10424 8432 10452
rect 8300 10406 8352 10412
rect 8206 10367 8262 10376
rect 8206 10296 8262 10305
rect 8036 10254 8156 10282
rect 8022 10160 8078 10169
rect 8022 10095 8078 10104
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7944 4826 7972 9862
rect 8036 9382 8064 10095
rect 8128 9926 8156 10254
rect 8206 10231 8262 10240
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 8838 8064 9046
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8128 3126 8156 6802
rect 8220 6322 8248 10231
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8312 7478 8340 10066
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8298 6216 8354 6225
rect 8298 6151 8300 6160
rect 8352 6151 8354 6160
rect 8300 6122 8352 6128
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5846 8248 6054
rect 8404 5930 8432 8978
rect 8312 5902 8432 5930
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8206 5672 8262 5681
rect 8206 5607 8262 5616
rect 8220 4078 8248 5607
rect 8312 4826 8340 5902
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8404 5234 8432 5714
rect 8496 5642 8524 12038
rect 8588 8974 8616 13670
rect 8680 11014 8708 17614
rect 8772 13530 8800 18702
rect 8864 14414 8892 19306
rect 8956 15910 8984 20538
rect 9048 19689 9076 24142
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9416 23798 9444 24006
rect 9404 23792 9456 23798
rect 9404 23734 9456 23740
rect 9508 23730 9536 24074
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9404 23588 9456 23594
rect 9404 23530 9456 23536
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22642 9352 23054
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 21554 9168 22442
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9034 19680 9090 19689
rect 9034 19615 9090 19624
rect 9036 19508 9088 19514
rect 9140 19496 9168 20266
rect 9220 19848 9272 19854
rect 9218 19816 9220 19825
rect 9272 19816 9274 19825
rect 9218 19751 9274 19760
rect 9088 19468 9168 19496
rect 9036 19450 9088 19456
rect 9126 19374 9182 19383
rect 9048 19318 9126 19334
rect 9048 19309 9182 19318
rect 9048 19306 9168 19309
rect 9048 18873 9076 19306
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9034 18864 9090 18873
rect 9034 18799 9090 18808
rect 9140 18714 9168 19110
rect 9232 18834 9260 19246
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9140 18686 9260 18714
rect 9232 18630 9260 18686
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9034 17504 9090 17513
rect 9034 17439 9090 17448
rect 9048 17202 9076 17439
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9140 16454 9168 18566
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8758 13424 8814 13433
rect 8758 13359 8814 13368
rect 8772 11370 8800 13359
rect 8864 12442 8892 13806
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8772 11342 8892 11370
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8666 10840 8722 10849
rect 8666 10775 8722 10784
rect 8680 9518 8708 10775
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8772 8906 8800 11222
rect 8864 9450 8892 11342
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8574 8528 8630 8537
rect 8574 8463 8630 8472
rect 8588 8362 8616 8463
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8588 6662 8616 8298
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8666 6896 8722 6905
rect 8666 6831 8722 6840
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8588 5545 8616 5850
rect 8574 5536 8630 5545
rect 8574 5471 8630 5480
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8298 4040 8354 4049
rect 8298 3975 8354 3984
rect 8312 3942 8340 3975
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 7470 2952 7526 2961
rect 7470 2887 7526 2896
rect 8404 800 8432 4558
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8496 3398 8524 3606
rect 8588 3398 8616 5471
rect 8680 5302 8708 6831
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8772 4321 8800 8230
rect 8850 5944 8906 5953
rect 8850 5879 8852 5888
rect 8904 5879 8906 5888
rect 8852 5850 8904 5856
rect 8758 4312 8814 4321
rect 8758 4247 8814 4256
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8574 3224 8630 3233
rect 8574 3159 8630 3168
rect 8588 3126 8616 3159
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8956 2378 8984 14962
rect 9048 13734 9076 16118
rect 9140 16046 9168 16118
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 9036 13728 9088 13734
rect 9140 13705 9168 15574
rect 9232 15337 9260 18226
rect 9218 15328 9274 15337
rect 9218 15263 9274 15272
rect 9218 15056 9274 15065
rect 9218 14991 9274 15000
rect 9232 14657 9260 14991
rect 9218 14648 9274 14657
rect 9218 14583 9274 14592
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9036 13670 9088 13676
rect 9126 13696 9182 13705
rect 9126 13631 9182 13640
rect 9034 13560 9090 13569
rect 9034 13495 9090 13504
rect 9128 13524 9180 13530
rect 9048 11830 9076 13495
rect 9128 13466 9180 13472
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 9034 11656 9090 11665
rect 9034 11591 9090 11600
rect 9048 11558 9076 11591
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11257 9076 11494
rect 9034 11248 9090 11257
rect 9034 11183 9090 11192
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 6458 9076 10950
rect 9140 10538 9168 13466
rect 9232 13190 9260 14418
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9232 12782 9260 12922
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11218 9260 11562
rect 9324 11354 9352 22578
rect 9416 22574 9444 23530
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9508 19145 9536 23666
rect 9600 19174 9628 24618
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 10152 24206 10180 24550
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10244 24018 10272 24550
rect 10152 23990 10272 24018
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9678 21040 9734 21049
rect 9678 20975 9734 20984
rect 9692 20942 9720 20975
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9680 20800 9732 20806
rect 9678 20768 9680 20777
rect 9732 20768 9734 20777
rect 9678 20703 9734 20712
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9588 19168 9640 19174
rect 9494 19136 9550 19145
rect 9588 19110 9640 19116
rect 9494 19071 9550 19080
rect 9692 18986 9720 20470
rect 9600 18958 9720 18986
rect 9494 18864 9550 18873
rect 9494 18799 9550 18808
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9416 17270 9444 17818
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9402 16824 9458 16833
rect 9402 16759 9458 16768
rect 9416 16658 9444 16759
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16425 9444 16458
rect 9402 16416 9458 16425
rect 9402 16351 9458 16360
rect 9508 15881 9536 18799
rect 9600 16402 9628 18958
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 16708 9720 18022
rect 9784 17610 9812 22374
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9876 20369 9904 21354
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9876 16810 9904 18090
rect 9968 17746 9996 22034
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10060 20534 10088 20742
rect 10048 20528 10100 20534
rect 10048 20470 10100 20476
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10060 17218 10088 19994
rect 10152 18834 10180 23990
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10244 22778 10272 23122
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10336 21554 10364 23190
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10232 20936 10284 20942
rect 10428 20890 10456 31826
rect 11072 30734 11100 37130
rect 14844 37126 14872 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 14924 37256 14976 37262
rect 14922 37224 14924 37233
rect 14976 37224 14978 37233
rect 14922 37159 14978 37168
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 14832 37120 14884 37126
rect 14832 37062 14884 37068
rect 11716 31958 11744 37062
rect 11796 36916 11848 36922
rect 11796 36858 11848 36864
rect 11808 36786 11836 36858
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10968 30660 11020 30666
rect 10968 30602 11020 30608
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10520 23798 10548 30194
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10704 24614 10732 29446
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10980 24274 11008 30602
rect 11164 30122 11192 30738
rect 11152 30116 11204 30122
rect 11152 30058 11204 30064
rect 11808 28558 11836 36722
rect 12360 32502 12388 37062
rect 12544 35834 12572 37062
rect 12532 35828 12584 35834
rect 12532 35770 12584 35776
rect 13912 35692 13964 35698
rect 13912 35634 13964 35640
rect 13924 32570 13952 35634
rect 13912 32564 13964 32570
rect 13912 32506 13964 32512
rect 12348 32496 12400 32502
rect 12348 32438 12400 32444
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12452 26450 12480 26930
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 11520 26308 11572 26314
rect 11520 26250 11572 26256
rect 11244 25220 11296 25226
rect 11244 25162 11296 25168
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10888 24177 10916 24210
rect 11256 24206 11284 25162
rect 11244 24200 11296 24206
rect 10874 24168 10930 24177
rect 11244 24142 11296 24148
rect 10874 24103 10930 24112
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10508 23792 10560 23798
rect 10508 23734 10560 23740
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10704 22778 10732 23054
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10284 20884 10456 20890
rect 10232 20878 10456 20884
rect 10244 20862 10456 20878
rect 10520 20874 10548 22374
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9968 17190 10088 17218
rect 9968 16998 9996 17190
rect 10140 17128 10192 17134
rect 10046 17096 10102 17105
rect 10140 17070 10192 17076
rect 10046 17031 10048 17040
rect 10100 17031 10102 17040
rect 10048 17002 10100 17008
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9876 16782 10088 16810
rect 9692 16680 9996 16708
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9876 16425 9904 16458
rect 9862 16416 9918 16425
rect 9600 16374 9720 16402
rect 9692 16232 9720 16374
rect 9862 16351 9918 16360
rect 9600 16204 9720 16232
rect 9494 15872 9550 15881
rect 9494 15807 9550 15816
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9508 15162 9536 15574
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 13682 9444 14758
rect 9508 13841 9536 14962
rect 9494 13832 9550 13841
rect 9494 13767 9550 13776
rect 9416 13654 9536 13682
rect 9402 13560 9458 13569
rect 9402 13495 9458 13504
rect 9416 12986 9444 13495
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9416 12306 9444 12718
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9416 11218 9444 12242
rect 9508 11558 9536 13654
rect 9600 13569 9628 16204
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9586 13560 9642 13569
rect 9586 13495 9642 13504
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9600 12986 9628 13194
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9600 11150 9628 12922
rect 9692 12345 9720 15982
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15434 9812 15914
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9770 15192 9826 15201
rect 9770 15127 9826 15136
rect 9784 13394 9812 15127
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9772 13252 9824 13258
rect 9876 13240 9904 15642
rect 9968 15434 9996 16680
rect 10060 16182 10088 16782
rect 10048 16176 10100 16182
rect 10048 16118 10100 16124
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 14226 10088 15302
rect 10152 14657 10180 17070
rect 10138 14648 10194 14657
rect 10138 14583 10194 14592
rect 10244 14482 10272 20334
rect 10428 19786 10456 20862
rect 10508 20868 10560 20874
rect 10508 20810 10560 20816
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18086 10364 18906
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10336 16726 10364 17682
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10322 15736 10378 15745
rect 10322 15671 10378 15680
rect 10336 15366 10364 15671
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10428 14804 10456 17750
rect 10520 17270 10548 19314
rect 10508 17264 10560 17270
rect 10508 17206 10560 17212
rect 10612 17082 10640 21830
rect 10704 19446 10732 22714
rect 10796 21962 10824 22918
rect 10784 21956 10836 21962
rect 10784 21898 10836 21904
rect 10888 21570 10916 23802
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 11072 22778 11100 23598
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10966 21720 11022 21729
rect 11072 21690 11100 22714
rect 10966 21655 10968 21664
rect 11020 21655 11022 21664
rect 11060 21684 11112 21690
rect 10968 21626 11020 21632
rect 11060 21626 11112 21632
rect 10888 21542 11100 21570
rect 11072 21418 11100 21542
rect 11164 21486 11192 24006
rect 11348 22710 11376 24006
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11336 22704 11388 22710
rect 11336 22646 11388 22652
rect 11440 22506 11468 22714
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 11428 22500 11480 22506
rect 11428 22442 11480 22448
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10704 18306 10732 19382
rect 10796 19378 10824 21286
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10888 20777 10916 20810
rect 10874 20768 10930 20777
rect 10874 20703 10930 20712
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 19446 10916 19654
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10980 18737 11008 19790
rect 11072 18834 11100 21014
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10966 18728 11022 18737
rect 10784 18692 10836 18698
rect 10966 18663 11022 18672
rect 10784 18634 10836 18640
rect 10796 18426 10824 18634
rect 10966 18456 11022 18465
rect 10784 18420 10836 18426
rect 10966 18391 11022 18400
rect 11060 18420 11112 18426
rect 10784 18362 10836 18368
rect 10704 18278 10824 18306
rect 10980 18290 11008 18391
rect 11060 18362 11112 18368
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10704 17542 10732 17750
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10704 17105 10732 17206
rect 10336 14776 10456 14804
rect 10520 17054 10640 17082
rect 10690 17096 10746 17105
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 14385 10272 14418
rect 10230 14376 10286 14385
rect 10230 14311 10286 14320
rect 9968 14198 10088 14226
rect 9968 13938 9996 14198
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10060 13394 10088 14039
rect 10140 14000 10192 14006
rect 10138 13968 10140 13977
rect 10192 13968 10194 13977
rect 10138 13903 10194 13912
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9824 13212 9904 13240
rect 9772 13194 9824 13200
rect 10060 13025 10088 13330
rect 10046 13016 10102 13025
rect 10046 12951 10102 12960
rect 9770 12880 9826 12889
rect 9770 12815 9826 12824
rect 9678 12336 9734 12345
rect 9784 12306 9812 12815
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9678 12271 9734 12280
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 12170 9904 12242
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9508 10985 9536 11086
rect 9494 10976 9550 10985
rect 9494 10911 9550 10920
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9416 10470 9444 10610
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9218 9888 9274 9897
rect 9218 9823 9274 9832
rect 9126 9752 9182 9761
rect 9232 9722 9260 9823
rect 9126 9687 9182 9696
rect 9220 9716 9272 9722
rect 9140 8294 9168 9687
rect 9220 9658 9272 9664
rect 9310 9616 9366 9625
rect 9310 9551 9366 9560
rect 9324 9382 9352 9551
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9402 9344 9458 9353
rect 9402 9279 9458 9288
rect 9416 9178 9444 9279
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9508 9058 9536 10911
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9232 9030 9536 9058
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9232 6798 9260 9030
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7002 9352 7686
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5778 9168 6258
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9232 4622 9260 6734
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9232 4282 9260 4422
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9416 3738 9444 8434
rect 9494 8256 9550 8265
rect 9494 8191 9550 8200
rect 9508 5642 9536 8191
rect 9600 6730 9628 10406
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9722 9720 9998
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9692 9081 9720 9658
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9784 9353 9812 9454
rect 9770 9344 9826 9353
rect 9770 9279 9826 9288
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9680 8832 9732 8838
rect 9876 8820 9904 12106
rect 10060 10266 10088 12718
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9732 8792 9904 8820
rect 9680 8774 9732 8780
rect 9678 8664 9734 8673
rect 9678 8599 9680 8608
rect 9732 8599 9734 8608
rect 9680 8570 9732 8576
rect 9692 6866 9720 8570
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 7342 9812 7482
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9126 3496 9182 3505
rect 9126 3431 9182 3440
rect 9404 3460 9456 3466
rect 9140 3398 9168 3431
rect 9404 3402 9456 3408
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9416 3074 9444 3402
rect 9324 3058 9444 3074
rect 9312 3052 9444 3058
rect 9364 3046 9444 3052
rect 9312 2994 9364 3000
rect 9508 2854 9536 4694
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4214 9812 4626
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9784 3602 9812 4150
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9588 3120 9640 3126
rect 9784 3074 9812 3538
rect 9640 3068 9812 3074
rect 9588 3062 9812 3068
rect 9600 3046 9812 3062
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9784 2514 9812 3046
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9876 2394 9904 7210
rect 9968 6730 9996 9930
rect 10046 9072 10102 9081
rect 10046 9007 10102 9016
rect 10060 8906 10088 9007
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10152 8090 10180 13670
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10244 12170 10272 12582
rect 10336 12306 10364 14776
rect 10520 14634 10548 17054
rect 10690 17031 10746 17040
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10428 14606 10548 14634
rect 10428 12782 10456 14606
rect 10506 14376 10562 14385
rect 10506 14311 10562 14320
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10232 12164 10284 12170
rect 10232 12106 10284 12112
rect 10428 11937 10456 12378
rect 10414 11928 10470 11937
rect 10414 11863 10470 11872
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 10169 10272 10610
rect 10230 10160 10286 10169
rect 10230 10095 10286 10104
rect 10232 9648 10284 9654
rect 10230 9616 10232 9625
rect 10284 9616 10286 9625
rect 10230 9551 10286 9560
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10244 7478 10272 8434
rect 10232 7472 10284 7478
rect 10232 7414 10284 7420
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 10060 4690 10088 7278
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10046 4584 10102 4593
rect 10046 4519 10048 4528
rect 10100 4519 10102 4528
rect 10048 4490 10100 4496
rect 10060 3942 10088 4490
rect 10152 4162 10180 7346
rect 10336 5302 10364 11018
rect 10520 10674 10548 14311
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8945 10456 8978
rect 10414 8936 10470 8945
rect 10414 8871 10470 8880
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10520 7546 10548 8570
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10520 6866 10548 7482
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10152 4134 10272 4162
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10152 3466 10180 4014
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 9956 3120 10008 3126
rect 10244 3108 10272 4134
rect 10008 3080 10272 3108
rect 9956 3062 10008 3068
rect 10428 2774 10456 5714
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 9692 2366 9904 2394
rect 10336 2746 10456 2774
rect 9956 2372 10008 2378
rect 9692 800 9720 2366
rect 9956 2314 10008 2320
rect 9968 1834 9996 2314
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 10336 800 10364 2746
rect 10612 2310 10640 16526
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10704 15638 10732 16050
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10704 14385 10732 15574
rect 10690 14376 10746 14385
rect 10690 14311 10746 14320
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10796 14226 10824 18278
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10888 17882 10916 18226
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 15638 10916 16390
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10874 15056 10930 15065
rect 10874 14991 10930 15000
rect 10888 14346 10916 14991
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10704 9330 10732 14214
rect 10796 14198 10916 14226
rect 10888 11082 10916 14198
rect 10980 12617 11008 17546
rect 11072 16833 11100 18362
rect 11058 16824 11114 16833
rect 11058 16759 11114 16768
rect 11072 16658 11100 16759
rect 11164 16697 11192 21082
rect 11256 20534 11284 22442
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11256 16708 11284 17070
rect 11348 16810 11376 18566
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11440 17270 11468 18022
rect 11532 17762 11560 26250
rect 12164 24336 12216 24342
rect 12164 24278 12216 24284
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21690 11744 21898
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11624 19514 11652 19722
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11624 19145 11652 19246
rect 11610 19136 11666 19145
rect 11610 19071 11666 19080
rect 11716 18426 11744 19450
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11716 18057 11744 18226
rect 11702 18048 11758 18057
rect 11702 17983 11758 17992
rect 11808 17882 11836 19926
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11532 17734 11744 17762
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11348 16782 11560 16810
rect 11336 16720 11388 16726
rect 11150 16688 11206 16697
rect 11060 16652 11112 16658
rect 11256 16680 11336 16708
rect 11336 16662 11388 16668
rect 11150 16623 11206 16632
rect 11060 16594 11112 16600
rect 11244 16584 11296 16590
rect 11150 16552 11206 16561
rect 11244 16526 11296 16532
rect 11150 16487 11206 16496
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11072 15706 11100 15982
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11164 14278 11192 16487
rect 11256 15026 11284 16526
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 13326 11100 13806
rect 11256 13546 11284 14282
rect 11348 13734 11376 16662
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11440 15337 11468 15370
rect 11426 15328 11482 15337
rect 11426 15263 11482 15272
rect 11426 14512 11482 14521
rect 11426 14447 11482 14456
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11256 13518 11376 13546
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12918 11100 13262
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11072 12646 11100 12854
rect 11060 12640 11112 12646
rect 10966 12608 11022 12617
rect 11060 12582 11112 12588
rect 10966 12543 11022 12552
rect 11060 12096 11112 12102
rect 11058 12064 11060 12073
rect 11112 12064 11114 12073
rect 11058 11999 11114 12008
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10980 10674 11008 10950
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10704 9302 10824 9330
rect 10690 7984 10746 7993
rect 10690 7919 10746 7928
rect 10704 6254 10732 7919
rect 10796 6322 10824 9302
rect 10888 7478 10916 10406
rect 11072 9586 11100 11630
rect 11164 10180 11192 13194
rect 11256 12850 11284 13398
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 11830 11284 12582
rect 11348 12442 11376 13518
rect 11440 12617 11468 14447
rect 11532 13258 11560 16782
rect 11624 15502 11652 17614
rect 11716 16454 11744 17734
rect 11794 17504 11850 17513
rect 11794 17439 11850 17448
rect 11808 16658 11836 17439
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11624 14906 11652 15438
rect 11808 14958 11836 16594
rect 11900 15570 11928 22578
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 17785 12020 20334
rect 11978 17776 12034 17785
rect 11978 17711 12034 17720
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11992 17202 12020 17614
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11796 14952 11848 14958
rect 11624 14878 11744 14906
rect 11796 14894 11848 14900
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12753 11560 12786
rect 11518 12744 11574 12753
rect 11518 12679 11574 12688
rect 11426 12608 11482 12617
rect 11426 12543 11482 12552
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11334 12200 11390 12209
rect 11334 12135 11390 12144
rect 11348 12102 11376 12135
rect 11336 12096 11388 12102
rect 11388 12044 11468 12050
rect 11336 12038 11468 12044
rect 11348 12022 11468 12038
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11256 11218 11284 11766
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11348 11082 11376 11834
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11244 10192 11296 10198
rect 11164 10152 11244 10180
rect 11244 10134 11296 10140
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 10966 9480 11022 9489
rect 11348 9466 11376 9658
rect 10966 9415 11022 9424
rect 11072 9438 11376 9466
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10690 3768 10746 3777
rect 10690 3703 10746 3712
rect 10704 2990 10732 3703
rect 10796 3602 10824 5850
rect 10980 5778 11008 9415
rect 11072 5846 11100 9438
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11164 9178 11192 9318
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11244 8288 11296 8294
rect 11150 8256 11206 8265
rect 11244 8230 11296 8236
rect 11150 8191 11206 8200
rect 11164 7410 11192 8191
rect 11256 7818 11284 8230
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 11164 6118 11192 6831
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11164 5370 11192 6054
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10968 4208 11020 4214
rect 10966 4176 10968 4185
rect 11020 4176 11022 4185
rect 10966 4111 11022 4120
rect 11348 4078 11376 9318
rect 11440 7206 11468 12022
rect 11532 7732 11560 12679
rect 11624 12306 11652 14486
rect 11716 13161 11744 14878
rect 11992 14260 12020 17138
rect 12084 16182 12112 23190
rect 12176 22574 12204 24278
rect 12346 24168 12402 24177
rect 12346 24103 12348 24112
rect 12400 24103 12402 24112
rect 12348 24074 12400 24080
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12268 21894 12296 22034
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12348 21888 12400 21894
rect 12348 21830 12400 21836
rect 12360 21570 12388 21830
rect 12268 21542 12388 21570
rect 12268 20806 12296 21542
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12360 21010 12388 21422
rect 12348 21004 12400 21010
rect 12348 20946 12400 20952
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12254 20088 12310 20097
rect 12254 20023 12310 20032
rect 12348 20052 12400 20058
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12176 18290 12204 18702
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12084 14482 12112 16118
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15434 12204 15846
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11900 14232 12020 14260
rect 11702 13152 11758 13161
rect 11702 13087 11758 13096
rect 11900 12986 11928 14232
rect 12268 14226 12296 20023
rect 12348 19994 12400 20000
rect 12360 19446 12388 19994
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12360 18834 12388 19246
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12348 17672 12400 17678
rect 12346 17640 12348 17649
rect 12400 17640 12402 17649
rect 12346 17575 12402 17584
rect 12452 17241 12480 26386
rect 12820 25906 12848 26726
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 12808 24336 12860 24342
rect 12808 24278 12860 24284
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12728 23118 12756 23598
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12544 22030 12572 22986
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12728 22234 12756 22918
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12636 21010 12664 22034
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12728 20602 12756 21422
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12544 18290 12572 19858
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 17377 12572 17478
rect 12530 17368 12586 17377
rect 12530 17303 12586 17312
rect 12438 17232 12494 17241
rect 12438 17167 12494 17176
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12360 14346 12388 15574
rect 12452 15094 12480 16050
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12176 14198 12296 14226
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11716 12714 11744 12922
rect 12084 12918 12112 14010
rect 12176 13938 12204 14198
rect 12530 14104 12586 14113
rect 12530 14039 12586 14048
rect 12544 14006 12572 14039
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11716 11694 11744 12650
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12254 12608 12310 12617
rect 12084 12424 12112 12582
rect 12254 12543 12310 12552
rect 11992 12396 12112 12424
rect 12162 12472 12218 12481
rect 12162 12407 12218 12416
rect 11794 12336 11850 12345
rect 11794 12271 11850 12280
rect 11808 12170 11836 12271
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11624 10606 11652 11154
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11702 10432 11758 10441
rect 11624 8566 11652 10406
rect 11702 10367 11758 10376
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11532 7704 11652 7732
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11426 7032 11482 7041
rect 11426 6967 11482 6976
rect 11440 6662 11468 6967
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11336 4072 11388 4078
rect 11058 4040 11114 4049
rect 11336 4014 11388 4020
rect 11058 3975 11060 3984
rect 11112 3975 11114 3984
rect 11060 3946 11112 3952
rect 11060 3664 11112 3670
rect 11058 3632 11060 3641
rect 11112 3632 11114 3641
rect 10784 3596 10836 3602
rect 11058 3567 11114 3576
rect 10784 3538 10836 3544
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10888 2990 10916 3334
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10980 1290 11008 3062
rect 11532 1850 11560 5170
rect 11624 3058 11652 7704
rect 11716 4826 11744 10367
rect 11808 5574 11836 12106
rect 11900 11830 11928 12174
rect 11992 12102 12020 12396
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 11900 11286 11928 11562
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11978 9480 12034 9489
rect 11978 9415 12034 9424
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11900 8945 11928 8978
rect 11886 8936 11942 8945
rect 11886 8871 11942 8880
rect 11900 8566 11928 8871
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11900 7478 11928 7754
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11992 6866 12020 9415
rect 12084 7750 12112 11562
rect 12176 11082 12204 12407
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12268 8906 12296 12543
rect 12360 12170 12388 13126
rect 12438 13016 12494 13025
rect 12438 12951 12440 12960
rect 12492 12951 12494 12960
rect 12440 12922 12492 12928
rect 12544 12220 12572 13194
rect 12636 12782 12664 20402
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 16522 12756 18566
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12820 15910 12848 24278
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13004 20602 13032 21966
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12912 19514 12940 19926
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12912 18154 12940 19450
rect 13004 18834 13032 19994
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 12900 18148 12952 18154
rect 12900 18090 12952 18096
rect 13096 17320 13124 25162
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 22098 13216 22918
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13280 21622 13308 22170
rect 13268 21616 13320 21622
rect 13268 21558 13320 21564
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13188 18601 13216 20402
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13280 19378 13308 20198
rect 13372 19922 13400 30534
rect 14108 29170 14136 37062
rect 15568 36848 15620 36854
rect 15568 36790 15620 36796
rect 15476 36576 15528 36582
rect 15476 36518 15528 36524
rect 15016 32428 15068 32434
rect 15016 32370 15068 32376
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14096 28416 14148 28422
rect 14096 28358 14148 28364
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13740 26382 13768 26726
rect 14004 26512 14056 26518
rect 14004 26454 14056 26460
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 13832 23730 13860 24686
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13924 23662 13952 25094
rect 14016 23730 14044 26454
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13268 19236 13320 19242
rect 13372 19224 13400 19654
rect 13320 19196 13400 19224
rect 13268 19178 13320 19184
rect 13464 18873 13492 20402
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19786 13584 20198
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13450 18864 13506 18873
rect 13450 18799 13506 18808
rect 13174 18592 13230 18601
rect 13174 18527 13230 18536
rect 12912 17292 13124 17320
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12728 14618 12756 14758
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12714 14376 12770 14385
rect 12714 14311 12770 14320
rect 12728 13530 12756 14311
rect 12820 13530 12848 14758
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 13190 12848 13466
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12452 12192 12572 12220
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12360 9722 12388 11766
rect 12452 11354 12480 12192
rect 12636 11830 12664 12718
rect 12912 11914 12940 17292
rect 13188 17048 13216 18527
rect 13450 18456 13506 18465
rect 13450 18391 13506 18400
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13280 17610 13308 17750
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13096 17020 13216 17048
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 13004 14929 13032 15030
rect 12990 14920 13046 14929
rect 12990 14855 12992 14864
rect 13044 14855 13046 14864
rect 12992 14826 13044 14832
rect 13004 14795 13032 14826
rect 13096 14362 13124 17020
rect 13280 16946 13308 17138
rect 13188 16918 13308 16946
rect 13188 16046 13216 16918
rect 13266 16824 13322 16833
rect 13266 16759 13268 16768
rect 13320 16759 13322 16768
rect 13268 16730 13320 16736
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13188 14482 13216 15982
rect 13280 15570 13308 16390
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13266 15328 13322 15337
rect 13266 15263 13322 15272
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13096 14334 13216 14362
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12728 11886 12940 11914
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12728 10690 12756 11886
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12820 10810 12848 11766
rect 13004 11286 13032 13738
rect 13096 11694 13124 14214
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 13188 11218 13216 14334
rect 13280 12889 13308 15263
rect 13372 15094 13400 18022
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13372 13161 13400 14894
rect 13464 14278 13492 18391
rect 13556 18222 13584 19110
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13648 17252 13676 22578
rect 13740 22574 13768 23462
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13728 22432 13780 22438
rect 13728 22374 13780 22380
rect 13740 21010 13768 22374
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 13832 21486 13860 21558
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13910 21448 13966 21457
rect 13910 21383 13966 21392
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13726 20904 13782 20913
rect 13726 20839 13782 20848
rect 13740 19922 13768 20839
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13740 19417 13768 19858
rect 13726 19408 13782 19417
rect 13726 19343 13782 19352
rect 13924 19334 13952 21383
rect 13924 19306 14044 19334
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13556 17224 13676 17252
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13358 13152 13414 13161
rect 13358 13087 13414 13096
rect 13266 12880 13322 12889
rect 13266 12815 13322 12824
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13280 10810 13308 12815
rect 13464 11354 13492 13942
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 12728 10662 12848 10690
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 9994 12664 10474
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12532 9920 12584 9926
rect 12584 9868 12664 9874
rect 12532 9862 12664 9868
rect 12544 9846 12664 9862
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12176 8362 12204 8842
rect 12348 8492 12400 8498
rect 12400 8452 12480 8480
rect 12348 8434 12400 8440
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12070 6896 12126 6905
rect 11980 6860 12032 6866
rect 12070 6831 12072 6840
rect 11980 6802 12032 6808
rect 12124 6831 12126 6840
rect 12072 6802 12124 6808
rect 12084 5658 12112 6802
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12162 6488 12218 6497
rect 12268 6458 12296 6734
rect 12452 6730 12480 8452
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12162 6423 12218 6432
rect 12256 6452 12308 6458
rect 12176 6186 12204 6423
rect 12256 6394 12308 6400
rect 12268 6322 12296 6394
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 11992 5642 12112 5658
rect 11980 5636 12112 5642
rect 12032 5630 12112 5636
rect 11980 5578 12032 5584
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 12268 5234 12296 6258
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 11704 4820 11756 4826
rect 11756 4780 11836 4808
rect 11704 4762 11756 4768
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11716 4146 11744 4626
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11808 3890 11836 4780
rect 11886 4720 11942 4729
rect 12268 4690 12296 5170
rect 11886 4655 11942 4664
rect 12256 4684 12308 4690
rect 11716 3862 11836 3890
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11624 2825 11652 2858
rect 11610 2816 11666 2825
rect 11610 2751 11666 2760
rect 11716 2774 11744 3862
rect 11900 3738 11928 4655
rect 12256 4626 12308 4632
rect 12360 4554 12388 6598
rect 12438 6488 12494 6497
rect 12438 6423 12440 6432
rect 12492 6423 12494 6432
rect 12440 6394 12492 6400
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 11980 4072 12032 4078
rect 12544 4026 12572 7754
rect 12636 5166 12664 9846
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 11980 4014 12032 4020
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11716 2746 11836 2774
rect 11532 1822 11652 1850
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 11624 800 11652 1822
rect 11808 1766 11836 2746
rect 11900 2582 11928 3062
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11992 1086 12020 4014
rect 12452 3998 12572 4026
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12452 3482 12480 3998
rect 12530 3632 12586 3641
rect 12530 3567 12586 3576
rect 12176 3466 12480 3482
rect 12544 3466 12572 3567
rect 12164 3460 12480 3466
rect 12216 3454 12480 3460
rect 12532 3460 12584 3466
rect 12164 3402 12216 3408
rect 12532 3402 12584 3408
rect 12636 3126 12664 4014
rect 12728 3777 12756 10406
rect 12820 8022 12848 10662
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12912 9042 12940 10610
rect 13268 10600 13320 10606
rect 12990 10568 13046 10577
rect 13268 10542 13320 10548
rect 12990 10503 13046 10512
rect 13004 9586 13032 10503
rect 13280 10198 13308 10542
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 9602 13308 10134
rect 13188 9586 13308 9602
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13176 9580 13308 9586
rect 13228 9574 13308 9580
rect 13176 9522 13228 9528
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12912 7886 12940 8978
rect 13188 8498 13216 9522
rect 13372 9364 13400 11086
rect 13450 10976 13506 10985
rect 13450 10911 13506 10920
rect 13464 10742 13492 10911
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13450 10024 13506 10033
rect 13450 9959 13506 9968
rect 13280 9353 13400 9364
rect 13266 9344 13400 9353
rect 13322 9336 13400 9344
rect 13266 9279 13322 9288
rect 13464 9194 13492 9959
rect 13556 9926 13584 17224
rect 13740 17134 13768 18838
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13648 15366 13676 15846
rect 13740 15638 13768 16934
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13726 14648 13782 14657
rect 13726 14583 13782 14592
rect 13740 14550 13768 14583
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13726 14376 13782 14385
rect 13726 14311 13728 14320
rect 13780 14311 13782 14320
rect 13728 14282 13780 14288
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13740 12646 13768 13670
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12434 13768 12582
rect 13648 12406 13768 12434
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13542 9616 13598 9625
rect 13542 9551 13598 9560
rect 13280 9166 13492 9194
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 7954 13216 8434
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12900 7880 12952 7886
rect 13280 7834 13308 9166
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13464 8566 13492 9046
rect 13556 8566 13584 9551
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13544 8424 13596 8430
rect 13648 8378 13676 12406
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 10062 13768 12242
rect 13832 11830 13860 17614
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13924 15094 13952 16730
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 14016 14822 14044 19306
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14108 13977 14136 28358
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14200 24682 14228 25230
rect 14384 24886 14412 26250
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14372 24880 14424 24886
rect 14372 24822 14424 24828
rect 14188 24676 14240 24682
rect 14188 24618 14240 24624
rect 14200 17678 14228 24618
rect 14476 24138 14504 25638
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14464 24132 14516 24138
rect 14464 24074 14516 24080
rect 14384 23594 14412 24074
rect 14372 23588 14424 23594
rect 14372 23530 14424 23536
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14384 20398 14412 21354
rect 14568 21010 14596 27814
rect 15028 24818 15056 32370
rect 15384 32224 15436 32230
rect 15384 32166 15436 32172
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15120 26314 15148 26930
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 15028 24274 15056 24754
rect 15120 24682 15148 26250
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15016 24268 15068 24274
rect 15016 24210 15068 24216
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14660 21978 14688 22578
rect 14752 22098 14780 22918
rect 15120 22778 15148 23734
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 14660 21950 14780 21978
rect 14752 21049 14780 21950
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14844 21729 14872 21898
rect 14830 21720 14886 21729
rect 14830 21655 14886 21664
rect 14738 21040 14794 21049
rect 14556 21004 14608 21010
rect 14738 20975 14794 20984
rect 14556 20946 14608 20952
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14280 19848 14332 19854
rect 14278 19816 14280 19825
rect 14332 19816 14334 19825
rect 14278 19751 14334 19760
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14292 17116 14320 19654
rect 14476 18766 14504 20198
rect 14568 19922 14596 20946
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19553 14688 19654
rect 14646 19544 14702 19553
rect 14646 19479 14702 19488
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14554 19272 14610 19281
rect 14554 19207 14556 19216
rect 14608 19207 14610 19216
rect 14556 19178 14608 19184
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14476 18193 14504 18702
rect 14568 18358 14596 18838
rect 14660 18834 14688 19382
rect 14752 19258 14780 20975
rect 14936 19446 14964 22034
rect 15028 21010 15056 22374
rect 15212 21706 15240 28970
rect 15396 27146 15424 32166
rect 15488 29170 15516 36518
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15580 28082 15608 36790
rect 15936 29096 15988 29102
rect 15936 29038 15988 29044
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15396 27118 15700 27146
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15120 21678 15240 21706
rect 15120 21468 15148 21678
rect 15200 21616 15252 21622
rect 15304 21570 15332 25094
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 23662 15424 24754
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15488 24274 15516 24550
rect 15580 24274 15608 26454
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15568 24268 15620 24274
rect 15568 24210 15620 24216
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15396 22094 15424 23598
rect 15396 22066 15516 22094
rect 15252 21564 15332 21570
rect 15200 21558 15332 21564
rect 15212 21542 15332 21558
rect 15200 21480 15252 21486
rect 15120 21440 15200 21468
rect 15200 21422 15252 21428
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15014 20360 15070 20369
rect 15014 20295 15016 20304
rect 15068 20295 15070 20304
rect 15016 20266 15068 20272
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14752 19230 14964 19258
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14556 18352 14608 18358
rect 14556 18294 14608 18300
rect 14462 18184 14518 18193
rect 14462 18119 14518 18128
rect 14556 18148 14608 18154
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14200 17088 14320 17116
rect 14200 16046 14228 17088
rect 14384 16726 14412 17818
rect 14476 16980 14504 18119
rect 14556 18090 14608 18096
rect 14568 17134 14596 18090
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14476 16952 14596 16980
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14462 16688 14518 16697
rect 14462 16623 14464 16632
rect 14516 16623 14518 16632
rect 14464 16594 14516 16600
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 15910 14228 15982
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14200 14006 14228 14554
rect 14188 14000 14240 14006
rect 14094 13968 14150 13977
rect 13912 13932 13964 13938
rect 14188 13942 14240 13948
rect 14094 13903 14150 13912
rect 13912 13874 13964 13880
rect 13924 13274 13952 13874
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14108 13569 14136 13806
rect 14094 13560 14150 13569
rect 14094 13495 14150 13504
rect 13924 13246 14228 13274
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13832 10810 13860 11630
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13924 9654 13952 12106
rect 14016 10606 14044 13126
rect 14200 12442 14228 13246
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13596 8372 13676 8378
rect 13544 8366 13676 8372
rect 13556 8350 13676 8366
rect 12900 7822 12952 7828
rect 13188 7806 13308 7834
rect 12806 7032 12862 7041
rect 12806 6967 12862 6976
rect 12820 5710 12848 6967
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 13188 5302 13216 7806
rect 13266 7712 13322 7721
rect 13266 7647 13322 7656
rect 13280 7478 13308 7647
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 13280 5030 13308 7239
rect 13740 6662 13768 8774
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 5914 13676 6258
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13084 3936 13136 3942
rect 12806 3904 12862 3913
rect 13084 3878 13136 3884
rect 12806 3839 12862 3848
rect 12714 3768 12770 3777
rect 12820 3738 12848 3839
rect 12714 3703 12770 3712
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12360 2514 12388 2926
rect 12636 2825 12664 2926
rect 12622 2816 12678 2825
rect 12622 2751 12678 2760
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12176 1494 12204 2314
rect 12164 1488 12216 1494
rect 12164 1430 12216 1436
rect 11980 1080 12032 1086
rect 11980 1022 12032 1028
rect 12912 800 12940 3674
rect 13096 3641 13124 3878
rect 13082 3632 13138 3641
rect 13082 3567 13138 3576
rect 13280 1222 13308 4150
rect 13556 4078 13584 5782
rect 13726 5672 13782 5681
rect 13726 5607 13782 5616
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13648 3482 13676 4966
rect 13740 4078 13768 5607
rect 13832 4758 13860 9279
rect 14108 6390 14136 12310
rect 14292 12050 14320 15438
rect 14568 15201 14596 16952
rect 14554 15192 14610 15201
rect 14554 15127 14610 15136
rect 14660 15065 14688 17614
rect 14646 15056 14702 15065
rect 14646 14991 14702 15000
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14482 14596 14758
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14462 14240 14518 14249
rect 14462 14175 14518 14184
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14384 13258 14412 13466
rect 14476 13258 14504 14175
rect 14648 14000 14700 14006
rect 14646 13968 14648 13977
rect 14700 13968 14702 13977
rect 14646 13903 14702 13912
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14752 12918 14780 19110
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 16454 14872 17478
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14200 12022 14320 12050
rect 14462 12064 14518 12073
rect 14200 11694 14228 12022
rect 14462 11999 14518 12008
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14200 9178 14228 11630
rect 14292 11218 14320 11766
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 14292 9178 14320 10678
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14384 8634 14412 11698
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14002 5264 14058 5273
rect 14002 5199 14058 5208
rect 14016 5098 14044 5199
rect 14384 5166 14412 5510
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 13820 4752 13872 4758
rect 13818 4720 13820 4729
rect 13872 4720 13874 4729
rect 13818 4655 13874 4664
rect 14278 4720 14334 4729
rect 14278 4655 14334 4664
rect 14292 4622 14320 4655
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13740 3670 13768 4014
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13544 3460 13596 3466
rect 13648 3454 13768 3482
rect 13544 3402 13596 3408
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13372 1578 13400 2790
rect 13556 2009 13584 3402
rect 13740 3398 13768 3454
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 14476 3126 14504 11999
rect 14568 11762 14596 12786
rect 14752 12374 14780 12854
rect 14740 12368 14792 12374
rect 14646 12336 14702 12345
rect 14740 12310 14792 12316
rect 14646 12271 14702 12280
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14556 11620 14608 11626
rect 14660 11608 14688 12271
rect 14608 11580 14688 11608
rect 14556 11562 14608 11568
rect 14554 11384 14610 11393
rect 14554 11319 14610 11328
rect 14568 11218 14596 11319
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14844 11121 14872 14282
rect 14830 11112 14886 11121
rect 14830 11047 14886 11056
rect 14740 11008 14792 11014
rect 14738 10976 14740 10985
rect 14792 10976 14794 10985
rect 14738 10911 14794 10920
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14752 7818 14780 9930
rect 14844 9353 14872 11047
rect 14830 9344 14886 9353
rect 14830 9279 14886 9288
rect 14936 8294 14964 19230
rect 15028 10849 15056 20266
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 17882 15148 19722
rect 15212 19446 15240 21422
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15396 20398 15424 20878
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15292 18624 15344 18630
rect 15396 18612 15424 20334
rect 15344 18584 15424 18612
rect 15292 18566 15344 18572
rect 15304 18426 15332 18566
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15120 17338 15148 17546
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15120 17066 15148 17274
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15212 16114 15240 16934
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15014 10840 15070 10849
rect 15014 10775 15070 10784
rect 15014 10160 15070 10169
rect 15014 10095 15070 10104
rect 15028 9586 15056 10095
rect 15120 9994 15148 14010
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15212 13258 15240 13874
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15304 12209 15332 16186
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15396 13870 15424 15506
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15382 13696 15438 13705
rect 15382 13631 15438 13640
rect 15396 13530 15424 13631
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15290 12200 15346 12209
rect 15290 12135 15346 12144
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 10577 15240 12038
rect 15198 10568 15254 10577
rect 15198 10503 15254 10512
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15106 9888 15162 9897
rect 15212 9874 15240 10134
rect 15304 9926 15332 12135
rect 15162 9846 15240 9874
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15106 9823 15162 9832
rect 15396 9738 15424 9862
rect 15120 9710 15424 9738
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14752 6866 14780 7754
rect 15028 7698 15056 8570
rect 15120 8090 15148 9710
rect 15488 9178 15516 22066
rect 15580 21350 15608 23802
rect 15672 22778 15700 27118
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15764 22710 15792 24550
rect 15856 24342 15884 24686
rect 15844 24336 15896 24342
rect 15844 24278 15896 24284
rect 15752 22704 15804 22710
rect 15948 22658 15976 29038
rect 16132 23730 16160 37266
rect 16500 37210 16528 39222
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 16580 37664 16632 37670
rect 16580 37606 16632 37612
rect 16592 37398 16620 37606
rect 16580 37392 16632 37398
rect 16580 37334 16632 37340
rect 16500 37194 16620 37210
rect 16500 37188 16632 37194
rect 16500 37182 16580 37188
rect 16580 37130 16632 37136
rect 16776 36786 16804 39200
rect 18064 37262 18092 39200
rect 19156 37664 19208 37670
rect 19156 37606 19208 37612
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 16764 36780 16816 36786
rect 16764 36722 16816 36728
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16304 27056 16356 27062
rect 16304 26998 16356 27004
rect 16316 24070 16344 26998
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 15752 22646 15804 22652
rect 15856 22630 15976 22658
rect 15856 22574 15884 22630
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15580 19666 15608 21286
rect 15856 21010 15884 22510
rect 16316 22098 16344 24006
rect 16592 23254 16620 29582
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16960 24886 16988 25094
rect 16948 24880 17000 24886
rect 16948 24822 17000 24828
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 24274 16988 24550
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16304 22092 16356 22098
rect 16304 22034 16356 22040
rect 16028 21956 16080 21962
rect 16028 21898 16080 21904
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16040 21350 16068 21898
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16040 21078 16068 21286
rect 16028 21072 16080 21078
rect 16028 21014 16080 21020
rect 16120 21072 16172 21078
rect 16120 21014 16172 21020
rect 15844 21004 15896 21010
rect 15844 20946 15896 20952
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15672 19854 15700 19994
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15580 19638 15700 19666
rect 15566 19544 15622 19553
rect 15566 19479 15622 19488
rect 15580 19446 15608 19479
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 16522 15608 18566
rect 15672 17814 15700 19638
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15672 16697 15700 17070
rect 15658 16688 15714 16697
rect 15658 16623 15714 16632
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15764 16250 15792 20402
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 18834 15884 20198
rect 16132 19922 16160 21014
rect 16316 20466 16344 21490
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16592 20058 16620 21286
rect 16684 20534 16712 21898
rect 16868 21010 16896 22374
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16776 20602 16804 20810
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16026 18864 16082 18873
rect 15844 18828 15896 18834
rect 16026 18799 16082 18808
rect 15844 18770 15896 18776
rect 16040 18766 16068 18799
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16132 18465 16160 18702
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16118 18456 16174 18465
rect 16118 18391 16174 18400
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16224 17882 16252 18090
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16316 17270 16344 18566
rect 16684 18222 16712 19178
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16304 17264 16356 17270
rect 16304 17206 16356 17212
rect 16118 17096 16174 17105
rect 16118 17031 16174 17040
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 13852 15608 15574
rect 15672 15162 15700 15642
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15672 14074 15700 14282
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15764 14006 15792 14214
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15844 13864 15896 13870
rect 15580 13824 15792 13852
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15672 12306 15700 12922
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 10606 15700 12242
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10130 15700 10542
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 15476 8900 15528 8906
rect 15580 8888 15608 9114
rect 15528 8860 15608 8888
rect 15476 8842 15528 8848
rect 15382 8528 15438 8537
rect 15382 8463 15438 8472
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14936 7670 15056 7698
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14752 6730 14780 6802
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5710 14688 6054
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14646 5400 14702 5409
rect 14646 5335 14648 5344
rect 14700 5335 14702 5344
rect 14648 5306 14700 5312
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14568 4078 14596 4558
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14568 3602 14596 4014
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14568 3058 14596 3538
rect 14752 3534 14780 6666
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13542 2000 13598 2009
rect 13648 1970 13676 2586
rect 13740 2553 13768 2994
rect 13726 2544 13782 2553
rect 14568 2514 14596 2994
rect 13726 2479 13782 2488
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13542 1935 13598 1944
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 13740 1873 13768 2314
rect 13726 1864 13782 1873
rect 13726 1799 13782 1808
rect 13372 1550 13584 1578
rect 13268 1216 13320 1222
rect 13268 1158 13320 1164
rect 13556 800 13584 1550
rect 14844 800 14872 4422
rect 14936 4214 14964 7670
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15028 7449 15056 7482
rect 15014 7440 15070 7449
rect 15014 7375 15016 7384
rect 15068 7375 15070 7384
rect 15016 7346 15068 7352
rect 15120 7206 15148 7754
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6798 15148 7142
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 5710 15148 6734
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 5166 15148 5646
rect 15304 5642 15332 6258
rect 15396 5642 15424 8463
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14936 2854 14964 4150
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 15396 2774 15424 5578
rect 15764 5302 15792 13824
rect 15844 13806 15896 13812
rect 15856 13258 15884 13806
rect 15948 13462 15976 16118
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15856 9654 15884 13194
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15948 10849 15976 11154
rect 15934 10840 15990 10849
rect 15934 10775 15990 10784
rect 16040 9674 16068 16662
rect 16132 13530 16160 17031
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 11558 16160 12718
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15948 9646 16068 9674
rect 15948 6610 15976 9646
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 9042 16160 9386
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16132 8498 16160 8978
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 7954 16160 8434
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 15856 6582 15976 6610
rect 15856 6322 15884 6582
rect 16224 6474 16252 16050
rect 16408 15570 16436 17478
rect 16500 16522 16528 18090
rect 16776 18086 16804 20402
rect 16960 19922 16988 21286
rect 17052 21078 17080 31962
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17316 28960 17368 28966
rect 17316 28902 17368 28908
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17236 25294 17264 26182
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 17144 22710 17172 25094
rect 17132 22704 17184 22710
rect 17132 22646 17184 22652
rect 17328 22094 17356 28902
rect 17880 25906 17908 30194
rect 18064 28558 18092 37062
rect 18432 36922 18460 37198
rect 18420 36916 18472 36922
rect 18420 36858 18472 36864
rect 18236 31884 18288 31890
rect 18236 31826 18288 31832
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 18144 28416 18196 28422
rect 18144 28358 18196 28364
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 18064 25226 18092 25638
rect 18052 25220 18104 25226
rect 18052 25162 18104 25168
rect 18064 24750 18092 25162
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17972 24138 18000 24618
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17420 22166 17448 22442
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17236 22066 17356 22094
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17236 19786 17264 22066
rect 17420 21010 17448 22102
rect 17512 21690 17540 23258
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17604 20913 17632 21082
rect 17590 20904 17646 20913
rect 17500 20868 17552 20874
rect 17590 20839 17646 20848
rect 17500 20810 17552 20816
rect 17512 20097 17540 20810
rect 17696 20330 17724 22170
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17788 21418 17816 21898
rect 17880 21690 17908 23598
rect 17972 23594 18000 24074
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17498 20088 17554 20097
rect 17498 20023 17554 20032
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17236 19666 17264 19722
rect 17144 19638 17264 19666
rect 16946 19136 17002 19145
rect 16946 19071 17002 19080
rect 16960 18970 16988 19071
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16408 15026 16436 15506
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16500 14958 16528 16458
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16316 14006 16344 14486
rect 16500 14482 16528 14894
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16316 12866 16344 13466
rect 16408 12986 16436 14282
rect 16500 13190 16528 14282
rect 16592 13258 16620 16934
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 14958 16712 16594
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16776 15706 16804 15914
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16868 15570 16896 18906
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16948 18352 17000 18358
rect 17052 18340 17080 18566
rect 17000 18312 17080 18340
rect 16948 18294 17000 18300
rect 17144 17678 17172 19638
rect 17512 19417 17540 19722
rect 17604 19446 17632 19722
rect 17592 19440 17644 19446
rect 17498 19408 17554 19417
rect 17592 19382 17644 19388
rect 17696 19378 17724 20266
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17498 19343 17554 19352
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17222 19272 17278 19281
rect 17222 19207 17224 19216
rect 17276 19207 17278 19216
rect 17224 19178 17276 19184
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17236 17202 17264 18702
rect 17420 18358 17448 18770
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17316 18216 17368 18222
rect 17314 18184 17316 18193
rect 17368 18184 17370 18193
rect 17314 18119 17370 18128
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17224 17196 17276 17202
rect 17224 17138 17276 17144
rect 17132 16584 17184 16590
rect 16946 16552 17002 16561
rect 17132 16526 17184 16532
rect 16946 16487 17002 16496
rect 16856 15564 16908 15570
rect 16856 15506 16908 15512
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16684 13530 16712 13738
rect 16776 13705 16804 14418
rect 16762 13696 16818 13705
rect 16762 13631 16818 13640
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16316 12838 16528 12866
rect 16868 12850 16896 14758
rect 16316 12782 16344 12838
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16316 11898 16344 12378
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16408 11937 16436 12106
rect 16394 11928 16450 11937
rect 16304 11892 16356 11898
rect 16394 11863 16450 11872
rect 16304 11834 16356 11840
rect 16500 10742 16528 12838
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16672 12300 16724 12306
rect 16868 12288 16896 12786
rect 16724 12260 16896 12288
rect 16672 12242 16724 12248
rect 16684 11762 16712 12242
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 9353 16344 9522
rect 16302 9344 16358 9353
rect 16302 9279 16358 9288
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 15948 6458 16252 6474
rect 15936 6452 16252 6458
rect 15988 6446 16252 6452
rect 15936 6394 15988 6400
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16132 6225 16160 6258
rect 16118 6216 16174 6225
rect 16118 6151 16174 6160
rect 15842 5944 15898 5953
rect 15842 5879 15898 5888
rect 15856 5778 15884 5879
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15396 2746 15516 2774
rect 15488 2650 15516 2746
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15948 1578 15976 5714
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4690 16344 4966
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16408 4570 16436 8978
rect 16500 7993 16528 10406
rect 16672 9988 16724 9994
rect 16672 9930 16724 9936
rect 16684 9518 16712 9930
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16578 9208 16634 9217
rect 16868 9178 16896 11290
rect 16578 9143 16580 9152
rect 16632 9143 16634 9152
rect 16856 9172 16908 9178
rect 16580 9114 16632 9120
rect 16856 9114 16908 9120
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8634 16712 8910
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16960 8430 16988 16487
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 14006 17080 16390
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17052 13025 17080 13126
rect 17038 13016 17094 13025
rect 17038 12951 17094 12960
rect 17040 12776 17092 12782
rect 17038 12744 17040 12753
rect 17092 12744 17094 12753
rect 17038 12679 17094 12688
rect 17040 11688 17092 11694
rect 17040 11630 17092 11636
rect 17052 11014 17080 11630
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17144 10606 17172 16526
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 10470 17172 10542
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17132 9512 17184 9518
rect 17130 9480 17132 9489
rect 17184 9480 17186 9489
rect 17130 9415 17186 9424
rect 17236 9382 17264 17138
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17328 14822 17356 16050
rect 17420 15094 17448 17478
rect 17512 16250 17540 17546
rect 17604 17513 17632 17546
rect 17590 17504 17646 17513
rect 17590 17439 17646 17448
rect 17682 17368 17738 17377
rect 17682 17303 17738 17312
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17604 16794 17632 16934
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17604 15910 17632 16526
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17408 15088 17460 15094
rect 17408 15030 17460 15036
rect 17498 15056 17554 15065
rect 17498 14991 17554 15000
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17328 14414 17356 14758
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17328 11082 17356 13330
rect 17420 13258 17448 14554
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17512 11354 17540 14991
rect 17696 14958 17724 17303
rect 17788 15978 17816 20198
rect 17880 19310 17908 21626
rect 18050 19816 18106 19825
rect 18050 19751 18106 19760
rect 18064 19446 18092 19751
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17880 16046 17908 19110
rect 17972 16522 18000 19382
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17270 18092 18022
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 16153 18092 16390
rect 18050 16144 18106 16153
rect 17960 16108 18012 16114
rect 18050 16079 18106 16088
rect 17960 16050 18012 16056
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17776 15972 17828 15978
rect 17776 15914 17828 15920
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15434 17908 15846
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17972 15337 18000 16050
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 17958 15328 18014 15337
rect 17958 15263 18014 15272
rect 18064 15178 18092 15982
rect 18156 15570 18184 28358
rect 18248 22098 18276 31826
rect 19064 26376 19116 26382
rect 19064 26318 19116 26324
rect 19076 25906 19104 26318
rect 19064 25900 19116 25906
rect 19064 25842 19116 25848
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 18340 25226 18368 25638
rect 18328 25220 18380 25226
rect 18328 25162 18380 25168
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18340 23050 18368 24006
rect 18892 23730 18920 24142
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18512 23588 18564 23594
rect 18512 23530 18564 23536
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 18236 22092 18288 22098
rect 18236 22034 18288 22040
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18248 17610 18276 19246
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18248 15337 18276 16050
rect 18234 15328 18290 15337
rect 18234 15263 18290 15272
rect 18064 15150 18276 15178
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17604 10470 17632 14894
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17314 9752 17370 9761
rect 17314 9687 17370 9696
rect 17500 9716 17552 9722
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16486 7984 16542 7993
rect 16960 7970 16988 8366
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 16960 7942 17080 7970
rect 16486 7919 16542 7928
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 7200 16816 7206
rect 16486 7168 16542 7177
rect 16764 7142 16816 7148
rect 16486 7103 16542 7112
rect 16500 5710 16528 7103
rect 16670 6760 16726 6769
rect 16670 6695 16672 6704
rect 16724 6695 16726 6704
rect 16672 6666 16724 6672
rect 16776 6254 16804 7142
rect 16868 6458 16896 7278
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16868 6322 16896 6394
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16316 4542 16436 4570
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16040 2514 16068 2926
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16132 2310 16160 3402
rect 16316 2990 16344 4542
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16316 1698 16344 2246
rect 16304 1692 16356 1698
rect 16304 1634 16356 1640
rect 15948 1550 16160 1578
rect 16132 800 16160 1550
rect 16408 1154 16436 4150
rect 16592 3913 16620 4626
rect 16578 3904 16634 3913
rect 16578 3839 16634 3848
rect 16578 3632 16634 3641
rect 16684 3602 16712 6054
rect 16764 5840 16816 5846
rect 16764 5782 16816 5788
rect 16578 3567 16580 3576
rect 16632 3567 16634 3576
rect 16672 3596 16724 3602
rect 16580 3538 16632 3544
rect 16672 3538 16724 3544
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16500 2825 16528 3062
rect 16486 2816 16542 2825
rect 16486 2751 16542 2760
rect 16396 1148 16448 1154
rect 16396 1090 16448 1096
rect 16776 800 16804 5782
rect 17052 5778 17080 7942
rect 17144 6254 17172 8026
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17236 6254 17264 6326
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17328 4690 17356 9687
rect 17500 9658 17552 9664
rect 17512 9518 17540 9658
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8430 17632 9318
rect 17696 8906 17724 14758
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17788 14482 17816 14554
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17788 10810 17816 13942
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17774 9208 17830 9217
rect 17880 9178 17908 13194
rect 17960 12776 18012 12782
rect 18012 12736 18092 12764
rect 17960 12718 18012 12724
rect 18064 11762 18092 12736
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18064 11286 18092 11698
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 18156 10198 18184 13874
rect 18248 12782 18276 15150
rect 18340 13258 18368 22374
rect 18432 21962 18460 23462
rect 18524 23186 18552 23530
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18420 21956 18472 21962
rect 18420 21898 18472 21904
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18616 21457 18644 21490
rect 18602 21448 18658 21457
rect 18602 21383 18658 21392
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18432 18057 18460 18226
rect 18418 18048 18474 18057
rect 18418 17983 18474 17992
rect 18524 17678 18552 18702
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18418 16824 18474 16833
rect 18418 16759 18474 16768
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18248 12345 18276 12718
rect 18234 12336 18290 12345
rect 18234 12271 18290 12280
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11608 18368 12038
rect 18248 11580 18368 11608
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 17774 9143 17830 9152
rect 17868 9172 17920 9178
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17696 6662 17724 8026
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17498 5808 17554 5817
rect 17498 5743 17554 5752
rect 17512 5710 17540 5743
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17144 4214 17172 4490
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16868 3058 16896 4014
rect 17788 3670 17816 9143
rect 17868 9114 17920 9120
rect 18248 9081 18276 11580
rect 18326 11384 18382 11393
rect 18326 11319 18328 11328
rect 18380 11319 18382 11328
rect 18328 11290 18380 11296
rect 18432 9110 18460 16759
rect 18524 16726 18552 17614
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18616 15178 18644 20538
rect 18694 18592 18750 18601
rect 18694 18527 18750 18536
rect 18708 18290 18736 18527
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18524 15150 18644 15178
rect 18524 13190 18552 15150
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18616 12170 18644 15030
rect 18708 13734 18736 16526
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 9104 18472 9110
rect 18234 9072 18290 9081
rect 18290 9030 18368 9058
rect 18420 9046 18472 9052
rect 18234 9007 18290 9016
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17868 5160 17920 5166
rect 17866 5128 17868 5137
rect 17920 5128 17922 5137
rect 17866 5063 17922 5072
rect 17972 4622 18000 6598
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18064 4486 18092 7686
rect 18156 5409 18184 7958
rect 18234 6896 18290 6905
rect 18234 6831 18290 6840
rect 18248 6322 18276 6831
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18340 6186 18368 9030
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18142 5400 18198 5409
rect 18142 5335 18198 5344
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17788 3194 17816 3470
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17144 2514 17172 2994
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 17328 2038 17356 2314
rect 17316 2032 17368 2038
rect 17316 1974 17368 1980
rect 17972 1902 18000 3402
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18156 2774 18184 3334
rect 18432 2854 18460 8910
rect 18524 7886 18552 11630
rect 18708 10062 18736 12718
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18616 8362 18644 9318
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18616 7342 18644 8298
rect 18708 8022 18736 9318
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18800 7818 18828 15642
rect 18892 12102 18920 23666
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18984 16726 19012 17070
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18984 14278 19012 15914
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18878 11520 18934 11529
rect 18878 11455 18934 11464
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18694 7304 18750 7313
rect 18694 7239 18750 7248
rect 18708 7002 18736 7239
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18616 4690 18644 4966
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18708 4026 18736 6938
rect 18800 6361 18828 7142
rect 18786 6352 18842 6361
rect 18786 6287 18842 6296
rect 18892 5114 18920 11455
rect 18984 9382 19012 13126
rect 19076 11694 19104 25842
rect 19168 20602 19196 37606
rect 19352 36922 19380 39200
rect 19996 37126 20024 39200
rect 21284 37262 21312 39200
rect 22572 37330 22600 39200
rect 22560 37324 22612 37330
rect 22560 37266 22612 37272
rect 21272 37256 21324 37262
rect 21272 37198 21324 37204
rect 21088 37188 21140 37194
rect 21088 37130 21140 37136
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 20352 37120 20404 37126
rect 20352 37062 20404 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19352 22710 19380 25162
rect 19444 23322 19472 36722
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19628 24138 19656 24210
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19168 20466 19196 20538
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 19168 17338 19196 17546
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19260 16794 19288 17206
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19260 15026 19288 16118
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19168 14074 19196 14894
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19260 14006 19288 14282
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19352 13870 19380 21558
rect 19444 20058 19472 21830
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 19720 21350 19748 21490
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19628 20874 19656 21286
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19444 18034 19472 19382
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19536 18834 19564 19246
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19444 18006 19564 18034
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19444 17066 19472 17818
rect 19536 17678 19564 18006
rect 19628 17678 19656 18226
rect 19524 17672 19576 17678
rect 19522 17640 19524 17649
rect 19616 17672 19668 17678
rect 19576 17640 19578 17649
rect 19616 17614 19668 17620
rect 19996 17626 20024 33798
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 20088 22098 20116 31826
rect 20364 31822 20392 37062
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20640 31822 20668 34886
rect 20812 32292 20864 32298
rect 20812 32234 20864 32240
rect 20824 31822 20852 32234
rect 20352 31816 20404 31822
rect 20352 31758 20404 31764
rect 20628 31816 20680 31822
rect 20628 31758 20680 31764
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 21100 31754 21128 37130
rect 23020 37120 23072 37126
rect 23216 37108 23244 39200
rect 23572 37392 23624 37398
rect 23572 37334 23624 37340
rect 23216 37080 23520 37108
rect 23020 37062 23072 37068
rect 21640 36576 21692 36582
rect 21640 36518 21692 36524
rect 21652 31822 21680 36518
rect 23032 31822 23060 37062
rect 23492 36786 23520 37080
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 20916 31726 21128 31754
rect 20536 26920 20588 26926
rect 20536 26862 20588 26868
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20180 22098 20208 24210
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 20272 22642 20300 22918
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20364 22574 20392 26522
rect 20548 24274 20576 26862
rect 20536 24268 20588 24274
rect 20536 24210 20588 24216
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20180 20806 20208 22034
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20456 20584 20484 23598
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20180 20556 20484 20584
rect 20180 20330 20208 20556
rect 20548 20482 20576 22646
rect 20640 22642 20668 23122
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20272 20454 20576 20482
rect 20640 20466 20668 22578
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20732 21010 20760 21354
rect 20824 21350 20852 23054
rect 20916 21554 20944 31726
rect 23124 28966 23152 31962
rect 23584 30394 23612 37334
rect 24504 37262 24532 39200
rect 24860 37324 24912 37330
rect 24860 37266 24912 37272
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23112 28960 23164 28966
rect 23112 28902 23164 28908
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21652 23118 21680 25298
rect 21640 23112 21692 23118
rect 21638 23080 21640 23089
rect 21692 23080 21694 23089
rect 21638 23015 21694 23024
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21468 22642 21496 22918
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 21008 21010 21036 22374
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21100 21690 21128 21898
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20996 21004 21048 21010
rect 20996 20946 21048 20952
rect 20628 20460 20680 20466
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 19996 17598 20116 17626
rect 19522 17575 19578 17584
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19812 16794 19840 17070
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19904 16794 19932 16934
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 14278 19472 15846
rect 19996 15434 20024 17478
rect 20088 16658 20116 17598
rect 20272 17338 20300 20454
rect 20628 20402 20680 20408
rect 20640 20346 20668 20402
rect 20732 20398 20760 20946
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20548 20318 20668 20346
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 20058 20392 20198
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19536 14346 19564 15098
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19812 14822 19840 14962
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19248 13864 19300 13870
rect 19246 13832 19248 13841
rect 19340 13864 19392 13870
rect 19300 13832 19302 13841
rect 19340 13806 19392 13812
rect 19246 13767 19302 13776
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 19798 13424 19854 13433
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18984 8294 19012 9046
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18984 7750 19012 7890
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18970 6080 19026 6089
rect 18970 6015 19026 6024
rect 18800 5098 18920 5114
rect 18788 5092 18920 5098
rect 18840 5086 18920 5092
rect 18788 5034 18840 5040
rect 18800 4554 18828 5034
rect 18984 4672 19012 6015
rect 19076 5302 19104 11018
rect 19168 10742 19196 13398
rect 19798 13359 19854 13368
rect 19812 13258 19840 13359
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19800 13252 19852 13258
rect 19800 13194 19852 13200
rect 19444 12646 19472 13194
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19432 12368 19484 12374
rect 19430 12336 19432 12345
rect 19484 12336 19486 12345
rect 19430 12271 19486 12280
rect 19708 12164 19760 12170
rect 19352 12124 19708 12152
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11286 19288 12038
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19260 10606 19288 11222
rect 19352 10810 19380 12124
rect 19708 12106 19760 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19536 10996 19564 11766
rect 19444 10968 19564 10996
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19168 7721 19196 9386
rect 19260 9024 19288 10542
rect 19444 10198 19472 10968
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19444 9518 19472 9998
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9654 20024 14214
rect 20088 10606 20116 15302
rect 20180 15162 20208 17002
rect 20364 16182 20392 18566
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20456 17270 20484 18022
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20548 17116 20576 20318
rect 20824 20058 20852 20742
rect 21100 20534 21128 21490
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20640 17626 20668 19994
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20916 18766 20944 19178
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20640 17598 20760 17626
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20456 17088 20576 17116
rect 20456 16538 20484 17088
rect 20534 16688 20590 16697
rect 20534 16623 20536 16632
rect 20588 16623 20590 16632
rect 20536 16594 20588 16600
rect 20456 16510 20576 16538
rect 20640 16522 20668 17478
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20444 16176 20496 16182
rect 20444 16118 20496 16124
rect 20456 15502 20484 16118
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20180 13734 20208 14826
rect 20272 14362 20300 15098
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20350 14512 20406 14521
rect 20350 14447 20352 14456
rect 20404 14447 20406 14456
rect 20352 14418 20404 14424
rect 20272 14334 20392 14362
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19340 9036 19392 9042
rect 19260 8996 19340 9024
rect 19340 8978 19392 8984
rect 19444 8634 19472 9454
rect 19708 9104 19760 9110
rect 19706 9072 19708 9081
rect 19760 9072 19762 9081
rect 19706 9007 19762 9016
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19536 8498 19564 8570
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19536 7954 19564 8434
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 7732 19564 7890
rect 19890 7848 19946 7857
rect 19890 7783 19892 7792
rect 19944 7783 19946 7792
rect 19892 7754 19944 7760
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 19444 7704 19564 7732
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19352 6458 19380 7278
rect 19444 6866 19472 7704
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19800 7472 19852 7478
rect 19996 7460 20024 9590
rect 19800 7414 19852 7420
rect 19904 7432 20024 7460
rect 19812 7342 19840 7414
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19522 6896 19578 6905
rect 19432 6860 19484 6866
rect 19522 6831 19578 6840
rect 19432 6802 19484 6808
rect 19536 6746 19564 6831
rect 19444 6718 19564 6746
rect 19904 6730 19932 7432
rect 19892 6724 19944 6730
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19352 6254 19380 6394
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19064 5296 19116 5302
rect 19064 5238 19116 5244
rect 18892 4644 19012 4672
rect 19156 4684 19208 4690
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18616 3998 18736 4026
rect 18616 3942 18644 3998
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18064 2746 18184 2774
rect 17960 1896 18012 1902
rect 17960 1838 18012 1844
rect 18064 800 18092 2746
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18432 1766 18460 2518
rect 18892 1834 18920 4644
rect 19156 4626 19208 4632
rect 18972 4548 19024 4554
rect 18972 4490 19024 4496
rect 18984 4078 19012 4490
rect 19168 4146 19196 4626
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19076 2990 19104 4014
rect 19168 3602 19196 4082
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19168 3058 19196 3538
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19168 2514 19196 2994
rect 19260 2666 19288 6190
rect 19352 5778 19380 6190
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5302 19380 5714
rect 19444 5302 19472 6718
rect 19892 6666 19944 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 20088 6458 20116 10542
rect 20180 9722 20208 13194
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20180 8809 20208 8842
rect 20166 8800 20222 8809
rect 20166 8735 20222 8744
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 19982 5536 20038 5545
rect 19574 5468 19882 5477
rect 19982 5471 20038 5480
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19352 4622 19380 5238
rect 19430 4992 19486 5001
rect 19430 4927 19486 4936
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4214 19380 4422
rect 19444 4214 19472 4927
rect 19996 4554 20024 5471
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19984 3460 20036 3466
rect 20088 3448 20116 5607
rect 20168 4208 20220 4214
rect 20272 4196 20300 14010
rect 20364 13802 20392 14334
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20364 13569 20392 13738
rect 20350 13560 20406 13569
rect 20350 13495 20406 13504
rect 20350 13288 20406 13297
rect 20350 13223 20406 13232
rect 20364 12782 20392 13223
rect 20456 12850 20484 14962
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20364 7002 20392 12718
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20456 7698 20484 12582
rect 20548 12102 20576 16510
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20732 16402 20760 17598
rect 20824 16658 20852 17750
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20916 16561 20944 16594
rect 20902 16552 20958 16561
rect 20902 16487 20958 16496
rect 20640 16374 20760 16402
rect 20640 16182 20668 16374
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20720 15496 20772 15502
rect 20718 15464 20720 15473
rect 20772 15464 20774 15473
rect 20718 15399 20774 15408
rect 20732 14618 20760 15399
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20810 14104 20866 14113
rect 20810 14039 20866 14048
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20640 9874 20668 13806
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20732 13258 20760 13738
rect 20824 13394 20852 14039
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20718 12880 20774 12889
rect 20718 12815 20720 12824
rect 20772 12815 20774 12824
rect 20720 12786 20772 12792
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12170 20852 12582
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20548 9846 20668 9874
rect 20548 8673 20576 9846
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20534 8664 20590 8673
rect 20534 8599 20590 8608
rect 20456 7670 20576 7698
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20456 7002 20484 7482
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20350 6624 20406 6633
rect 20350 6559 20406 6568
rect 20364 5273 20392 6559
rect 20350 5264 20406 5273
rect 20350 5199 20406 5208
rect 20220 4168 20300 4196
rect 20168 4150 20220 4156
rect 20548 3942 20576 7670
rect 20640 6905 20668 9658
rect 20732 9625 20760 12038
rect 20916 11694 20944 15506
rect 21008 12434 21036 18634
rect 21100 18290 21128 18906
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 21192 15094 21220 21898
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21284 21146 21312 21490
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19854 21496 20198
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21456 18284 21508 18290
rect 21456 18226 21508 18232
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21284 16046 21312 17070
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21284 14890 21312 15982
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21088 14816 21140 14822
rect 21140 14764 21220 14770
rect 21088 14758 21220 14764
rect 21100 14742 21220 14758
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 21100 13172 21128 13942
rect 21192 13410 21220 14742
rect 21376 13870 21404 15982
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21468 13682 21496 18226
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 13977 21588 14350
rect 21546 13968 21602 13977
rect 21546 13903 21602 13912
rect 21468 13654 21588 13682
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21192 13382 21404 13410
rect 21376 13326 21404 13382
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 13184 21324 13190
rect 21100 13144 21272 13172
rect 21272 13126 21324 13132
rect 21468 12850 21496 13466
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21008 12406 21404 12434
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21100 11937 21128 12310
rect 21284 12209 21312 12310
rect 21270 12200 21326 12209
rect 21270 12135 21326 12144
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21086 11928 21142 11937
rect 21284 11898 21312 12038
rect 21086 11863 21142 11872
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21086 11792 21142 11801
rect 21086 11727 21142 11736
rect 21270 11792 21326 11801
rect 21270 11727 21326 11736
rect 21100 11694 21128 11727
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20718 9616 20774 9625
rect 20718 9551 20774 9560
rect 20732 7970 20760 9551
rect 20916 9450 20944 11630
rect 21284 11558 21312 11727
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21376 11354 21404 12406
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21086 11248 21142 11257
rect 21086 11183 21142 11192
rect 21100 11150 21128 11183
rect 21088 11144 21140 11150
rect 21284 11121 21312 11290
rect 21088 11086 21140 11092
rect 21270 11112 21326 11121
rect 21270 11047 21326 11056
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21178 10704 21234 10713
rect 21178 10639 21234 10648
rect 21192 10606 21220 10639
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21192 9926 21220 10542
rect 21284 10198 21312 10746
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 21376 9382 21404 11290
rect 21468 10742 21496 11834
rect 21560 11506 21588 13654
rect 21652 12102 21680 20402
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21744 16522 21772 16662
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21560 11478 21680 11506
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21454 9344 21510 9353
rect 21454 9279 21510 9288
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21192 9081 21220 9114
rect 21178 9072 21234 9081
rect 21178 9007 21234 9016
rect 21468 8974 21496 9279
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21362 8800 21418 8809
rect 21100 8430 21128 8774
rect 21362 8735 21418 8744
rect 21376 8430 21404 8735
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20732 7954 20852 7970
rect 20732 7948 20864 7954
rect 20732 7942 20812 7948
rect 20812 7890 20864 7896
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20626 6896 20682 6905
rect 20626 6831 20682 6840
rect 20732 6780 20760 7142
rect 20640 6752 20760 6780
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20036 3420 20116 3448
rect 19984 3402 20036 3408
rect 19260 2638 19380 2666
rect 19444 2650 19472 3402
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19904 2689 19932 3130
rect 19890 2680 19946 2689
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 18880 1828 18932 1834
rect 18880 1770 18932 1776
rect 18420 1760 18472 1766
rect 18420 1702 18472 1708
rect 19352 800 19380 2638
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19524 2644 19576 2650
rect 19890 2615 19946 2624
rect 19524 2586 19576 2592
rect 19536 2310 19564 2586
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19984 1692 20036 1698
rect 19984 1634 20036 1640
rect 19996 800 20024 1634
rect 20456 1358 20484 3878
rect 20640 3641 20668 6752
rect 20824 6304 20852 7890
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21100 7585 21128 7754
rect 21192 7750 21220 8026
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21086 7576 21142 7585
rect 21192 7546 21220 7686
rect 21086 7511 21142 7520
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6662 20944 7142
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 21008 6497 21036 7414
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 20994 6488 21050 6497
rect 20994 6423 21050 6432
rect 20996 6316 21048 6322
rect 20824 6276 20996 6304
rect 20996 6258 21048 6264
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20732 5778 20760 6122
rect 21100 5953 21128 6870
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21192 6186 21220 6802
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21086 5944 21142 5953
rect 21086 5879 21142 5888
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 21100 5574 21128 5782
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 21100 5166 21128 5510
rect 21284 5234 21312 7482
rect 21560 6848 21588 11290
rect 21652 9518 21680 11478
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21640 8560 21692 8566
rect 21640 8502 21692 8508
rect 21652 7041 21680 8502
rect 21638 7032 21694 7041
rect 21638 6967 21694 6976
rect 21376 6820 21588 6848
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21192 4826 21220 5102
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21086 4584 21142 4593
rect 20996 4548 21048 4554
rect 21086 4519 21142 4528
rect 20996 4490 21048 4496
rect 21008 3738 21036 4490
rect 21100 4486 21128 4519
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 21284 3670 21312 5170
rect 21376 5137 21404 6820
rect 21744 6746 21772 12582
rect 21836 12345 21864 19722
rect 22112 18222 22140 27814
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22480 18834 22508 27066
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 23730 22692 24006
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22756 23186 22784 24754
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 22848 23730 22876 24550
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 23032 22778 23060 23462
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22756 21962 22784 22374
rect 22652 21956 22704 21962
rect 22652 21898 22704 21904
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22664 21690 22692 21898
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 23032 21554 23060 22714
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23308 21078 23336 22034
rect 23296 21072 23348 21078
rect 23296 21014 23348 21020
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22572 18698 22600 19110
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 23204 18692 23256 18698
rect 23204 18634 23256 18640
rect 22192 18352 22244 18358
rect 22192 18294 22244 18300
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22112 17746 22140 18158
rect 22204 17882 22232 18294
rect 23216 18086 23244 18634
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 23216 17610 23244 18022
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16522 22232 16934
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22296 16504 22324 16730
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22376 16516 22428 16522
rect 22296 16476 22376 16504
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22112 16250 22140 16390
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 14952 21968 14958
rect 21914 14920 21916 14929
rect 21968 14920 21970 14929
rect 21914 14855 21970 14864
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21928 13977 21956 14418
rect 22020 14278 22048 16050
rect 22190 15056 22246 15065
rect 22190 14991 22246 15000
rect 22204 14550 22232 14991
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22112 14006 22140 14486
rect 22100 14000 22152 14006
rect 21914 13968 21970 13977
rect 22100 13942 22152 13948
rect 21914 13903 21970 13912
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 21928 13326 21956 13670
rect 22112 13433 22140 13670
rect 22098 13424 22154 13433
rect 22098 13359 22154 13368
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22020 12434 22048 13126
rect 21928 12406 22048 12434
rect 21822 12336 21878 12345
rect 21822 12271 21878 12280
rect 21836 10538 21864 12271
rect 21928 10742 21956 12406
rect 22008 12368 22060 12374
rect 22008 12310 22060 12316
rect 22020 11354 22048 12310
rect 22112 11898 22140 13126
rect 22296 12730 22324 16476
rect 22376 16458 22428 16464
rect 22468 16516 22520 16522
rect 22468 16458 22520 16464
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22388 15638 22416 15846
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22480 15094 22508 16458
rect 22664 16114 22692 16526
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22756 15570 22784 17274
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22848 16182 22876 16390
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22940 15706 22968 16118
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 23032 14958 23060 15642
rect 23124 15638 23152 15982
rect 23112 15632 23164 15638
rect 23112 15574 23164 15580
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22376 14884 22428 14890
rect 22376 14826 22428 14832
rect 22388 12918 22416 14826
rect 22744 14816 22796 14822
rect 23216 14804 23244 17546
rect 23308 16250 23336 18158
rect 23400 17270 23428 24278
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22710 23520 22918
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 24044 22574 24072 31078
rect 24872 30258 24900 37266
rect 25792 37262 25820 39200
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 26332 37256 26384 37262
rect 26332 37198 26384 37204
rect 24952 30592 25004 30598
rect 24952 30534 25004 30540
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24964 23254 24992 30534
rect 25964 30048 26016 30054
rect 25964 29990 26016 29996
rect 24952 23248 25004 23254
rect 24952 23190 25004 23196
rect 24964 22574 24992 23190
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 24032 22568 24084 22574
rect 24032 22510 24084 22516
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24952 22568 25004 22574
rect 24952 22510 25004 22516
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23768 21554 23796 21830
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 20602 23888 21490
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24044 20874 24072 21286
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24032 20868 24084 20874
rect 24032 20810 24084 20816
rect 24136 20602 24164 20878
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23400 16250 23428 17206
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23308 14958 23336 16186
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23400 15502 23428 15914
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 22744 14758 22796 14764
rect 23032 14776 23244 14804
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22664 12782 22692 13262
rect 22652 12776 22704 12782
rect 22296 12702 22416 12730
rect 22652 12718 22704 12724
rect 22388 12306 22416 12702
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22098 11520 22154 11529
rect 22098 11455 22154 11464
rect 22112 11354 22140 11455
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 22020 10674 22048 11086
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 22020 10062 22048 10610
rect 22204 10305 22232 11698
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 11082 22324 11630
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22388 11121 22416 11494
rect 22374 11112 22430 11121
rect 22284 11076 22336 11082
rect 22756 11082 22784 14758
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 22848 13870 22876 14282
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22374 11047 22430 11056
rect 22744 11076 22796 11082
rect 22284 11018 22336 11024
rect 22190 10296 22246 10305
rect 22190 10231 22246 10240
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21822 9072 21878 9081
rect 21822 9007 21824 9016
rect 21876 9007 21878 9016
rect 21824 8978 21876 8984
rect 21822 8936 21878 8945
rect 21822 8871 21824 8880
rect 21876 8871 21878 8880
rect 21824 8842 21876 8848
rect 21560 6718 21772 6746
rect 21456 6656 21508 6662
rect 21560 6644 21588 6718
rect 21508 6616 21588 6644
rect 21456 6598 21508 6604
rect 21362 5128 21418 5137
rect 21362 5063 21418 5072
rect 21376 4146 21404 5063
rect 21468 5001 21496 6598
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21560 5574 21588 6394
rect 21836 6089 21864 8842
rect 21928 7274 21956 9930
rect 22020 9042 22048 9998
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 21916 7268 21968 7274
rect 21916 7210 21968 7216
rect 21822 6080 21878 6089
rect 21822 6015 21878 6024
rect 21928 5692 21956 7210
rect 22020 6118 22048 7278
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6662 22140 7142
rect 22282 6896 22338 6905
rect 22282 6831 22338 6840
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 22100 6656 22152 6662
rect 22204 6633 22232 6666
rect 22296 6662 22324 6831
rect 22284 6656 22336 6662
rect 22100 6598 22152 6604
rect 22190 6624 22246 6633
rect 22284 6598 22336 6604
rect 22190 6559 22246 6568
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22008 5704 22060 5710
rect 21928 5664 22008 5692
rect 22008 5646 22060 5652
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 22008 5568 22060 5574
rect 22112 5556 22140 6122
rect 22060 5528 22140 5556
rect 22008 5510 22060 5516
rect 22020 5234 22048 5510
rect 22098 5400 22154 5409
rect 22098 5335 22154 5344
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21454 4992 21510 5001
rect 22112 4978 22140 5335
rect 21454 4927 21510 4936
rect 22020 4950 22140 4978
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21272 3664 21324 3670
rect 20626 3632 20682 3641
rect 21272 3606 21324 3612
rect 20626 3567 20682 3576
rect 20640 3482 20668 3567
rect 21180 3528 21232 3534
rect 20640 3476 21180 3482
rect 20640 3470 21232 3476
rect 20640 3454 21220 3470
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21008 1834 21036 2926
rect 21376 2922 21404 3878
rect 21560 3369 21588 4558
rect 22020 4554 22048 4950
rect 22008 4548 22060 4554
rect 22008 4490 22060 4496
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22112 4214 22140 4422
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 21546 3360 21602 3369
rect 21546 3295 21602 3304
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21928 2922 21956 3062
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 20996 1828 21048 1834
rect 20996 1770 21048 1776
rect 21192 1426 21220 2586
rect 22204 2446 22232 6122
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22296 3913 22324 5238
rect 22388 3942 22416 11047
rect 22744 11018 22796 11024
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22664 10690 22692 10746
rect 22664 10662 22784 10690
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22558 9480 22614 9489
rect 22558 9415 22614 9424
rect 22572 9382 22600 9415
rect 22560 9376 22612 9382
rect 22560 9318 22612 9324
rect 22468 8900 22520 8906
rect 22468 8842 22520 8848
rect 22480 6322 22508 8842
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22664 5522 22692 9658
rect 22756 7954 22784 10662
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 22848 7886 22876 13262
rect 22928 12708 22980 12714
rect 22928 12650 22980 12656
rect 22940 12238 22968 12650
rect 23032 12306 23060 14776
rect 23112 14000 23164 14006
rect 23112 13942 23164 13948
rect 23124 13734 23152 13942
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 23308 13546 23336 14894
rect 23386 14512 23442 14521
rect 23492 14482 23520 19450
rect 23768 18766 23796 19654
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23768 18290 23796 18566
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23386 14447 23442 14456
rect 23480 14476 23532 14482
rect 23400 14362 23428 14447
rect 23480 14418 23532 14424
rect 23400 14334 23520 14362
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23124 13518 23336 13546
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22940 10606 22968 12174
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11830 23060 12038
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23124 11694 23152 13518
rect 23400 13326 23428 13806
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23400 12850 23428 13262
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23112 11688 23164 11694
rect 23112 11630 23164 11636
rect 23110 11520 23166 11529
rect 23110 11455 23166 11464
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 23124 10130 23152 11455
rect 23216 10198 23244 12174
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23308 9738 23336 12174
rect 23400 11898 23428 12786
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23492 11778 23520 14334
rect 23400 11750 23520 11778
rect 23400 11370 23428 11750
rect 23480 11552 23532 11558
rect 23478 11520 23480 11529
rect 23532 11520 23534 11529
rect 23478 11455 23534 11464
rect 23400 11342 23520 11370
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23400 10130 23428 10474
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23032 9710 23336 9738
rect 23032 8430 23060 9710
rect 23492 9674 23520 11342
rect 23584 10606 23612 15098
rect 23676 10996 23704 15506
rect 23848 15496 23900 15502
rect 23846 15464 23848 15473
rect 23900 15464 23902 15473
rect 23846 15399 23902 15408
rect 23860 14940 23888 15399
rect 23940 15360 23992 15366
rect 23938 15328 23940 15337
rect 24032 15360 24084 15366
rect 23992 15328 23994 15337
rect 24032 15302 24084 15308
rect 23938 15263 23994 15272
rect 24044 15094 24072 15302
rect 24032 15088 24084 15094
rect 24032 15030 24084 15036
rect 23860 14912 23980 14940
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 12442 23796 13262
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23756 11008 23808 11014
rect 23676 10968 23756 10996
rect 23756 10950 23808 10956
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23400 9646 23520 9674
rect 23400 9586 23428 9646
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23112 9376 23164 9382
rect 23112 9318 23164 9324
rect 23124 8498 23152 9318
rect 23386 8664 23442 8673
rect 23204 8628 23256 8634
rect 23386 8599 23442 8608
rect 23204 8570 23256 8576
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22756 5914 22784 7686
rect 23020 6384 23072 6390
rect 23020 6326 23072 6332
rect 23032 6186 23060 6326
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 23018 6080 23074 6089
rect 23018 6015 23074 6024
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 22572 5494 22692 5522
rect 22572 5409 22600 5494
rect 22558 5400 22614 5409
rect 22558 5335 22614 5344
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22664 5001 22692 5306
rect 22650 4992 22706 5001
rect 22650 4927 22706 4936
rect 23032 4078 23060 6015
rect 23216 5370 23244 8570
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 23294 4448 23350 4457
rect 23294 4383 23350 4392
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 22652 4004 22704 4010
rect 22652 3946 22704 3952
rect 22376 3936 22428 3942
rect 22282 3904 22338 3913
rect 22376 3878 22428 3884
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22282 3839 22338 3848
rect 22376 2984 22428 2990
rect 22374 2952 22376 2961
rect 22428 2952 22430 2961
rect 22374 2887 22430 2896
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22468 2372 22520 2378
rect 22468 2314 22520 2320
rect 22480 2106 22508 2314
rect 22468 2100 22520 2106
rect 22468 2042 22520 2048
rect 21272 1556 21324 1562
rect 21272 1498 21324 1504
rect 21180 1420 21232 1426
rect 21180 1362 21232 1368
rect 20444 1352 20496 1358
rect 20444 1294 20496 1300
rect 21284 800 21312 1498
rect 22572 800 22600 3878
rect 22664 2990 22692 3946
rect 23308 3466 23336 4383
rect 23400 4078 23428 8599
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23492 7342 23520 8298
rect 23480 7336 23532 7342
rect 23480 7278 23532 7284
rect 23492 6934 23520 7278
rect 23480 6928 23532 6934
rect 23480 6870 23532 6876
rect 23584 6254 23612 10542
rect 23768 10266 23796 10950
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23756 9988 23808 9994
rect 23860 9976 23888 10950
rect 23808 9948 23888 9976
rect 23756 9930 23808 9936
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23676 8566 23704 9862
rect 23952 9674 23980 14912
rect 24030 13560 24086 13569
rect 24030 13495 24086 13504
rect 23860 9646 23980 9674
rect 23756 9104 23808 9110
rect 23754 9072 23756 9081
rect 23808 9072 23810 9081
rect 23754 9007 23810 9016
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23768 5681 23796 7346
rect 23860 5953 23888 9646
rect 24044 8430 24072 13495
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 24044 7342 24072 7414
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24136 7274 24164 15846
rect 24228 14929 24256 17070
rect 24214 14920 24270 14929
rect 24214 14855 24270 14864
rect 24228 12986 24256 14855
rect 24320 14113 24348 22510
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24596 21146 24624 21966
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24584 21140 24636 21146
rect 24584 21082 24636 21088
rect 24688 21010 24716 21286
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 24780 20466 24808 20878
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24504 16182 24532 16390
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24412 15706 24440 15982
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24596 14770 24624 17138
rect 24688 17105 24716 18770
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24780 17218 24808 18702
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24872 18358 24900 18566
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24872 17746 24900 18158
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 25056 17338 25084 22646
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25516 21146 25544 21490
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 25516 17270 25544 18566
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25504 17264 25556 17270
rect 24780 17190 24900 17218
rect 25504 17206 25556 17212
rect 24872 17134 24900 17190
rect 24860 17128 24912 17134
rect 24674 17096 24730 17105
rect 24860 17070 24912 17076
rect 24674 17031 24730 17040
rect 24872 15502 24900 17070
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24860 15496 24912 15502
rect 24860 15438 24912 15444
rect 24780 15094 24808 15438
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24504 14742 24624 14770
rect 24306 14104 24362 14113
rect 24306 14039 24362 14048
rect 24320 13870 24348 14039
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24308 13728 24360 13734
rect 24308 13670 24360 13676
rect 24320 13258 24348 13670
rect 24308 13252 24360 13258
rect 24308 13194 24360 13200
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12646 24348 12786
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24228 11257 24256 12582
rect 24412 12434 24440 13806
rect 24320 12406 24440 12434
rect 24214 11248 24270 11257
rect 24214 11183 24270 11192
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24228 7954 24256 9522
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24228 7478 24256 7754
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 23846 5944 23902 5953
rect 23846 5879 23902 5888
rect 23860 5710 23888 5879
rect 23848 5704 23900 5710
rect 23754 5672 23810 5681
rect 23848 5646 23900 5652
rect 23754 5607 23810 5616
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23480 5092 23532 5098
rect 23480 5034 23532 5040
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23296 3460 23348 3466
rect 23296 3402 23348 3408
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22664 2514 22692 2926
rect 23492 2650 23520 5034
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4758 23612 4966
rect 23572 4752 23624 4758
rect 23572 4694 23624 4700
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23204 1624 23256 1630
rect 23204 1566 23256 1572
rect 23216 800 23244 1566
rect 23308 1562 23336 2382
rect 23676 1970 23704 5510
rect 23756 5024 23808 5030
rect 23754 4992 23756 5001
rect 23808 4992 23810 5001
rect 23754 4927 23810 4936
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 23860 3602 23888 4422
rect 23952 4078 23980 7210
rect 24320 5778 24348 12406
rect 24398 11928 24454 11937
rect 24398 11863 24454 11872
rect 24412 11762 24440 11863
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24504 11336 24532 14742
rect 24584 13796 24636 13802
rect 24584 13738 24636 13744
rect 24412 11308 24532 11336
rect 24412 10062 24440 11308
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24412 8090 24440 9998
rect 24596 9897 24624 13738
rect 24688 11626 24716 14894
rect 24872 13297 24900 15438
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25044 13524 25096 13530
rect 25044 13466 25096 13472
rect 24858 13288 24914 13297
rect 24858 13223 24914 13232
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24676 11620 24728 11626
rect 24676 11562 24728 11568
rect 24676 11348 24728 11354
rect 24676 11290 24728 11296
rect 24582 9888 24638 9897
rect 24582 9823 24638 9832
rect 24688 9674 24716 11290
rect 24596 9646 24716 9674
rect 24780 9654 24808 12922
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9654 24900 9862
rect 24768 9648 24820 9654
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24504 8974 24532 9318
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24490 7848 24546 7857
rect 24490 7783 24546 7792
rect 24504 6322 24532 7783
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24308 5772 24360 5778
rect 24308 5714 24360 5720
rect 24398 5672 24454 5681
rect 24398 5607 24454 5616
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24044 4554 24072 4966
rect 24032 4548 24084 4554
rect 24032 4490 24084 4496
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23952 3602 23980 3878
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 23938 3224 23994 3233
rect 23938 3159 23994 3168
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23860 2650 23888 2994
rect 23952 2922 23980 3159
rect 24320 2922 24348 3334
rect 24412 3097 24440 5607
rect 24504 5234 24532 6258
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24490 3768 24546 3777
rect 24490 3703 24546 3712
rect 24504 3534 24532 3703
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 24398 3088 24454 3097
rect 24596 3058 24624 9646
rect 24768 9590 24820 9596
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24780 9178 24808 9454
rect 24964 9450 24992 12174
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24688 8974 24716 9114
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24860 8424 24912 8430
rect 24766 8392 24822 8401
rect 24860 8366 24912 8372
rect 24766 8327 24822 8336
rect 24780 8022 24808 8327
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24780 6730 24808 7647
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24688 5914 24716 6666
rect 24780 6497 24808 6666
rect 24766 6488 24822 6497
rect 24766 6423 24822 6432
rect 24872 6322 24900 8366
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24964 7546 24992 7754
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25056 7274 25084 13466
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 25042 6896 25098 6905
rect 25042 6831 25098 6840
rect 24950 6624 25006 6633
rect 24950 6559 25006 6568
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24860 6180 24912 6186
rect 24860 6122 24912 6128
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24780 5642 24808 6054
rect 24872 5778 24900 6122
rect 24964 5778 24992 6559
rect 25056 6322 25084 6831
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24674 5400 24730 5409
rect 24674 5335 24730 5344
rect 24688 4554 24716 5335
rect 24676 4548 24728 4554
rect 24676 4490 24728 4496
rect 24766 4312 24822 4321
rect 24766 4247 24822 4256
rect 24674 3632 24730 3641
rect 24674 3567 24730 3576
rect 24398 3023 24454 3032
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 23940 2916 23992 2922
rect 23940 2858 23992 2864
rect 24308 2916 24360 2922
rect 24308 2858 24360 2864
rect 24688 2774 24716 3567
rect 24780 3466 24808 4247
rect 24872 4010 24900 5714
rect 25044 5296 25096 5302
rect 25044 5238 25096 5244
rect 25056 5137 25084 5238
rect 25042 5128 25098 5137
rect 25042 5063 25098 5072
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24964 3754 24992 4082
rect 24872 3726 24992 3754
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24872 3369 24900 3726
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 24858 3360 24914 3369
rect 24858 3295 24914 3304
rect 24504 2746 24716 2774
rect 24964 2774 24992 3606
rect 25056 2922 25084 4082
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 24964 2746 25084 2774
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 23296 1556 23348 1562
rect 23296 1498 23348 1504
rect 24504 800 24532 2746
rect 25056 2689 25084 2746
rect 24858 2680 24914 2689
rect 24858 2615 24860 2624
rect 24912 2615 24914 2624
rect 25042 2680 25098 2689
rect 25042 2615 25098 2624
rect 24860 2586 24912 2592
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24780 2038 24808 2382
rect 24768 2032 24820 2038
rect 24768 1974 24820 1980
rect 25148 1426 25176 11698
rect 25240 11665 25268 14350
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25332 14006 25360 14214
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25226 11656 25282 11665
rect 25226 11591 25282 11600
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25240 9722 25268 9998
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25240 8566 25268 8774
rect 25332 8673 25360 12922
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25424 11150 25452 11834
rect 25608 11354 25636 14350
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 12986 25728 13194
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25424 8974 25452 9522
rect 25700 9217 25728 11698
rect 25686 9208 25742 9217
rect 25686 9143 25742 9152
rect 25792 9110 25820 17614
rect 25976 17270 26004 29990
rect 26344 29646 26372 37198
rect 26436 37126 26464 39200
rect 27724 37330 27752 39200
rect 27712 37324 27764 37330
rect 27712 37266 27764 37272
rect 29012 37262 29040 39200
rect 29656 37330 29684 39200
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 28080 37256 28132 37262
rect 28080 37198 28132 37204
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26528 22710 26556 31622
rect 27172 30258 27200 37062
rect 28092 36854 28120 37198
rect 30944 37126 30972 39200
rect 31024 37256 31076 37262
rect 31024 37198 31076 37204
rect 32128 37256 32180 37262
rect 32128 37198 32180 37204
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 28080 36848 28132 36854
rect 28080 36790 28132 36796
rect 27160 30252 27212 30258
rect 27160 30194 27212 30200
rect 27712 28960 27764 28966
rect 27712 28902 27764 28908
rect 27068 25900 27120 25906
rect 27068 25842 27120 25848
rect 26516 22704 26568 22710
rect 26516 22646 26568 22652
rect 27080 21486 27108 25842
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27540 21622 27568 21830
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 26240 19984 26292 19990
rect 26240 19926 26292 19932
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26068 17882 26096 18294
rect 26160 18222 26188 19654
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 26056 17264 26108 17270
rect 26056 17206 26108 17212
rect 26068 16794 26096 17206
rect 26056 16788 26108 16794
rect 26056 16730 26108 16736
rect 26056 16176 26108 16182
rect 26056 16118 26108 16124
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25976 14385 26004 15846
rect 26068 14618 26096 16118
rect 26160 16046 26188 18158
rect 26252 18086 26280 19926
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 26516 18896 26568 18902
rect 26516 18838 26568 18844
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26252 17746 26280 18022
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26344 17610 26372 18566
rect 26332 17604 26384 17610
rect 26332 17546 26384 17552
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26252 14618 26280 15098
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 25962 14376 26018 14385
rect 25962 14311 26018 14320
rect 25976 13818 26004 14311
rect 25976 13790 26096 13818
rect 25962 13696 26018 13705
rect 25962 13631 26018 13640
rect 25976 13394 26004 13631
rect 25872 13388 25924 13394
rect 25872 13330 25924 13336
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25884 9586 25912 13330
rect 26068 12434 26096 13790
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 25976 12406 26096 12434
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 25872 9104 25924 9110
rect 25872 9046 25924 9052
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25318 8664 25374 8673
rect 25318 8599 25374 8608
rect 25332 8566 25360 8599
rect 25228 8560 25280 8566
rect 25228 8502 25280 8508
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25320 6928 25372 6934
rect 25320 6870 25372 6876
rect 25424 6882 25452 8910
rect 25884 8106 25912 9046
rect 25976 8430 26004 12406
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26160 9110 26188 11630
rect 26344 11626 26372 13194
rect 26332 11620 26384 11626
rect 26332 11562 26384 11568
rect 26148 9104 26200 9110
rect 26148 9046 26200 9052
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26148 8900 26200 8906
rect 26148 8842 26200 8848
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 26054 8528 26110 8537
rect 26054 8463 26056 8472
rect 26108 8463 26110 8472
rect 26056 8434 26108 8440
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 25884 8078 26004 8106
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25332 5030 25360 6870
rect 25424 6854 25636 6882
rect 25410 6488 25466 6497
rect 25410 6423 25466 6432
rect 25424 5710 25452 6423
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 25424 4622 25452 5646
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25320 4004 25372 4010
rect 25320 3946 25372 3952
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 25240 1494 25268 3878
rect 25332 3126 25360 3946
rect 25410 3496 25466 3505
rect 25410 3431 25466 3440
rect 25320 3120 25372 3126
rect 25320 3062 25372 3068
rect 25424 2774 25452 3431
rect 25516 3233 25544 5170
rect 25608 4146 25636 6854
rect 25792 6186 25820 7890
rect 25870 7576 25926 7585
rect 25870 7511 25926 7520
rect 25884 6322 25912 7511
rect 25976 6730 26004 8078
rect 26160 7954 26188 8842
rect 26148 7948 26200 7954
rect 26148 7890 26200 7896
rect 26148 7812 26200 7818
rect 26148 7754 26200 7760
rect 26160 7426 26188 7754
rect 26252 7546 26280 8842
rect 26332 8084 26384 8090
rect 26332 8026 26384 8032
rect 26344 7750 26372 8026
rect 26332 7744 26384 7750
rect 26332 7686 26384 7692
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 26160 7398 26280 7426
rect 26252 7342 26280 7398
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26148 7268 26200 7274
rect 26148 7210 26200 7216
rect 26160 6798 26188 7210
rect 26330 7032 26386 7041
rect 26330 6967 26386 6976
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 25964 6724 26016 6730
rect 25964 6666 26016 6672
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 25780 6180 25832 6186
rect 25780 6122 25832 6128
rect 25686 5944 25742 5953
rect 25686 5879 25742 5888
rect 25700 5710 25728 5879
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25700 4622 25728 5646
rect 25688 4616 25740 4622
rect 25688 4558 25740 4564
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 25608 4049 25636 4082
rect 25594 4040 25650 4049
rect 25594 3975 25650 3984
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25596 3392 25648 3398
rect 25596 3334 25648 3340
rect 25502 3224 25558 3233
rect 25502 3159 25558 3168
rect 25608 3126 25636 3334
rect 25700 3126 25728 3606
rect 25976 3505 26004 6666
rect 26054 6488 26110 6497
rect 26054 6423 26110 6432
rect 25962 3496 26018 3505
rect 25962 3431 25964 3440
rect 26016 3431 26018 3440
rect 25964 3402 26016 3408
rect 25976 3371 26004 3402
rect 26068 3346 26096 6423
rect 26160 6254 26188 6734
rect 26148 6248 26200 6254
rect 26148 6190 26200 6196
rect 26160 5556 26188 6190
rect 26344 5778 26372 6967
rect 26436 6322 26464 8978
rect 26528 6338 26556 18838
rect 26700 18692 26752 18698
rect 26700 18634 26752 18640
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26620 17134 26648 18158
rect 26608 17128 26660 17134
rect 26608 17070 26660 17076
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26620 8430 26648 14554
rect 26712 10810 26740 18634
rect 27264 18358 27292 19722
rect 27540 18834 27568 20266
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 27252 18352 27304 18358
rect 27252 18294 27304 18300
rect 27160 17604 27212 17610
rect 27160 17546 27212 17552
rect 27068 17128 27120 17134
rect 27068 17070 27120 17076
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26804 11898 26832 12854
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26608 8424 26660 8430
rect 26608 8366 26660 8372
rect 26804 7478 26832 11086
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26698 7304 26754 7313
rect 26896 7290 26924 12174
rect 26974 11928 27030 11937
rect 26974 11863 27030 11872
rect 26754 7262 26924 7290
rect 26698 7239 26754 7248
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26620 6458 26648 6598
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26424 6316 26476 6322
rect 26528 6310 26648 6338
rect 26424 6258 26476 6264
rect 26424 6180 26476 6186
rect 26424 6122 26476 6128
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26160 5528 26372 5556
rect 26148 5160 26200 5166
rect 26148 5102 26200 5108
rect 26160 4622 26188 5102
rect 26344 4865 26372 5528
rect 26436 5234 26464 6122
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26330 4856 26386 4865
rect 26330 4791 26386 4800
rect 26148 4616 26200 4622
rect 26148 4558 26200 4564
rect 26148 4480 26200 4486
rect 26240 4480 26292 4486
rect 26148 4422 26200 4428
rect 26238 4448 26240 4457
rect 26292 4448 26294 4457
rect 26160 4282 26188 4422
rect 26238 4383 26294 4392
rect 26148 4276 26200 4282
rect 26148 4218 26200 4224
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26252 4162 26280 4218
rect 26160 4134 26280 4162
rect 26160 3534 26188 4134
rect 26344 3618 26372 4791
rect 26528 4554 26556 6054
rect 26620 5370 26648 6310
rect 26712 6254 26740 7239
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26790 5944 26846 5953
rect 26790 5879 26846 5888
rect 26804 5710 26832 5879
rect 26988 5794 27016 11863
rect 27080 7721 27108 17070
rect 27172 16590 27200 17546
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 16250 27292 16390
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27632 15162 27660 21558
rect 27724 21078 27752 28902
rect 28092 28082 28120 36790
rect 28448 36780 28500 36786
rect 28448 36722 28500 36728
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28000 22098 28028 25230
rect 28368 23866 28396 32846
rect 28460 27062 28488 36722
rect 29840 31346 29868 37062
rect 31036 36922 31064 37198
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 29828 30592 29880 30598
rect 29828 30534 29880 30540
rect 29840 27130 29868 30534
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 29184 26376 29236 26382
rect 29184 26318 29236 26324
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 29196 22778 29224 26318
rect 30748 24404 30800 24410
rect 30748 24346 30800 24352
rect 30760 23866 30788 24346
rect 30748 23860 30800 23866
rect 30748 23802 30800 23808
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 29184 22772 29236 22778
rect 29184 22714 29236 22720
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 27988 22092 28040 22098
rect 27988 22034 28040 22040
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27816 19854 27844 20810
rect 28724 20256 28776 20262
rect 28724 20198 28776 20204
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 28632 19780 28684 19786
rect 28632 19722 28684 19728
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 27724 17678 27752 18566
rect 28368 18290 28396 18566
rect 28552 18290 28580 19110
rect 28356 18284 28408 18290
rect 28356 18226 28408 18232
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27816 16182 27844 18090
rect 27896 17536 27948 17542
rect 27896 17478 27948 17484
rect 27908 17270 27936 17478
rect 27896 17264 27948 17270
rect 27896 17206 27948 17212
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27816 15178 27844 16118
rect 27620 15156 27672 15162
rect 27816 15150 27936 15178
rect 27620 15098 27672 15104
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27264 14414 27292 14758
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27724 14414 27752 14554
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27712 14408 27764 14414
rect 27712 14350 27764 14356
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 27356 14226 27384 14282
rect 27264 14198 27384 14226
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27158 13968 27214 13977
rect 27158 13903 27214 13912
rect 27172 13258 27200 13903
rect 27264 13870 27292 14198
rect 27724 14006 27752 14214
rect 27344 14000 27396 14006
rect 27344 13942 27396 13948
rect 27712 14000 27764 14006
rect 27712 13942 27764 13948
rect 27252 13864 27304 13870
rect 27252 13806 27304 13812
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 27172 8514 27200 13194
rect 27264 11830 27292 13806
rect 27356 12442 27384 13942
rect 27908 13938 27936 15150
rect 28264 15020 28316 15026
rect 28264 14962 28316 14968
rect 28172 14272 28224 14278
rect 28172 14214 28224 14220
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27988 13456 28040 13462
rect 27988 13398 28040 13404
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27344 12436 27396 12442
rect 27344 12378 27396 12384
rect 27252 11824 27304 11830
rect 27252 11766 27304 11772
rect 27344 11824 27396 11830
rect 27344 11766 27396 11772
rect 27434 11792 27490 11801
rect 27356 11354 27384 11766
rect 27434 11727 27490 11736
rect 27448 11694 27476 11727
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 27448 9654 27476 9862
rect 27436 9648 27488 9654
rect 27436 9590 27488 9596
rect 27172 8486 27292 8514
rect 27066 7712 27122 7721
rect 27066 7647 27122 7656
rect 27158 7440 27214 7449
rect 27158 7375 27160 7384
rect 27212 7375 27214 7384
rect 27160 7346 27212 7352
rect 27264 7342 27292 8486
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 27264 6458 27292 6938
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 26896 5766 27016 5794
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26516 4548 26568 4554
rect 26516 4490 26568 4496
rect 26516 3936 26568 3942
rect 26516 3878 26568 3884
rect 26344 3590 26464 3618
rect 26436 3534 26464 3590
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26148 3392 26200 3398
rect 26068 3340 26148 3346
rect 26068 3334 26200 3340
rect 26068 3318 26188 3334
rect 26344 3233 26372 3470
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26330 3224 26386 3233
rect 26436 3194 26464 3334
rect 26330 3159 26386 3168
rect 26424 3188 26476 3194
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 25688 3120 25740 3126
rect 25688 3062 25740 3068
rect 25872 2984 25924 2990
rect 25872 2926 25924 2932
rect 25332 2746 25452 2774
rect 25332 2281 25360 2746
rect 25884 2446 25912 2926
rect 26344 2650 26372 3159
rect 26424 3130 26476 3136
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26160 2310 26188 2382
rect 25780 2304 25832 2310
rect 25318 2272 25374 2281
rect 25780 2246 25832 2252
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 25318 2207 25374 2216
rect 25228 1488 25280 1494
rect 25228 1430 25280 1436
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 25792 800 25820 2246
rect 26528 1737 26556 3878
rect 26620 3126 26648 5306
rect 26896 4622 26924 5766
rect 27264 5545 27292 6258
rect 27540 5778 27568 12582
rect 27632 12306 27660 12718
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27632 8090 27660 11630
rect 27802 11112 27858 11121
rect 27802 11047 27858 11056
rect 27620 8084 27672 8090
rect 27620 8026 27672 8032
rect 27620 7812 27672 7818
rect 27620 7754 27672 7760
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 27344 5636 27396 5642
rect 27344 5578 27396 5584
rect 27250 5536 27306 5545
rect 27250 5471 27306 5480
rect 26884 4616 26936 4622
rect 26884 4558 26936 4564
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26804 4214 26832 4422
rect 26792 4208 26844 4214
rect 26792 4150 26844 4156
rect 26896 4026 26924 4422
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 26712 3998 26924 4026
rect 26608 3120 26660 3126
rect 26608 3062 26660 3068
rect 26712 2825 26740 3998
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26698 2816 26754 2825
rect 26698 2751 26754 2760
rect 26804 2106 26832 3878
rect 26884 3528 26936 3534
rect 26882 3496 26884 3505
rect 26936 3496 26938 3505
rect 26882 3431 26938 3440
rect 27066 2816 27122 2825
rect 27066 2751 27122 2760
rect 26792 2100 26844 2106
rect 26792 2042 26844 2048
rect 26514 1728 26570 1737
rect 26514 1663 26570 1672
rect 27080 800 27108 2751
rect 27172 1086 27200 4082
rect 27250 3224 27306 3233
rect 27250 3159 27306 3168
rect 27264 2990 27292 3159
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 27356 2774 27384 5578
rect 27540 4842 27568 5714
rect 27448 4814 27568 4842
rect 27448 4214 27476 4814
rect 27528 4752 27580 4758
rect 27528 4694 27580 4700
rect 27540 4554 27568 4694
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27436 4208 27488 4214
rect 27436 4150 27488 4156
rect 27632 3942 27660 7754
rect 27816 6866 27844 11047
rect 28000 9518 28028 13398
rect 28184 13258 28212 14214
rect 28080 13252 28132 13258
rect 28080 13194 28132 13200
rect 28172 13252 28224 13258
rect 28172 13194 28224 13200
rect 28092 10606 28120 13194
rect 28276 12238 28304 14962
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 14414 28396 14894
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 28276 11898 28304 12174
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28080 10600 28132 10606
rect 28080 10542 28132 10548
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28448 10532 28500 10538
rect 28448 10474 28500 10480
rect 28460 10198 28488 10474
rect 28448 10192 28500 10198
rect 28448 10134 28500 10140
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 27988 9512 28040 9518
rect 27988 9454 28040 9460
rect 28000 9110 28028 9454
rect 27988 9104 28040 9110
rect 27988 9046 28040 9052
rect 28368 8634 28396 9590
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28460 8514 28488 10134
rect 28552 8634 28580 10542
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28356 8492 28408 8498
rect 28460 8486 28580 8514
rect 28356 8434 28408 8440
rect 28368 8294 28396 8434
rect 28448 8356 28500 8362
rect 28448 8298 28500 8304
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 27816 6662 27844 6802
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27908 6458 27936 7686
rect 28460 6798 28488 8298
rect 28552 7954 28580 8486
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 27896 6452 27948 6458
rect 27896 6394 27948 6400
rect 28264 5772 28316 5778
rect 28264 5714 28316 5720
rect 27804 5704 27856 5710
rect 27802 5672 27804 5681
rect 27988 5704 28040 5710
rect 27856 5672 27858 5681
rect 27988 5646 28040 5652
rect 27802 5607 27858 5616
rect 28000 4622 28028 5646
rect 28276 5302 28304 5714
rect 28264 5296 28316 5302
rect 28264 5238 28316 5244
rect 28460 5166 28488 6734
rect 28540 5636 28592 5642
rect 28540 5578 28592 5584
rect 28552 5302 28580 5578
rect 28540 5296 28592 5302
rect 28540 5238 28592 5244
rect 28448 5160 28500 5166
rect 28448 5102 28500 5108
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 27816 4298 27844 4558
rect 28264 4548 28316 4554
rect 28264 4490 28316 4496
rect 28080 4480 28132 4486
rect 28080 4422 28132 4428
rect 27816 4270 28028 4298
rect 28000 4146 28028 4270
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 27988 4140 28040 4146
rect 27988 4082 28040 4088
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 3369 27660 3878
rect 27618 3360 27674 3369
rect 27618 3295 27674 3304
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27264 2746 27384 2774
rect 27264 2417 27292 2746
rect 27344 2440 27396 2446
rect 27250 2408 27306 2417
rect 27344 2382 27396 2388
rect 27250 2343 27306 2352
rect 27356 1698 27384 2382
rect 27344 1692 27396 1698
rect 27344 1634 27396 1640
rect 27448 1630 27476 3062
rect 27632 2922 27660 3295
rect 27620 2916 27672 2922
rect 27620 2858 27672 2864
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27436 1624 27488 1630
rect 27436 1566 27488 1572
rect 27160 1080 27212 1086
rect 27160 1022 27212 1028
rect 27724 800 27752 2382
rect 27816 1766 27844 4082
rect 27896 2916 27948 2922
rect 27896 2858 27948 2864
rect 27908 2514 27936 2858
rect 27896 2508 27948 2514
rect 27896 2450 27948 2456
rect 28092 1873 28120 4422
rect 28276 3534 28304 4490
rect 28552 4214 28580 4558
rect 28540 4208 28592 4214
rect 28540 4150 28592 4156
rect 28356 4072 28408 4078
rect 28552 4026 28580 4150
rect 28356 4014 28408 4020
rect 28368 3942 28396 4014
rect 28460 3998 28580 4026
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 28460 3534 28488 3998
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 28552 3738 28580 3878
rect 28540 3732 28592 3738
rect 28540 3674 28592 3680
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 28264 3528 28316 3534
rect 28264 3470 28316 3476
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28172 3392 28224 3398
rect 28172 3334 28224 3340
rect 28184 2854 28212 3334
rect 28552 3058 28580 3538
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28644 2514 28672 19722
rect 28736 19378 28764 20198
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17066 29040 18022
rect 29104 17746 29132 22578
rect 29460 21344 29512 21350
rect 29460 21286 29512 21292
rect 29184 20460 29236 20466
rect 29184 20402 29236 20408
rect 29196 19854 29224 20402
rect 29184 19848 29236 19854
rect 29184 19790 29236 19796
rect 29092 17740 29144 17746
rect 29092 17682 29144 17688
rect 29104 17270 29132 17682
rect 29196 17678 29224 19790
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29276 17536 29328 17542
rect 29276 17478 29328 17484
rect 29092 17264 29144 17270
rect 29092 17206 29144 17212
rect 29288 17202 29316 17478
rect 29276 17196 29328 17202
rect 29276 17138 29328 17144
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29012 15502 29040 15846
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 29368 14544 29420 14550
rect 29368 14486 29420 14492
rect 29380 13870 29408 14486
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29380 12986 29408 13806
rect 29472 13190 29500 21286
rect 30116 19378 30144 23666
rect 30840 21480 30892 21486
rect 30840 21422 30892 21428
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29644 15972 29696 15978
rect 29644 15914 29696 15920
rect 29656 13870 29684 15914
rect 29840 15570 29868 17070
rect 29828 15564 29880 15570
rect 29828 15506 29880 15512
rect 29920 15428 29972 15434
rect 29920 15370 29972 15376
rect 29932 14074 29960 15370
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 30024 14482 30052 14894
rect 30012 14476 30064 14482
rect 30012 14418 30064 14424
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 29644 13864 29696 13870
rect 29644 13806 29696 13812
rect 29460 13184 29512 13190
rect 29460 13126 29512 13132
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 28828 12434 28856 12718
rect 29012 12442 29040 12718
rect 28736 12406 28856 12434
rect 29000 12436 29052 12442
rect 28736 4570 28764 12406
rect 29000 12378 29052 12384
rect 29276 11144 29328 11150
rect 29276 11086 29328 11092
rect 29184 9988 29236 9994
rect 29184 9930 29236 9936
rect 28816 9648 28868 9654
rect 28814 9616 28816 9625
rect 28868 9616 28870 9625
rect 28814 9551 28870 9560
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 28814 7168 28870 7177
rect 28814 7103 28870 7112
rect 28828 5302 28856 7103
rect 29104 6798 29132 8434
rect 29092 6792 29144 6798
rect 28998 6760 29054 6769
rect 29092 6734 29144 6740
rect 28998 6695 29054 6704
rect 28908 6384 28960 6390
rect 28906 6352 28908 6361
rect 28960 6352 28962 6361
rect 28906 6287 28962 6296
rect 29012 5914 29040 6695
rect 29196 6458 29224 9930
rect 29288 9450 29316 11086
rect 29656 9586 29684 13806
rect 29828 12164 29880 12170
rect 29828 12106 29880 12112
rect 29840 9994 29868 12106
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 29826 9888 29882 9897
rect 29826 9823 29882 9832
rect 29644 9580 29696 9586
rect 29644 9522 29696 9528
rect 29276 9444 29328 9450
rect 29276 9386 29328 9392
rect 29288 7954 29316 9386
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29092 6180 29144 6186
rect 29092 6122 29144 6128
rect 29000 5908 29052 5914
rect 29000 5850 29052 5856
rect 29104 5710 29132 6122
rect 29288 5778 29316 7890
rect 29840 6458 29868 9823
rect 29932 9722 29960 9930
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30024 9722 30052 9862
rect 29920 9716 29972 9722
rect 29920 9658 29972 9664
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 29920 9376 29972 9382
rect 29920 9318 29972 9324
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 29460 6316 29512 6322
rect 29460 6258 29512 6264
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 29092 5704 29144 5710
rect 29092 5646 29144 5652
rect 28816 5296 28868 5302
rect 28816 5238 28868 5244
rect 28814 5128 28870 5137
rect 28814 5063 28870 5072
rect 28828 5030 28856 5063
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28920 4622 28948 5646
rect 29000 5092 29052 5098
rect 29000 5034 29052 5040
rect 28908 4616 28960 4622
rect 28736 4542 28856 4570
rect 28908 4558 28960 4564
rect 28828 3777 28856 4542
rect 29012 4282 29040 5034
rect 29276 4616 29328 4622
rect 29276 4558 29328 4564
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 29104 4146 29224 4162
rect 29288 4146 29316 4558
rect 29472 4282 29500 6258
rect 29932 5710 29960 9318
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29920 5704 29972 5710
rect 29920 5646 29972 5652
rect 29656 5234 29684 5646
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 29092 4140 29224 4146
rect 29144 4134 29224 4140
rect 29092 4082 29144 4088
rect 28920 4026 28948 4082
rect 28920 3998 29132 4026
rect 28814 3768 28870 3777
rect 28724 3732 28776 3738
rect 28814 3703 28870 3712
rect 28724 3674 28776 3680
rect 28736 3534 28764 3674
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28736 2854 28764 3470
rect 28828 3398 28856 3703
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28920 3097 28948 3538
rect 29104 3534 29132 3998
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29196 3346 29224 4134
rect 29276 4140 29328 4146
rect 29276 4082 29328 4088
rect 29276 4004 29328 4010
rect 29276 3946 29328 3952
rect 29288 3670 29316 3946
rect 29368 3936 29420 3942
rect 29368 3878 29420 3884
rect 29276 3664 29328 3670
rect 29276 3606 29328 3612
rect 29012 3318 29224 3346
rect 28906 3088 28962 3097
rect 28906 3023 28962 3032
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 29012 2689 29040 3318
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 28998 2680 29054 2689
rect 28998 2615 29054 2624
rect 28632 2508 28684 2514
rect 28632 2450 28684 2456
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 28078 1864 28134 1873
rect 28078 1799 28134 1808
rect 27804 1760 27856 1766
rect 27804 1702 27856 1708
rect 29012 800 29040 2382
rect 29104 1902 29132 2858
rect 29380 2774 29408 3878
rect 29288 2746 29408 2774
rect 29092 1896 29144 1902
rect 29092 1838 29144 1844
rect 29288 1222 29316 2746
rect 29564 2310 29592 5170
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29920 5024 29972 5030
rect 29920 4966 29972 4972
rect 29734 4856 29790 4865
rect 29734 4791 29790 4800
rect 29748 4622 29776 4791
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29656 3738 29684 4014
rect 29840 3738 29868 4966
rect 29932 4486 29960 4966
rect 29920 4480 29972 4486
rect 29920 4422 29972 4428
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 29736 2984 29788 2990
rect 29734 2952 29736 2961
rect 29788 2952 29790 2961
rect 29734 2887 29790 2896
rect 30116 2774 30144 19314
rect 30208 17134 30236 19314
rect 30196 17128 30248 17134
rect 30196 17070 30248 17076
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30208 14482 30236 14758
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30852 12306 30880 21422
rect 32140 17882 32168 37198
rect 32232 37126 32260 39200
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32416 33114 32444 37198
rect 32876 37108 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 33140 37120 33192 37126
rect 32876 37080 33140 37108
rect 34440 37108 34468 39222
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34888 37256 34940 37262
rect 34888 37198 34940 37204
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 33140 37062 33192 37068
rect 34520 37062 34572 37068
rect 34900 36650 34928 37198
rect 35452 36786 35480 39200
rect 35532 37256 35584 37262
rect 35532 37198 35584 37204
rect 35440 36780 35492 36786
rect 35440 36722 35492 36728
rect 34888 36644 34940 36650
rect 34888 36586 34940 36592
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32416 26042 32444 31282
rect 33152 30802 33180 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 33324 36100 33376 36106
rect 33324 36042 33376 36048
rect 33336 31482 33364 36042
rect 34520 35488 34572 35494
rect 34520 35430 34572 35436
rect 33784 34604 33836 34610
rect 33784 34546 33836 34552
rect 33324 31476 33376 31482
rect 33324 31418 33376 31424
rect 33140 30796 33192 30802
rect 33140 30738 33192 30744
rect 33796 29850 33824 34546
rect 34532 30734 34560 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34520 30728 34572 30734
rect 34520 30670 34572 30676
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 33784 29844 33836 29850
rect 33784 29786 33836 29792
rect 32496 29640 32548 29646
rect 32496 29582 32548 29588
rect 35440 29640 35492 29646
rect 35440 29582 35492 29588
rect 32404 26036 32456 26042
rect 32404 25978 32456 25984
rect 32508 25498 32536 29582
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35348 28076 35400 28082
rect 35348 28018 35400 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27130 35388 28018
rect 35348 27124 35400 27130
rect 35348 27066 35400 27072
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35452 26586 35480 29582
rect 35544 28966 35572 37198
rect 36096 37126 36124 39200
rect 37384 37126 37412 39200
rect 38290 38856 38346 38865
rect 38290 38791 38346 38800
rect 38106 37496 38162 37505
rect 38106 37431 38162 37440
rect 37464 37256 37516 37262
rect 37464 37198 37516 37204
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 37372 37120 37424 37126
rect 37372 37062 37424 37068
rect 37476 36922 37504 37198
rect 37464 36916 37516 36922
rect 37464 36858 37516 36864
rect 38120 36854 38148 37431
rect 38108 36848 38160 36854
rect 38108 36790 38160 36796
rect 36360 36780 36412 36786
rect 36360 36722 36412 36728
rect 36268 29164 36320 29170
rect 36268 29106 36320 29112
rect 35532 28960 35584 28966
rect 35532 28902 35584 28908
rect 36280 28218 36308 29106
rect 36268 28212 36320 28218
rect 36268 28154 36320 28160
rect 35440 26580 35492 26586
rect 35440 26522 35492 26528
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 32496 25492 32548 25498
rect 32496 25434 32548 25440
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 33980 20466 34008 21082
rect 33968 20460 34020 20466
rect 33968 20402 34020 20408
rect 33508 20256 33560 20262
rect 33508 20198 33560 20204
rect 32128 17876 32180 17882
rect 32128 17818 32180 17824
rect 30840 12300 30892 12306
rect 30840 12242 30892 12248
rect 33232 11756 33284 11762
rect 33232 11698 33284 11704
rect 33244 11354 33272 11698
rect 33232 11348 33284 11354
rect 33232 11290 33284 11296
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32128 9172 32180 9178
rect 32128 9114 32180 9120
rect 31576 7744 31628 7750
rect 31576 7686 31628 7692
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30380 6384 30432 6390
rect 30380 6326 30432 6332
rect 30392 5710 30420 6326
rect 30470 6216 30526 6225
rect 30470 6151 30526 6160
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30484 5302 30512 6151
rect 30668 6089 30696 6598
rect 30654 6080 30710 6089
rect 30654 6015 30710 6024
rect 30654 5808 30710 5817
rect 30654 5743 30710 5752
rect 30564 5568 30616 5574
rect 30564 5510 30616 5516
rect 30472 5296 30524 5302
rect 30472 5238 30524 5244
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30378 4312 30434 4321
rect 30378 4247 30434 4256
rect 30392 3738 30420 4247
rect 30380 3732 30432 3738
rect 30380 3674 30432 3680
rect 30024 2746 30144 2774
rect 30024 2514 30052 2746
rect 30484 2553 30512 4422
rect 30576 4146 30604 5510
rect 30668 4486 30696 5743
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 31036 5098 31064 5646
rect 31588 5370 31616 7686
rect 31668 7336 31720 7342
rect 31668 7278 31720 7284
rect 31576 5364 31628 5370
rect 31576 5306 31628 5312
rect 31680 5234 31708 7278
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 31024 5092 31076 5098
rect 31024 5034 31076 5040
rect 31220 4622 31248 5170
rect 31298 4992 31354 5001
rect 31298 4927 31354 4936
rect 30748 4616 30800 4622
rect 31208 4616 31260 4622
rect 30748 4558 30800 4564
rect 31114 4584 31170 4593
rect 30656 4480 30708 4486
rect 30656 4422 30708 4428
rect 30760 4146 30788 4558
rect 31208 4558 31260 4564
rect 31114 4519 31116 4528
rect 31168 4519 31170 4528
rect 31116 4490 31168 4496
rect 30564 4140 30616 4146
rect 30564 4082 30616 4088
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30760 4049 30788 4082
rect 31116 4072 31168 4078
rect 30746 4040 30802 4049
rect 31116 4014 31168 4020
rect 30746 3975 30802 3984
rect 30564 3936 30616 3942
rect 30564 3878 30616 3884
rect 30470 2544 30526 2553
rect 30012 2508 30064 2514
rect 30470 2479 30526 2488
rect 30012 2450 30064 2456
rect 29552 2304 29604 2310
rect 29552 2246 29604 2252
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 29276 1216 29328 1222
rect 29276 1158 29328 1164
rect 30300 800 30328 2246
rect 30576 2009 30604 3878
rect 30656 3664 30708 3670
rect 30708 3612 30880 3618
rect 30656 3606 30880 3612
rect 30668 3590 30880 3606
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30760 2922 30788 3334
rect 30852 3058 30880 3590
rect 31128 3482 31156 4014
rect 31220 3534 31248 4558
rect 31312 3942 31340 4927
rect 31864 4826 31892 5646
rect 31852 4820 31904 4826
rect 31852 4762 31904 4768
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 31680 4214 31708 4558
rect 31668 4208 31720 4214
rect 31668 4150 31720 4156
rect 31576 4140 31628 4146
rect 31576 4082 31628 4088
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31036 3454 31156 3482
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 31392 3528 31444 3534
rect 31392 3470 31444 3476
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30748 2916 30800 2922
rect 30748 2858 30800 2864
rect 30852 2038 30880 2994
rect 31036 2774 31064 3454
rect 31220 3398 31248 3470
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 31208 3392 31260 3398
rect 31208 3334 31260 3340
rect 30944 2746 31064 2774
rect 30840 2032 30892 2038
rect 30562 2000 30618 2009
rect 30840 1974 30892 1980
rect 30562 1935 30618 1944
rect 30944 800 30972 2746
rect 31128 1970 31156 3334
rect 31220 2990 31248 3334
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 31116 1964 31168 1970
rect 31116 1906 31168 1912
rect 31404 1358 31432 3470
rect 31588 3074 31616 4082
rect 31588 3058 31708 3074
rect 31588 3052 31720 3058
rect 31588 3046 31668 3052
rect 31668 2994 31720 3000
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 31392 1352 31444 1358
rect 31392 1294 31444 1300
rect 31680 1018 31708 2790
rect 32140 2650 32168 9114
rect 32312 5840 32364 5846
rect 32312 5782 32364 5788
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 32324 2446 32352 5782
rect 32416 4146 32444 9522
rect 33048 9104 33100 9110
rect 33048 9046 33100 9052
rect 32496 6112 32548 6118
rect 32496 6054 32548 6060
rect 32508 4622 32536 6054
rect 32588 5296 32640 5302
rect 32588 5238 32640 5244
rect 32496 4616 32548 4622
rect 32496 4558 32548 4564
rect 32404 4140 32456 4146
rect 32404 4082 32456 4088
rect 32494 3632 32550 3641
rect 32494 3567 32550 3576
rect 32508 3534 32536 3567
rect 32600 3534 32628 5238
rect 32862 4176 32918 4185
rect 32862 4111 32918 4120
rect 32772 3596 32824 3602
rect 32772 3538 32824 3544
rect 32496 3528 32548 3534
rect 32496 3470 32548 3476
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 32784 3058 32812 3538
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32876 2854 32904 4111
rect 33060 4078 33088 9046
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 33048 3936 33100 3942
rect 32954 3904 33010 3913
rect 33048 3878 33100 3884
rect 32954 3839 33010 3848
rect 32968 3074 32996 3839
rect 33060 3194 33088 3878
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 32968 3046 33272 3074
rect 33140 2984 33192 2990
rect 33060 2932 33140 2938
rect 33060 2926 33192 2932
rect 33060 2910 33180 2926
rect 33244 2922 33272 3046
rect 33232 2916 33284 2922
rect 32404 2848 32456 2854
rect 32404 2790 32456 2796
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 31668 1012 31720 1018
rect 31668 954 31720 960
rect 32232 800 32260 2246
rect 32416 1154 32444 2790
rect 33060 2378 33088 2910
rect 33232 2858 33284 2864
rect 33520 2446 33548 20198
rect 34716 19854 34744 21830
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21004 34848 21010
rect 34796 20946 34848 20952
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34520 9716 34572 9722
rect 34520 9658 34572 9664
rect 34532 8974 34560 9658
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34520 7200 34572 7206
rect 34520 7142 34572 7148
rect 34336 6860 34388 6866
rect 34336 6802 34388 6808
rect 33784 5024 33836 5030
rect 33784 4966 33836 4972
rect 33600 4752 33652 4758
rect 33598 4720 33600 4729
rect 33652 4720 33654 4729
rect 33598 4655 33654 4664
rect 33796 4622 33824 4966
rect 33784 4616 33836 4622
rect 33784 4558 33836 4564
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33612 3233 33640 3334
rect 33598 3224 33654 3233
rect 33598 3159 33654 3168
rect 33704 3126 33732 3334
rect 34348 3194 34376 6802
rect 34532 6798 34560 7142
rect 34520 6792 34572 6798
rect 34520 6734 34572 6740
rect 34612 5568 34664 5574
rect 34612 5510 34664 5516
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34336 3188 34388 3194
rect 34336 3130 34388 3136
rect 33692 3120 33744 3126
rect 33692 3062 33744 3068
rect 34440 3058 34468 3402
rect 34428 3052 34480 3058
rect 34428 2994 34480 3000
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 33048 2372 33100 2378
rect 33048 2314 33100 2320
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 32404 1148 32456 1154
rect 32404 1090 32456 1096
rect 33520 800 33548 2246
rect 34164 800 34192 2246
rect 34532 1290 34560 2790
rect 34624 2514 34652 5510
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34716 2825 34744 3470
rect 34702 2816 34758 2825
rect 34702 2751 34758 2760
rect 34612 2508 34664 2514
rect 34612 2450 34664 2456
rect 34808 2446 34836 20946
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35992 18828 36044 18834
rect 35992 18770 36044 18776
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35622 5400 35678 5409
rect 35622 5335 35678 5344
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35636 3194 35664 5335
rect 35820 4010 35848 8434
rect 36004 6914 36032 18770
rect 36372 15570 36400 36722
rect 36820 36576 36872 36582
rect 36820 36518 36872 36524
rect 37280 36576 37332 36582
rect 37280 36518 37332 36524
rect 36832 36174 36860 36518
rect 36820 36168 36872 36174
rect 36820 36110 36872 36116
rect 37292 33862 37320 36518
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38016 35692 38068 35698
rect 38016 35634 38068 35640
rect 37280 33856 37332 33862
rect 37280 33798 37332 33804
rect 38028 33114 38056 35634
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38304 35086 38332 38791
rect 38672 35766 38700 39200
rect 39316 36378 39344 39200
rect 39304 36372 39356 36378
rect 39304 36314 39356 36320
rect 38660 35760 38712 35766
rect 38660 35702 38712 35708
rect 38292 35080 38344 35086
rect 38292 35022 38344 35028
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38016 33108 38068 33114
rect 38016 33050 38068 33056
rect 36820 32904 36872 32910
rect 36820 32846 36872 32852
rect 36832 32570 36860 32846
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 37832 32768 37884 32774
rect 38120 32745 38148 32778
rect 37832 32710 37884 32716
rect 38106 32736 38162 32745
rect 36820 32564 36872 32570
rect 36820 32506 36872 32512
rect 36728 32428 36780 32434
rect 36728 32370 36780 32376
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36740 12918 36768 32370
rect 37372 27328 37424 27334
rect 37372 27270 37424 27276
rect 37384 21554 37412 27270
rect 37740 27056 37792 27062
rect 37740 26998 37792 27004
rect 37464 24200 37516 24206
rect 37464 24142 37516 24148
rect 37476 23905 37504 24142
rect 37462 23896 37518 23905
rect 37462 23831 37518 23840
rect 37372 21548 37424 21554
rect 37372 21490 37424 21496
rect 37280 17672 37332 17678
rect 37280 17614 37332 17620
rect 37188 15496 37240 15502
rect 37188 15438 37240 15444
rect 37200 15065 37228 15438
rect 37186 15056 37242 15065
rect 37186 14991 37242 15000
rect 37292 13938 37320 17614
rect 37752 15570 37780 26998
rect 37844 20466 37872 32710
rect 38106 32671 38162 32680
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 38120 32065 38148 32370
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38106 32056 38162 32065
rect 38106 31991 38162 32000
rect 38212 31958 38240 32166
rect 38200 31952 38252 31958
rect 38200 31894 38252 31900
rect 38016 30728 38068 30734
rect 38016 30670 38068 30676
rect 38198 30696 38254 30705
rect 38028 30122 38056 30670
rect 38198 30631 38254 30640
rect 38212 30598 38240 30631
rect 38200 30592 38252 30598
rect 38200 30534 38252 30540
rect 38016 30116 38068 30122
rect 38016 30058 38068 30064
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38212 29345 38240 29446
rect 38198 29336 38254 29345
rect 38198 29271 38254 29280
rect 38200 29028 38252 29034
rect 38200 28970 38252 28976
rect 38212 28665 38240 28970
rect 38198 28656 38254 28665
rect 38198 28591 38254 28600
rect 38292 27464 38344 27470
rect 38292 27406 38344 27412
rect 38304 27305 38332 27406
rect 38290 27296 38346 27305
rect 38290 27231 38346 27240
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38108 26240 38160 26246
rect 38108 26182 38160 26188
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 37924 24200 37976 24206
rect 37924 24142 37976 24148
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37936 16574 37964 24142
rect 38028 23526 38056 25230
rect 38016 23520 38068 23526
rect 38016 23462 38068 23468
rect 38120 22030 38148 26182
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38290 25871 38346 25880
rect 38198 25256 38254 25265
rect 38198 25191 38254 25200
rect 38212 25158 38240 25191
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38108 22024 38160 22030
rect 38108 21966 38160 21972
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 38200 20800 38252 20806
rect 38200 20742 38252 20748
rect 38212 20505 38240 20742
rect 38198 20496 38254 20505
rect 38198 20431 38254 20440
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 38120 19145 38148 19314
rect 38200 19168 38252 19174
rect 38106 19136 38162 19145
rect 38200 19110 38252 19116
rect 38106 19071 38162 19080
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 38120 16658 38148 16934
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 37936 16546 38056 16574
rect 37740 15564 37792 15570
rect 37740 15506 37792 15512
rect 38028 15026 38056 16546
rect 38016 15020 38068 15026
rect 38016 14962 38068 14968
rect 37924 14816 37976 14822
rect 37924 14758 37976 14764
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 37188 13864 37240 13870
rect 37188 13806 37240 13812
rect 37200 13705 37228 13806
rect 37186 13696 37242 13705
rect 37186 13631 37242 13640
rect 36728 12912 36780 12918
rect 36728 12854 36780 12860
rect 36912 12844 36964 12850
rect 36912 12786 36964 12792
rect 36924 11898 36952 12786
rect 36912 11892 36964 11898
rect 36912 11834 36964 11840
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 37844 10266 37872 10610
rect 37832 10260 37884 10266
rect 37832 10202 37884 10208
rect 36084 8968 36136 8974
rect 36084 8910 36136 8916
rect 36096 8634 36124 8910
rect 36268 8832 36320 8838
rect 36268 8774 36320 8780
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 36280 8498 36308 8774
rect 36268 8492 36320 8498
rect 36268 8434 36320 8440
rect 35912 6886 36032 6914
rect 35808 4004 35860 4010
rect 35808 3946 35860 3952
rect 35716 3936 35768 3942
rect 35716 3878 35768 3884
rect 35728 3534 35756 3878
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 35624 3188 35676 3194
rect 35624 3130 35676 3136
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34520 1284 34572 1290
rect 34520 1226 34572 1232
rect 35452 800 35480 2926
rect 35544 2281 35572 2994
rect 35912 2446 35940 6886
rect 36728 6180 36780 6186
rect 36728 6122 36780 6128
rect 36740 3738 36768 6122
rect 36728 3732 36780 3738
rect 36728 3674 36780 3680
rect 37936 3534 37964 14758
rect 38028 14618 38056 14962
rect 38016 14612 38068 14618
rect 38016 14554 38068 14560
rect 38212 14346 38240 19110
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 38304 17105 38332 17138
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 38292 16108 38344 16114
rect 38292 16050 38344 16056
rect 38304 15745 38332 16050
rect 38290 15736 38346 15745
rect 38290 15671 38346 15680
rect 38200 14340 38252 14346
rect 38200 14282 38252 14288
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38016 11008 38068 11014
rect 38304 10985 38332 11086
rect 38016 10950 38068 10956
rect 38290 10976 38346 10985
rect 38028 10062 38056 10950
rect 38290 10911 38346 10920
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 38212 10305 38240 10406
rect 38198 10296 38254 10305
rect 38198 10231 38254 10240
rect 38016 10056 38068 10062
rect 38016 9998 38068 10004
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38212 7585 38240 7686
rect 38198 7576 38254 7585
rect 38198 7511 38254 7520
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38304 6905 38332 7346
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38014 6488 38070 6497
rect 38014 6423 38070 6432
rect 38028 5710 38056 6423
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 38016 5568 38068 5574
rect 38200 5568 38252 5574
rect 38016 5510 38068 5516
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38028 4622 38056 5510
rect 38198 5471 38254 5480
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 38212 4185 38240 4422
rect 38198 4176 38254 4185
rect 38198 4111 38254 4120
rect 38292 4140 38344 4146
rect 38292 4082 38344 4088
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37924 3528 37976 3534
rect 38304 3505 38332 4082
rect 37924 3470 37976 3476
rect 38290 3496 38346 3505
rect 36636 3392 36688 3398
rect 36636 3334 36688 3340
rect 36648 3058 36676 3334
rect 36636 3052 36688 3058
rect 36636 2994 36688 3000
rect 36176 2848 36228 2854
rect 36176 2790 36228 2796
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35530 2272 35586 2281
rect 35530 2207 35586 2216
rect 36188 1698 36216 2790
rect 37188 2576 37240 2582
rect 37188 2518 37240 2524
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36176 1692 36228 1698
rect 36176 1634 36228 1640
rect 36740 800 36768 2246
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 37200 105 37228 2518
rect 37384 800 37412 3470
rect 38290 3431 38346 3440
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37476 1465 37504 2382
rect 38212 2145 38240 3334
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38198 2136 38254 2145
rect 38198 2071 38254 2080
rect 37462 1456 37518 1465
rect 37462 1391 37518 1400
rect 38672 800 38700 2790
rect 37370 200 37426 800
rect 38658 200 38714 800
rect 37186 96 37242 105
rect 37186 31 37242 40
<< via2 >>
rect 3146 39480 3202 39536
rect 1582 38800 1638 38856
rect 1766 37440 1822 37496
rect 1766 36116 1768 36136
rect 1768 36116 1820 36136
rect 1820 36116 1822 36136
rect 1766 36080 1822 36116
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 1766 34040 1822 34096
rect 1766 32716 1768 32736
rect 1768 32716 1820 32736
rect 1820 32716 1822 32736
rect 1766 32680 1822 32716
rect 1766 32000 1822 32056
rect 1766 30640 1822 30696
rect 1766 29280 1822 29336
rect 1766 28600 1822 28656
rect 1766 27240 1822 27296
rect 1766 25880 1822 25936
rect 1766 24556 1768 24576
rect 1768 24556 1820 24576
rect 1820 24556 1822 24576
rect 1766 24520 1822 24556
rect 1766 23840 1822 23896
rect 1674 22480 1730 22536
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 2502 22500 2558 22536
rect 2502 22480 2504 22500
rect 2504 22480 2556 22500
rect 2556 22480 2558 22500
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1766 21120 1822 21176
rect 1766 20440 1822 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1766 19080 1822 19136
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1766 17720 1822 17776
rect 1582 17076 1584 17096
rect 1584 17076 1636 17096
rect 1636 17076 1638 17096
rect 1582 17040 1638 17076
rect 1582 16108 1638 16144
rect 1582 16088 1584 16108
rect 1584 16088 1636 16108
rect 1636 16088 1638 16108
rect 1766 15680 1822 15736
rect 2134 15272 2190 15328
rect 1766 14320 1822 14376
rect 1766 13676 1768 13696
rect 1768 13676 1820 13696
rect 1820 13676 1822 13696
rect 1766 13640 1822 13676
rect 1766 12280 1822 12336
rect 1582 10920 1638 10976
rect 1582 10784 1638 10840
rect 1766 10240 1822 10296
rect 1858 8200 1914 8256
rect 1582 6840 1638 6896
rect 2686 12960 2742 13016
rect 2686 8336 2742 8392
rect 2870 8916 2872 8936
rect 2872 8916 2924 8936
rect 2924 8916 2926 8936
rect 2870 8880 2926 8916
rect 2778 7520 2834 7576
rect 2778 4120 2834 4176
rect 2042 3596 2098 3632
rect 2042 3576 2044 3596
rect 2044 3576 2096 3596
rect 2096 3576 2098 3596
rect 4158 17040 4214 17096
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 2962 5480 3018 5536
rect 2870 3440 2926 3496
rect 2042 3304 2098 3360
rect 2778 2100 2834 2136
rect 2778 2080 2780 2100
rect 2780 2080 2832 2100
rect 2832 2080 2834 2100
rect 3606 6316 3662 6352
rect 3606 6296 3608 6316
rect 3608 6296 3660 6316
rect 3660 6296 3662 6316
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4342 15308 4344 15328
rect 4344 15308 4396 15328
rect 4396 15308 4398 15328
rect 4342 15272 4398 15308
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4618 14592 4674 14648
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4158 11056 4214 11112
rect 4894 16496 4950 16552
rect 4710 12688 4766 12744
rect 4710 12588 4712 12608
rect 4712 12588 4764 12608
rect 4764 12588 4766 12608
rect 4710 12552 4766 12588
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 3882 6704 3938 6760
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4710 10376 4766 10432
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4526 6568 4582 6624
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4526 4664 4582 4720
rect 4526 4256 4582 4312
rect 3790 3984 3846 4040
rect 3330 856 3386 912
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5262 16496 5318 16552
rect 4986 10920 5042 10976
rect 4894 10104 4950 10160
rect 4986 9460 4988 9480
rect 4988 9460 5040 9480
rect 5040 9460 5042 9480
rect 4986 9424 5042 9460
rect 4986 9172 5042 9208
rect 4986 9152 4988 9172
rect 4988 9152 5040 9172
rect 5040 9152 5042 9172
rect 5446 14048 5502 14104
rect 5630 13504 5686 13560
rect 5630 12688 5686 12744
rect 5354 12144 5410 12200
rect 5262 11872 5318 11928
rect 5262 9696 5318 9752
rect 4894 3460 4950 3496
rect 4894 3440 4896 3460
rect 4896 3440 4948 3460
rect 4948 3440 4950 3460
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 3974 1672 4030 1728
rect 5446 10920 5502 10976
rect 5814 14184 5870 14240
rect 6090 13640 6146 13696
rect 6090 13232 6146 13288
rect 6182 12552 6238 12608
rect 5538 4800 5594 4856
rect 6642 17740 6698 17776
rect 6642 17720 6644 17740
rect 6644 17720 6696 17740
rect 6696 17720 6698 17740
rect 6550 16652 6606 16688
rect 6550 16632 6552 16652
rect 6552 16632 6604 16652
rect 6604 16632 6606 16652
rect 6550 13640 6606 13696
rect 6918 15272 6974 15328
rect 6458 12144 6514 12200
rect 6090 4664 6146 4720
rect 6274 5752 6330 5808
rect 5262 2932 5264 2952
rect 5264 2932 5316 2952
rect 5316 2932 5318 2952
rect 5262 2896 5318 2932
rect 5906 2372 5962 2408
rect 5906 2352 5908 2372
rect 5908 2352 5960 2372
rect 5960 2352 5962 2372
rect 6734 10804 6790 10840
rect 6734 10784 6736 10804
rect 6736 10784 6788 10804
rect 6788 10784 6790 10804
rect 6734 10376 6790 10432
rect 6918 9696 6974 9752
rect 6826 8880 6882 8936
rect 7378 16244 7434 16280
rect 7378 16224 7380 16244
rect 7380 16224 7432 16244
rect 7432 16224 7434 16244
rect 7286 13948 7288 13968
rect 7288 13948 7340 13968
rect 7340 13948 7342 13968
rect 7286 13912 7342 13948
rect 7562 17740 7618 17776
rect 7562 17720 7564 17740
rect 7564 17720 7616 17740
rect 7616 17720 7618 17740
rect 6826 6160 6882 6216
rect 6734 5888 6790 5944
rect 6826 5616 6882 5672
rect 6826 3068 6828 3088
rect 6828 3068 6880 3088
rect 6880 3068 6882 3088
rect 6826 3032 6882 3068
rect 7838 15428 7894 15464
rect 7838 15408 7840 15428
rect 7840 15408 7892 15428
rect 7892 15408 7894 15428
rect 8206 17992 8262 18048
rect 8206 16532 8208 16552
rect 8208 16532 8260 16552
rect 8260 16532 8262 16552
rect 8206 16496 8262 16532
rect 8482 17448 8538 17504
rect 8482 17312 8538 17368
rect 8206 15272 8262 15328
rect 7930 13368 7986 13424
rect 7838 12144 7894 12200
rect 7562 11192 7618 11248
rect 7470 10784 7526 10840
rect 7378 6604 7380 6624
rect 7380 6604 7432 6624
rect 7432 6604 7434 6624
rect 7378 6568 7434 6604
rect 7286 5772 7342 5808
rect 7286 5752 7288 5772
rect 7288 5752 7340 5772
rect 7340 5752 7342 5772
rect 8574 15680 8630 15736
rect 8482 15544 8538 15600
rect 8482 14864 8538 14920
rect 8298 14728 8354 14784
rect 8206 14456 8262 14512
rect 8390 14592 8446 14648
rect 8482 14220 8484 14240
rect 8484 14220 8536 14240
rect 8536 14220 8538 14240
rect 8482 14184 8538 14220
rect 8390 13776 8446 13832
rect 8390 12416 8446 12472
rect 8114 11872 8170 11928
rect 8022 11464 8078 11520
rect 8206 10412 8208 10432
rect 8208 10412 8260 10432
rect 8260 10412 8262 10432
rect 8206 10376 8262 10412
rect 8022 10104 8078 10160
rect 8206 10240 8262 10296
rect 8298 6180 8354 6216
rect 8298 6160 8300 6180
rect 8300 6160 8352 6180
rect 8352 6160 8354 6180
rect 8206 5616 8262 5672
rect 9034 19624 9090 19680
rect 9218 19796 9220 19816
rect 9220 19796 9272 19816
rect 9272 19796 9274 19816
rect 9218 19760 9274 19796
rect 9126 19318 9182 19374
rect 9034 18808 9090 18864
rect 9034 17448 9090 17504
rect 8758 13368 8814 13424
rect 8666 10784 8722 10840
rect 8574 8472 8630 8528
rect 8666 6840 8722 6896
rect 8574 5480 8630 5536
rect 8298 3984 8354 4040
rect 7470 2896 7526 2952
rect 8850 5908 8906 5944
rect 8850 5888 8852 5908
rect 8852 5888 8904 5908
rect 8904 5888 8906 5908
rect 8758 4256 8814 4312
rect 8574 3168 8630 3224
rect 9218 15272 9274 15328
rect 9218 15000 9274 15056
rect 9218 14592 9274 14648
rect 9126 13640 9182 13696
rect 9034 13504 9090 13560
rect 9034 11600 9090 11656
rect 9034 11192 9090 11248
rect 9678 20984 9734 21040
rect 9678 20748 9680 20768
rect 9680 20748 9732 20768
rect 9732 20748 9734 20768
rect 9678 20712 9734 20748
rect 9494 19080 9550 19136
rect 9494 18808 9550 18864
rect 9402 16768 9458 16824
rect 9402 16360 9458 16416
rect 9862 20304 9918 20360
rect 14922 37204 14924 37224
rect 14924 37204 14976 37224
rect 14976 37204 14978 37224
rect 14922 37168 14978 37204
rect 10874 24112 10930 24168
rect 10046 17060 10102 17096
rect 10046 17040 10048 17060
rect 10048 17040 10100 17060
rect 10100 17040 10102 17060
rect 9862 16360 9918 16416
rect 9494 15816 9550 15872
rect 9494 13776 9550 13832
rect 9402 13504 9458 13560
rect 9586 13504 9642 13560
rect 9770 15136 9826 15192
rect 10138 14592 10194 14648
rect 10322 15680 10378 15736
rect 10966 21684 11022 21720
rect 10966 21664 10968 21684
rect 10968 21664 11020 21684
rect 11020 21664 11022 21684
rect 10874 20712 10930 20768
rect 10966 18672 11022 18728
rect 10966 18400 11022 18456
rect 10230 14320 10286 14376
rect 10046 14048 10102 14104
rect 10138 13948 10140 13968
rect 10140 13948 10192 13968
rect 10192 13948 10194 13968
rect 10138 13912 10194 13948
rect 10046 12960 10102 13016
rect 9770 12824 9826 12880
rect 9678 12280 9734 12336
rect 9494 10920 9550 10976
rect 9218 9832 9274 9888
rect 9126 9696 9182 9752
rect 9310 9560 9366 9616
rect 9402 9288 9458 9344
rect 9494 8200 9550 8256
rect 9770 9288 9826 9344
rect 9678 9016 9734 9072
rect 9678 8628 9734 8664
rect 9678 8608 9680 8628
rect 9680 8608 9732 8628
rect 9732 8608 9734 8628
rect 9126 3440 9182 3496
rect 10046 9016 10102 9072
rect 10690 17040 10746 17096
rect 10506 14320 10562 14376
rect 10414 11872 10470 11928
rect 10230 10104 10286 10160
rect 10230 9596 10232 9616
rect 10232 9596 10284 9616
rect 10284 9596 10286 9616
rect 10230 9560 10286 9596
rect 10046 4548 10102 4584
rect 10046 4528 10048 4548
rect 10048 4528 10100 4548
rect 10100 4528 10102 4548
rect 10414 8880 10470 8936
rect 10690 14320 10746 14376
rect 10874 15000 10930 15056
rect 11058 16768 11114 16824
rect 11610 19080 11666 19136
rect 11702 17992 11758 18048
rect 11150 16632 11206 16688
rect 11150 16496 11206 16552
rect 11426 15272 11482 15328
rect 11426 14456 11482 14512
rect 10966 12552 11022 12608
rect 11058 12044 11060 12064
rect 11060 12044 11112 12064
rect 11112 12044 11114 12064
rect 11058 12008 11114 12044
rect 10690 7928 10746 7984
rect 11794 17448 11850 17504
rect 11978 17720 12034 17776
rect 11518 12688 11574 12744
rect 11426 12552 11482 12608
rect 11334 12144 11390 12200
rect 10966 9424 11022 9480
rect 10690 3712 10746 3768
rect 11150 8200 11206 8256
rect 11150 6840 11206 6896
rect 10966 4156 10968 4176
rect 10968 4156 11020 4176
rect 11020 4156 11022 4176
rect 10966 4120 11022 4156
rect 12346 24132 12402 24168
rect 12346 24112 12348 24132
rect 12348 24112 12400 24132
rect 12400 24112 12402 24132
rect 12254 20032 12310 20088
rect 11702 13096 11758 13152
rect 12346 17620 12348 17640
rect 12348 17620 12400 17640
rect 12400 17620 12402 17640
rect 12346 17584 12402 17620
rect 12530 17312 12586 17368
rect 12438 17176 12494 17232
rect 12530 14048 12586 14104
rect 12254 12552 12310 12608
rect 12162 12416 12218 12472
rect 11794 12280 11850 12336
rect 11702 10376 11758 10432
rect 11426 6976 11482 7032
rect 11058 4004 11114 4040
rect 11058 3984 11060 4004
rect 11060 3984 11112 4004
rect 11112 3984 11114 4004
rect 11058 3612 11060 3632
rect 11060 3612 11112 3632
rect 11112 3612 11114 3632
rect 11058 3576 11114 3612
rect 11978 9424 12034 9480
rect 11886 8880 11942 8936
rect 12438 12980 12494 13016
rect 12438 12960 12440 12980
rect 12440 12960 12492 12980
rect 12492 12960 12494 12980
rect 13450 18808 13506 18864
rect 13174 18536 13230 18592
rect 12714 14320 12770 14376
rect 13450 18400 13506 18456
rect 12990 14884 13046 14920
rect 12990 14864 12992 14884
rect 12992 14864 13044 14884
rect 13044 14864 13046 14884
rect 13266 16788 13322 16824
rect 13266 16768 13268 16788
rect 13268 16768 13320 16788
rect 13320 16768 13322 16788
rect 13266 15272 13322 15328
rect 13910 21392 13966 21448
rect 13726 20848 13782 20904
rect 13726 19352 13782 19408
rect 13358 13096 13414 13152
rect 13266 12824 13322 12880
rect 12070 6860 12126 6896
rect 12070 6840 12072 6860
rect 12072 6840 12124 6860
rect 12124 6840 12126 6860
rect 12162 6432 12218 6488
rect 11886 4664 11942 4720
rect 11610 2760 11666 2816
rect 12438 6452 12494 6488
rect 12438 6432 12440 6452
rect 12440 6432 12492 6452
rect 12492 6432 12494 6452
rect 12530 3576 12586 3632
rect 12990 10512 13046 10568
rect 13450 10920 13506 10976
rect 13450 9968 13506 10024
rect 13266 9288 13322 9344
rect 13726 14592 13782 14648
rect 13726 14340 13782 14376
rect 13726 14320 13728 14340
rect 13728 14320 13780 14340
rect 13780 14320 13782 14340
rect 13542 9560 13598 9616
rect 14830 21664 14886 21720
rect 14738 20984 14794 21040
rect 14278 19796 14280 19816
rect 14280 19796 14332 19816
rect 14332 19796 14334 19816
rect 14278 19760 14334 19796
rect 14646 19488 14702 19544
rect 14554 19236 14610 19272
rect 14554 19216 14556 19236
rect 14556 19216 14608 19236
rect 14608 19216 14610 19236
rect 15014 20324 15070 20360
rect 15014 20304 15016 20324
rect 15016 20304 15068 20324
rect 15068 20304 15070 20324
rect 14462 18128 14518 18184
rect 14462 16652 14518 16688
rect 14462 16632 14464 16652
rect 14464 16632 14516 16652
rect 14516 16632 14518 16652
rect 14094 13912 14150 13968
rect 14094 13504 14150 13560
rect 13818 9288 13874 9344
rect 12806 6976 12862 7032
rect 13266 7656 13322 7712
rect 13266 7248 13322 7304
rect 12806 3848 12862 3904
rect 12714 3712 12770 3768
rect 12622 2760 12678 2816
rect 13082 3576 13138 3632
rect 13726 5616 13782 5672
rect 14554 15136 14610 15192
rect 14646 15000 14702 15056
rect 14462 14184 14518 14240
rect 14646 13948 14648 13968
rect 14648 13948 14700 13968
rect 14700 13948 14702 13968
rect 14646 13912 14702 13948
rect 14462 12008 14518 12064
rect 14002 5208 14058 5264
rect 13818 4700 13820 4720
rect 13820 4700 13872 4720
rect 13872 4700 13874 4720
rect 13818 4664 13874 4700
rect 14278 4664 14334 4720
rect 14646 12280 14702 12336
rect 14554 11328 14610 11384
rect 14830 11056 14886 11112
rect 14738 10956 14740 10976
rect 14740 10956 14792 10976
rect 14792 10956 14794 10976
rect 14738 10920 14794 10956
rect 14830 9288 14886 9344
rect 15014 10784 15070 10840
rect 15014 10104 15070 10160
rect 15382 13640 15438 13696
rect 15290 12144 15346 12200
rect 15198 10512 15254 10568
rect 15106 9832 15162 9888
rect 15566 19488 15622 19544
rect 15658 16632 15714 16688
rect 16026 18808 16082 18864
rect 16118 18400 16174 18456
rect 16118 17040 16174 17096
rect 15382 8472 15438 8528
rect 14646 5364 14702 5400
rect 14646 5344 14648 5364
rect 14648 5344 14700 5364
rect 14700 5344 14702 5364
rect 13542 1944 13598 2000
rect 13726 2488 13782 2544
rect 13726 1808 13782 1864
rect 15014 7404 15070 7440
rect 15014 7384 15016 7404
rect 15016 7384 15068 7404
rect 15068 7384 15070 7404
rect 15934 10784 15990 10840
rect 17590 20848 17646 20904
rect 17498 20032 17554 20088
rect 16946 19080 17002 19136
rect 17498 19352 17554 19408
rect 17222 19236 17278 19272
rect 17222 19216 17224 19236
rect 17224 19216 17276 19236
rect 17276 19216 17278 19236
rect 17314 18164 17316 18184
rect 17316 18164 17368 18184
rect 17368 18164 17370 18184
rect 17314 18128 17370 18164
rect 16946 16496 17002 16552
rect 16762 13640 16818 13696
rect 16394 11872 16450 11928
rect 16302 9288 16358 9344
rect 16118 6160 16174 6216
rect 15842 5888 15898 5944
rect 16578 9172 16634 9208
rect 16578 9152 16580 9172
rect 16580 9152 16632 9172
rect 16632 9152 16634 9172
rect 17038 12960 17094 13016
rect 17038 12724 17040 12744
rect 17040 12724 17092 12744
rect 17092 12724 17094 12744
rect 17038 12688 17094 12724
rect 17130 9460 17132 9480
rect 17132 9460 17184 9480
rect 17184 9460 17186 9480
rect 17130 9424 17186 9460
rect 17590 17448 17646 17504
rect 17682 17312 17738 17368
rect 17498 15000 17554 15056
rect 18050 19760 18106 19816
rect 18050 16088 18106 16144
rect 17958 15272 18014 15328
rect 18234 15272 18290 15328
rect 17314 9696 17370 9752
rect 16486 7928 16542 7984
rect 16486 7112 16542 7168
rect 16670 6724 16726 6760
rect 16670 6704 16672 6724
rect 16672 6704 16724 6724
rect 16724 6704 16726 6724
rect 16578 3848 16634 3904
rect 16578 3596 16634 3632
rect 16578 3576 16580 3596
rect 16580 3576 16632 3596
rect 16632 3576 16634 3596
rect 16486 2760 16542 2816
rect 17774 9152 17830 9208
rect 18602 21392 18658 21448
rect 18418 17992 18474 18048
rect 18418 16768 18474 16824
rect 18234 12280 18290 12336
rect 17498 5752 17554 5808
rect 18326 11348 18382 11384
rect 18326 11328 18328 11348
rect 18328 11328 18380 11348
rect 18380 11328 18382 11348
rect 18694 18536 18750 18592
rect 18234 9016 18290 9072
rect 17866 5108 17868 5128
rect 17868 5108 17920 5128
rect 17920 5108 17922 5128
rect 17866 5072 17922 5108
rect 18234 6840 18290 6896
rect 18142 5344 18198 5400
rect 18878 11464 18934 11520
rect 18694 7248 18750 7304
rect 18786 6296 18842 6352
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19522 17620 19524 17640
rect 19524 17620 19576 17640
rect 19576 17620 19578 17640
rect 19522 17584 19578 17620
rect 21638 23060 21640 23080
rect 21640 23060 21692 23080
rect 21692 23060 21694 23080
rect 21638 23024 21694 23060
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19246 13812 19248 13832
rect 19248 13812 19300 13832
rect 19300 13812 19302 13832
rect 19246 13776 19302 13812
rect 18970 6024 19026 6080
rect 19798 13368 19854 13424
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19430 12316 19432 12336
rect 19432 12316 19484 12336
rect 19484 12316 19486 12336
rect 19430 12280 19486 12316
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20534 16652 20590 16688
rect 20534 16632 20536 16652
rect 20536 16632 20588 16652
rect 20588 16632 20590 16652
rect 20350 14476 20406 14512
rect 20350 14456 20352 14476
rect 20352 14456 20404 14476
rect 20404 14456 20406 14476
rect 19706 9052 19708 9072
rect 19708 9052 19760 9072
rect 19760 9052 19762 9072
rect 19706 9016 19762 9052
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19890 7812 19946 7848
rect 19890 7792 19892 7812
rect 19892 7792 19944 7812
rect 19944 7792 19946 7812
rect 19154 7656 19210 7712
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19522 6840 19578 6896
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20166 8744 20222 8800
rect 20074 5616 20130 5672
rect 19982 5480 20038 5536
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19430 4936 19486 4992
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20350 13504 20406 13560
rect 20350 13232 20406 13288
rect 20902 16496 20958 16552
rect 20718 15444 20720 15464
rect 20720 15444 20772 15464
rect 20772 15444 20774 15464
rect 20718 15408 20774 15444
rect 20810 14048 20866 14104
rect 20718 12844 20774 12880
rect 20718 12824 20720 12844
rect 20720 12824 20772 12844
rect 20772 12824 20774 12844
rect 20534 8608 20590 8664
rect 20350 6568 20406 6624
rect 20350 5208 20406 5264
rect 21546 13912 21602 13968
rect 21270 12144 21326 12200
rect 21086 11872 21142 11928
rect 21086 11736 21142 11792
rect 21270 11736 21326 11792
rect 20718 9560 20774 9616
rect 21086 11192 21142 11248
rect 21270 11056 21326 11112
rect 21178 10648 21234 10704
rect 21454 9288 21510 9344
rect 21178 9016 21234 9072
rect 21362 8744 21418 8800
rect 20626 6840 20682 6896
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19890 2624 19946 2680
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21086 7520 21142 7576
rect 20994 6432 21050 6488
rect 21086 5888 21142 5944
rect 21638 6976 21694 7032
rect 21086 4528 21142 4584
rect 21914 14900 21916 14920
rect 21916 14900 21968 14920
rect 21968 14900 21970 14920
rect 21914 14864 21970 14900
rect 22190 15000 22246 15056
rect 21914 13912 21970 13968
rect 22098 13368 22154 13424
rect 21822 12280 21878 12336
rect 22098 11464 22154 11520
rect 22374 11056 22430 11112
rect 22190 10240 22246 10296
rect 21822 9036 21878 9072
rect 21822 9016 21824 9036
rect 21824 9016 21876 9036
rect 21876 9016 21878 9036
rect 21822 8900 21878 8936
rect 21822 8880 21824 8900
rect 21824 8880 21876 8900
rect 21876 8880 21878 8900
rect 21362 5072 21418 5128
rect 21822 6024 21878 6080
rect 22282 6840 22338 6896
rect 22190 6568 22246 6624
rect 22098 5344 22154 5400
rect 21454 4936 21510 4992
rect 20626 3576 20682 3632
rect 21546 3304 21602 3360
rect 22558 9424 22614 9480
rect 23386 14456 23442 14512
rect 23110 11464 23166 11520
rect 23478 11500 23480 11520
rect 23480 11500 23532 11520
rect 23532 11500 23534 11520
rect 23478 11464 23534 11500
rect 23846 15444 23848 15464
rect 23848 15444 23900 15464
rect 23900 15444 23902 15464
rect 23846 15408 23902 15444
rect 23938 15308 23940 15328
rect 23940 15308 23992 15328
rect 23992 15308 23994 15328
rect 23938 15272 23994 15308
rect 23386 8608 23442 8664
rect 23018 6024 23074 6080
rect 22558 5344 22614 5400
rect 22650 4936 22706 4992
rect 23294 4392 23350 4448
rect 22282 3848 22338 3904
rect 22374 2932 22376 2952
rect 22376 2932 22428 2952
rect 22428 2932 22430 2952
rect 22374 2896 22430 2932
rect 24030 13504 24086 13560
rect 23754 9052 23756 9072
rect 23756 9052 23808 9072
rect 23808 9052 23810 9072
rect 23754 9016 23810 9052
rect 24214 14864 24270 14920
rect 24674 17040 24730 17096
rect 24306 14048 24362 14104
rect 24214 11192 24270 11248
rect 23846 5888 23902 5944
rect 23754 5616 23810 5672
rect 23754 4972 23756 4992
rect 23756 4972 23808 4992
rect 23808 4972 23810 4992
rect 23754 4936 23810 4972
rect 24398 11872 24454 11928
rect 24858 13232 24914 13288
rect 24582 9832 24638 9888
rect 24490 7792 24546 7848
rect 24398 5616 24454 5672
rect 23938 3168 23994 3224
rect 24490 3712 24546 3768
rect 24398 3032 24454 3088
rect 24766 8336 24822 8392
rect 24766 7656 24822 7712
rect 24766 6432 24822 6488
rect 25042 6840 25098 6896
rect 24950 6568 25006 6624
rect 24674 5344 24730 5400
rect 24766 4256 24822 4312
rect 24674 3576 24730 3632
rect 25042 5072 25098 5128
rect 24858 3304 24914 3360
rect 24858 2644 24914 2680
rect 24858 2624 24860 2644
rect 24860 2624 24912 2644
rect 24912 2624 24914 2644
rect 25042 2624 25098 2680
rect 25226 11600 25282 11656
rect 25686 9152 25742 9208
rect 25962 14320 26018 14376
rect 25962 13640 26018 13696
rect 25318 8608 25374 8664
rect 26054 8492 26110 8528
rect 26054 8472 26056 8492
rect 26056 8472 26108 8492
rect 26108 8472 26110 8492
rect 25410 6432 25466 6488
rect 25410 3440 25466 3496
rect 25870 7520 25926 7576
rect 26330 6976 26386 7032
rect 25686 5888 25742 5944
rect 25594 3984 25650 4040
rect 25502 3168 25558 3224
rect 26054 6432 26110 6488
rect 25962 3460 26018 3496
rect 25962 3440 25964 3460
rect 25964 3440 26016 3460
rect 26016 3440 26018 3460
rect 26698 7248 26754 7304
rect 26974 11872 27030 11928
rect 26330 4800 26386 4856
rect 26238 4428 26240 4448
rect 26240 4428 26292 4448
rect 26292 4428 26294 4448
rect 26238 4392 26294 4428
rect 26790 5888 26846 5944
rect 27158 13912 27214 13968
rect 27434 11736 27490 11792
rect 27066 7656 27122 7712
rect 27158 7404 27214 7440
rect 27158 7384 27160 7404
rect 27160 7384 27212 7404
rect 27212 7384 27214 7404
rect 26330 3168 26386 3224
rect 25318 2216 25374 2272
rect 27802 11056 27858 11112
rect 27250 5480 27306 5536
rect 26698 2760 26754 2816
rect 26882 3476 26884 3496
rect 26884 3476 26936 3496
rect 26936 3476 26938 3496
rect 26882 3440 26938 3476
rect 27066 2760 27122 2816
rect 26514 1672 26570 1728
rect 27250 3168 27306 3224
rect 27802 5652 27804 5672
rect 27804 5652 27856 5672
rect 27856 5652 27858 5672
rect 27802 5616 27858 5652
rect 27618 3304 27674 3360
rect 27250 2352 27306 2408
rect 28814 9596 28816 9616
rect 28816 9596 28868 9616
rect 28868 9596 28870 9616
rect 28814 9560 28870 9596
rect 28814 7112 28870 7168
rect 28998 6704 29054 6760
rect 28906 6332 28908 6352
rect 28908 6332 28960 6352
rect 28960 6332 28962 6352
rect 28906 6296 28962 6332
rect 29826 9832 29882 9888
rect 28814 5072 28870 5128
rect 28814 3712 28870 3768
rect 28906 3032 28962 3088
rect 28998 2624 29054 2680
rect 28078 1808 28134 1864
rect 29734 4800 29790 4856
rect 29734 2932 29736 2952
rect 29736 2932 29788 2952
rect 29788 2932 29790 2952
rect 29734 2896 29790 2932
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 38290 38800 38346 38856
rect 38106 37440 38162 37496
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 30470 6160 30526 6216
rect 30654 6024 30710 6080
rect 30654 5752 30710 5808
rect 30378 4256 30434 4312
rect 31298 4936 31354 4992
rect 31114 4548 31170 4584
rect 31114 4528 31116 4548
rect 31116 4528 31168 4548
rect 31168 4528 31170 4548
rect 30746 3984 30802 4040
rect 30470 2488 30526 2544
rect 30562 1944 30618 2000
rect 32494 3576 32550 3632
rect 32862 4120 32918 4176
rect 32954 3848 33010 3904
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 33598 4700 33600 4720
rect 33600 4700 33652 4720
rect 33652 4700 33654 4720
rect 33598 4664 33654 4700
rect 33598 3168 33654 3224
rect 34702 2760 34758 2816
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35622 5344 35678 5400
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 34040 38254 34096
rect 37462 23840 37518 23896
rect 37186 15000 37242 15056
rect 38106 32680 38162 32736
rect 38106 32000 38162 32056
rect 38198 30640 38254 30696
rect 38198 29280 38254 29336
rect 38198 28600 38254 28656
rect 38290 27240 38346 27296
rect 38290 25880 38346 25936
rect 38198 25200 38254 25256
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38290 21800 38346 21856
rect 38198 20440 38254 20496
rect 38106 19080 38162 19136
rect 37186 13640 37242 13696
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 17040 38346 17096
rect 38290 15680 38346 15736
rect 38198 12280 38254 12336
rect 38290 10920 38346 10976
rect 38198 10240 38254 10296
rect 38198 8880 38254 8936
rect 38198 7520 38254 7576
rect 38290 6840 38346 6896
rect 38014 6432 38070 6488
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 38198 4120 38254 4176
rect 35530 2216 35586 2272
rect 38290 3440 38346 3496
rect 38198 2080 38254 2136
rect 37462 1400 37518 1456
rect 37186 40 37242 96
<< metal3 >>
rect 200 39538 800 39568
rect 3141 39538 3207 39541
rect 200 39536 3207 39538
rect 200 39480 3146 39536
rect 3202 39480 3207 39536
rect 200 39478 3207 39480
rect 200 39448 800 39478
rect 3141 39475 3207 39478
rect 200 38858 800 38888
rect 1577 38858 1643 38861
rect 200 38856 1643 38858
rect 200 38800 1582 38856
rect 1638 38800 1643 38856
rect 200 38798 1643 38800
rect 200 38768 800 38798
rect 1577 38795 1643 38798
rect 38285 38858 38351 38861
rect 39200 38858 39800 38888
rect 38285 38856 39800 38858
rect 38285 38800 38290 38856
rect 38346 38800 39800 38856
rect 38285 38798 39800 38800
rect 38285 38795 38351 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 1761 37498 1827 37501
rect 200 37496 1827 37498
rect 200 37440 1766 37496
rect 1822 37440 1827 37496
rect 200 37438 1827 37440
rect 200 37408 800 37438
rect 1761 37435 1827 37438
rect 38101 37498 38167 37501
rect 39200 37498 39800 37528
rect 38101 37496 39800 37498
rect 38101 37440 38106 37496
rect 38162 37440 39800 37496
rect 38101 37438 39800 37440
rect 38101 37435 38167 37438
rect 39200 37408 39800 37438
rect 14917 37228 14983 37229
rect 14917 37226 14964 37228
rect 14872 37224 14964 37226
rect 14872 37168 14922 37224
rect 14872 37166 14964 37168
rect 14917 37164 14964 37166
rect 15028 37164 15034 37228
rect 14917 37163 14983 37164
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 200 36138 800 36168
rect 1761 36138 1827 36141
rect 200 36136 1827 36138
rect 200 36080 1766 36136
rect 1822 36080 1827 36136
rect 200 36078 1827 36080
rect 200 36048 800 36078
rect 1761 36075 1827 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35368 800 35488
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 38101 32738 38167 32741
rect 39200 32738 39800 32768
rect 38101 32736 39800 32738
rect 38101 32680 38106 32736
rect 38162 32680 39800 32736
rect 38101 32678 39800 32680
rect 38101 32675 38167 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38101 32058 38167 32061
rect 39200 32058 39800 32088
rect 38101 32056 39800 32058
rect 38101 32000 38106 32056
rect 38162 32000 39800 32056
rect 38101 31998 39800 32000
rect 38101 31995 38167 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 38193 30698 38259 30701
rect 39200 30698 39800 30728
rect 38193 30696 39800 30698
rect 38193 30640 38198 30696
rect 38254 30640 39800 30696
rect 38193 30638 39800 30640
rect 38193 30635 38259 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 38193 29338 38259 29341
rect 39200 29338 39800 29368
rect 38193 29336 39800 29338
rect 38193 29280 38198 29336
rect 38254 29280 39800 29336
rect 38193 29278 39800 29280
rect 38193 29275 38259 29278
rect 39200 29248 39800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 38193 28658 38259 28661
rect 39200 28658 39800 28688
rect 38193 28656 39800 28658
rect 38193 28600 38198 28656
rect 38254 28600 39800 28656
rect 38193 28598 39800 28600
rect 38193 28595 38259 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38285 27298 38351 27301
rect 39200 27298 39800 27328
rect 38285 27296 39800 27298
rect 38285 27240 38290 27296
rect 38346 27240 39800 27296
rect 38285 27238 39800 27240
rect 38285 27235 38351 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1761 25938 1827 25941
rect 200 25936 1827 25938
rect 200 25880 1766 25936
rect 1822 25880 1827 25936
rect 200 25878 1827 25880
rect 200 25848 800 25878
rect 1761 25875 1827 25878
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 10869 24170 10935 24173
rect 12341 24170 12407 24173
rect 10869 24168 12407 24170
rect 10869 24112 10874 24168
rect 10930 24112 12346 24168
rect 12402 24112 12407 24168
rect 10869 24110 12407 24112
rect 10869 24107 10935 24110
rect 12341 24107 12407 24110
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 37457 23898 37523 23901
rect 39200 23898 39800 23928
rect 37457 23896 39800 23898
rect 37457 23840 37462 23896
rect 37518 23840 39800 23896
rect 37457 23838 39800 23840
rect 37457 23835 37523 23838
rect 39200 23808 39800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 21398 23020 21404 23084
rect 21468 23082 21474 23084
rect 21633 23082 21699 23085
rect 21468 23080 21699 23082
rect 21468 23024 21638 23080
rect 21694 23024 21699 23080
rect 21468 23022 21699 23024
rect 21468 23020 21474 23022
rect 21633 23019 21699 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1669 22538 1735 22541
rect 200 22536 1735 22538
rect 200 22480 1674 22536
rect 1730 22480 1735 22536
rect 200 22478 1735 22480
rect 200 22448 800 22478
rect 1669 22475 1735 22478
rect 1894 22476 1900 22540
rect 1964 22538 1970 22540
rect 2497 22538 2563 22541
rect 1964 22536 2563 22538
rect 1964 22480 2502 22536
rect 2558 22480 2563 22536
rect 1964 22478 2563 22480
rect 1964 22476 1970 22478
rect 2497 22475 2563 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 10961 21722 11027 21725
rect 14825 21722 14891 21725
rect 10961 21720 14891 21722
rect 10961 21664 10966 21720
rect 11022 21664 14830 21720
rect 14886 21664 14891 21720
rect 10961 21662 14891 21664
rect 10961 21659 11027 21662
rect 14825 21659 14891 21662
rect 13905 21450 13971 21453
rect 18597 21450 18663 21453
rect 13905 21448 18663 21450
rect 13905 21392 13910 21448
rect 13966 21392 18602 21448
rect 18658 21392 18663 21448
rect 13905 21390 18663 21392
rect 13905 21387 13971 21390
rect 18597 21387 18663 21390
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1761 21178 1827 21181
rect 200 21176 1827 21178
rect 200 21120 1766 21176
rect 1822 21120 1827 21176
rect 200 21118 1827 21120
rect 200 21088 800 21118
rect 1761 21115 1827 21118
rect 9673 21042 9739 21045
rect 14733 21042 14799 21045
rect 9673 21040 14799 21042
rect 9673 20984 9678 21040
rect 9734 20984 14738 21040
rect 14794 20984 14799 21040
rect 9673 20982 14799 20984
rect 9673 20979 9739 20982
rect 14733 20979 14799 20982
rect 13721 20906 13787 20909
rect 17585 20906 17651 20909
rect 13721 20904 17651 20906
rect 13721 20848 13726 20904
rect 13782 20848 17590 20904
rect 17646 20848 17651 20904
rect 13721 20846 17651 20848
rect 13721 20843 13787 20846
rect 17585 20843 17651 20846
rect 9673 20770 9739 20773
rect 10869 20770 10935 20773
rect 9673 20768 10935 20770
rect 9673 20712 9678 20768
rect 9734 20712 10874 20768
rect 10930 20712 10935 20768
rect 9673 20710 10935 20712
rect 9673 20707 9739 20710
rect 10869 20707 10935 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 38193 20498 38259 20501
rect 39200 20498 39800 20528
rect 38193 20496 39800 20498
rect 38193 20440 38198 20496
rect 38254 20440 39800 20496
rect 38193 20438 39800 20440
rect 38193 20435 38259 20438
rect 39200 20408 39800 20438
rect 9857 20362 9923 20365
rect 15009 20362 15075 20365
rect 9857 20360 15075 20362
rect 9857 20304 9862 20360
rect 9918 20304 15014 20360
rect 15070 20304 15075 20360
rect 9857 20302 15075 20304
rect 9857 20299 9923 20302
rect 15009 20299 15075 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 12249 20090 12315 20093
rect 17493 20090 17559 20093
rect 12249 20088 17559 20090
rect 12249 20032 12254 20088
rect 12310 20032 17498 20088
rect 17554 20032 17559 20088
rect 12249 20030 17559 20032
rect 12249 20027 12315 20030
rect 17493 20027 17559 20030
rect 7966 19756 7972 19820
rect 8036 19818 8042 19820
rect 9213 19818 9279 19821
rect 8036 19816 9279 19818
rect 8036 19760 9218 19816
rect 9274 19760 9279 19816
rect 8036 19758 9279 19760
rect 8036 19756 8042 19758
rect 9213 19755 9279 19758
rect 14273 19818 14339 19821
rect 18045 19818 18111 19821
rect 14273 19816 18111 19818
rect 14273 19760 14278 19816
rect 14334 19760 18050 19816
rect 18106 19760 18111 19816
rect 14273 19758 18111 19760
rect 14273 19755 14339 19758
rect 18045 19755 18111 19758
rect 9029 19682 9095 19685
rect 9029 19680 9138 19682
rect 9029 19624 9034 19680
rect 9090 19624 9138 19680
rect 9029 19619 9138 19624
rect 9078 19379 9138 19619
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 14641 19546 14707 19549
rect 15561 19546 15627 19549
rect 14641 19544 15627 19546
rect 14641 19488 14646 19544
rect 14702 19488 15566 19544
rect 15622 19488 15627 19544
rect 14641 19486 15627 19488
rect 14641 19483 14707 19486
rect 15561 19483 15627 19486
rect 13721 19412 13787 19413
rect 13670 19410 13676 19412
rect 9078 19374 9187 19379
rect 9078 19318 9126 19374
rect 9182 19318 9187 19374
rect 13630 19350 13676 19410
rect 13740 19408 13787 19412
rect 13782 19352 13787 19408
rect 13670 19348 13676 19350
rect 13740 19348 13787 19352
rect 13721 19347 13787 19348
rect 17493 19412 17559 19413
rect 17493 19408 17540 19412
rect 17604 19410 17610 19412
rect 17493 19352 17498 19408
rect 17493 19348 17540 19352
rect 17604 19350 17650 19410
rect 17604 19348 17610 19350
rect 17493 19347 17559 19348
rect 9078 19316 9187 19318
rect 9121 19313 9187 19316
rect 14549 19274 14615 19277
rect 17217 19274 17283 19277
rect 14549 19272 17283 19274
rect 14549 19216 14554 19272
rect 14610 19216 17222 19272
rect 17278 19216 17283 19272
rect 14549 19214 17283 19216
rect 14549 19211 14615 19214
rect 17217 19211 17283 19214
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 9489 19138 9555 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 9446 19136 9555 19138
rect 9446 19080 9494 19136
rect 9550 19080 9555 19136
rect 9446 19075 9555 19080
rect 11605 19138 11671 19141
rect 16941 19138 17007 19141
rect 11605 19136 17007 19138
rect 11605 19080 11610 19136
rect 11666 19080 16946 19136
rect 17002 19080 17007 19136
rect 11605 19078 17007 19080
rect 11605 19075 11671 19078
rect 16941 19075 17007 19078
rect 38101 19138 38167 19141
rect 39200 19138 39800 19168
rect 38101 19136 39800 19138
rect 38101 19080 38106 19136
rect 38162 19080 39800 19136
rect 38101 19078 39800 19080
rect 38101 19075 38167 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 9446 18869 9506 19075
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 7598 18804 7604 18868
rect 7668 18866 7674 18868
rect 9029 18866 9095 18869
rect 7668 18864 9095 18866
rect 7668 18808 9034 18864
rect 9090 18808 9095 18864
rect 7668 18806 9095 18808
rect 9446 18864 9555 18869
rect 9446 18808 9494 18864
rect 9550 18808 9555 18864
rect 9446 18806 9555 18808
rect 7668 18804 7674 18806
rect 9029 18803 9095 18806
rect 9489 18803 9555 18806
rect 13445 18866 13511 18869
rect 16021 18866 16087 18869
rect 13445 18864 16087 18866
rect 13445 18808 13450 18864
rect 13506 18808 16026 18864
rect 16082 18808 16087 18864
rect 13445 18806 16087 18808
rect 13445 18803 13511 18806
rect 16021 18803 16087 18806
rect 10961 18730 11027 18733
rect 21950 18730 21956 18732
rect 10961 18728 21956 18730
rect 10961 18672 10966 18728
rect 11022 18672 21956 18728
rect 10961 18670 21956 18672
rect 10961 18667 11027 18670
rect 21950 18668 21956 18670
rect 22020 18668 22026 18732
rect 13169 18594 13235 18597
rect 18689 18594 18755 18597
rect 13169 18592 18755 18594
rect 13169 18536 13174 18592
rect 13230 18536 18694 18592
rect 18750 18536 18755 18592
rect 13169 18534 18755 18536
rect 13169 18531 13235 18534
rect 18689 18531 18755 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 10961 18458 11027 18461
rect 13445 18458 13511 18461
rect 16113 18458 16179 18461
rect 10961 18456 16179 18458
rect 10961 18400 10966 18456
rect 11022 18400 13450 18456
rect 13506 18400 16118 18456
rect 16174 18400 16179 18456
rect 10961 18398 16179 18400
rect 10961 18395 11027 18398
rect 13445 18395 13511 18398
rect 16113 18395 16179 18398
rect 39200 18368 39800 18488
rect 14457 18186 14523 18189
rect 17309 18186 17375 18189
rect 14457 18184 17375 18186
rect 14457 18128 14462 18184
rect 14518 18128 17314 18184
rect 17370 18128 17375 18184
rect 14457 18126 17375 18128
rect 14457 18123 14523 18126
rect 17309 18123 17375 18126
rect 6862 17988 6868 18052
rect 6932 18050 6938 18052
rect 8201 18050 8267 18053
rect 6932 18048 8267 18050
rect 6932 17992 8206 18048
rect 8262 17992 8267 18048
rect 6932 17990 8267 17992
rect 6932 17988 6938 17990
rect 8201 17987 8267 17990
rect 11697 18050 11763 18053
rect 11830 18050 11836 18052
rect 11697 18048 11836 18050
rect 11697 17992 11702 18048
rect 11758 17992 11836 18048
rect 11697 17990 11836 17992
rect 11697 17987 11763 17990
rect 11830 17988 11836 17990
rect 11900 17988 11906 18052
rect 12934 17988 12940 18052
rect 13004 18050 13010 18052
rect 18413 18050 18479 18053
rect 13004 18048 18479 18050
rect 13004 17992 18418 18048
rect 18474 17992 18479 18048
rect 13004 17990 18479 17992
rect 13004 17988 13010 17990
rect 18413 17987 18479 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1761 17778 1827 17781
rect 200 17776 1827 17778
rect 200 17720 1766 17776
rect 1822 17720 1827 17776
rect 200 17718 1827 17720
rect 200 17688 800 17718
rect 1761 17715 1827 17718
rect 6637 17778 6703 17781
rect 7557 17778 7623 17781
rect 6637 17776 7623 17778
rect 6637 17720 6642 17776
rect 6698 17720 7562 17776
rect 7618 17720 7623 17776
rect 6637 17718 7623 17720
rect 6637 17715 6703 17718
rect 7557 17715 7623 17718
rect 11973 17778 12039 17781
rect 11973 17776 12266 17778
rect 11973 17720 11978 17776
rect 12034 17720 12266 17776
rect 11973 17718 12266 17720
rect 11973 17715 12039 17718
rect 12206 17644 12266 17718
rect 12198 17580 12204 17644
rect 12268 17642 12274 17644
rect 12341 17642 12407 17645
rect 12268 17640 12407 17642
rect 12268 17584 12346 17640
rect 12402 17584 12407 17640
rect 12268 17582 12407 17584
rect 12268 17580 12274 17582
rect 12341 17579 12407 17582
rect 18454 17580 18460 17644
rect 18524 17642 18530 17644
rect 19517 17642 19583 17645
rect 18524 17640 19583 17642
rect 18524 17584 19522 17640
rect 19578 17584 19583 17640
rect 18524 17582 19583 17584
rect 18524 17580 18530 17582
rect 19517 17579 19583 17582
rect 8477 17506 8543 17509
rect 9029 17506 9095 17509
rect 8477 17504 9095 17506
rect 8477 17448 8482 17504
rect 8538 17448 9034 17504
rect 9090 17448 9095 17504
rect 8477 17446 9095 17448
rect 8477 17443 8543 17446
rect 9029 17443 9095 17446
rect 11789 17506 11855 17509
rect 17585 17506 17651 17509
rect 11789 17504 17651 17506
rect 11789 17448 11794 17504
rect 11850 17448 17590 17504
rect 17646 17448 17651 17504
rect 11789 17446 17651 17448
rect 11789 17443 11855 17446
rect 17585 17443 17651 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 8477 17370 8543 17373
rect 12525 17370 12591 17373
rect 17677 17370 17743 17373
rect 8477 17368 17743 17370
rect 8477 17312 8482 17368
rect 8538 17312 12530 17368
rect 12586 17312 17682 17368
rect 17738 17312 17743 17368
rect 8477 17310 17743 17312
rect 8477 17307 8543 17310
rect 12525 17307 12591 17310
rect 17677 17307 17743 17310
rect 12433 17234 12499 17237
rect 13118 17234 13124 17236
rect 12433 17232 13124 17234
rect 12433 17176 12438 17232
rect 12494 17176 13124 17232
rect 12433 17174 13124 17176
rect 12433 17171 12499 17174
rect 13118 17172 13124 17174
rect 13188 17172 13194 17236
rect 200 17098 800 17128
rect 1577 17098 1643 17101
rect 200 17096 1643 17098
rect 200 17040 1582 17096
rect 1638 17040 1643 17096
rect 200 17038 1643 17040
rect 200 17008 800 17038
rect 1577 17035 1643 17038
rect 4153 17098 4219 17101
rect 5022 17098 5028 17100
rect 4153 17096 5028 17098
rect 4153 17040 4158 17096
rect 4214 17040 5028 17096
rect 4153 17038 5028 17040
rect 4153 17035 4219 17038
rect 5022 17036 5028 17038
rect 5092 17036 5098 17100
rect 10041 17098 10107 17101
rect 10685 17098 10751 17101
rect 10041 17096 10751 17098
rect 10041 17040 10046 17096
rect 10102 17040 10690 17096
rect 10746 17040 10751 17096
rect 10041 17038 10751 17040
rect 10041 17035 10107 17038
rect 10685 17035 10751 17038
rect 16113 17098 16179 17101
rect 24669 17098 24735 17101
rect 16113 17096 24735 17098
rect 16113 17040 16118 17096
rect 16174 17040 24674 17096
rect 24730 17040 24735 17096
rect 16113 17038 24735 17040
rect 16113 17035 16179 17038
rect 24669 17035 24735 17038
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 9397 16826 9463 16829
rect 11053 16826 11119 16829
rect 9397 16824 11119 16826
rect 9397 16768 9402 16824
rect 9458 16768 11058 16824
rect 11114 16768 11119 16824
rect 9397 16766 11119 16768
rect 9397 16763 9463 16766
rect 11053 16763 11119 16766
rect 13261 16826 13327 16829
rect 18413 16826 18479 16829
rect 13261 16824 18479 16826
rect 13261 16768 13266 16824
rect 13322 16768 18418 16824
rect 18474 16768 18479 16824
rect 13261 16766 18479 16768
rect 13261 16763 13327 16766
rect 18413 16763 18479 16766
rect 6545 16692 6611 16693
rect 6494 16690 6500 16692
rect 6454 16630 6500 16690
rect 6564 16688 6611 16692
rect 6606 16632 6611 16688
rect 6494 16628 6500 16630
rect 6564 16628 6611 16632
rect 6545 16627 6611 16628
rect 11145 16690 11211 16693
rect 14457 16692 14523 16693
rect 11278 16690 11284 16692
rect 11145 16688 11284 16690
rect 11145 16632 11150 16688
rect 11206 16632 11284 16688
rect 11145 16630 11284 16632
rect 11145 16627 11211 16630
rect 11278 16628 11284 16630
rect 11348 16628 11354 16692
rect 14406 16690 14412 16692
rect 14366 16630 14412 16690
rect 14476 16688 14523 16692
rect 14518 16632 14523 16688
rect 14406 16628 14412 16630
rect 14476 16628 14523 16632
rect 14457 16627 14523 16628
rect 15653 16692 15719 16693
rect 15653 16688 15700 16692
rect 15764 16690 15770 16692
rect 20529 16690 20595 16693
rect 23974 16690 23980 16692
rect 15653 16632 15658 16688
rect 15653 16628 15700 16632
rect 15764 16630 15810 16690
rect 20529 16688 23980 16690
rect 20529 16632 20534 16688
rect 20590 16632 23980 16688
rect 20529 16630 23980 16632
rect 15764 16628 15770 16630
rect 15653 16627 15719 16628
rect 20529 16627 20595 16630
rect 23974 16628 23980 16630
rect 24044 16628 24050 16692
rect 4654 16492 4660 16556
rect 4724 16554 4730 16556
rect 4889 16554 4955 16557
rect 5257 16556 5323 16557
rect 5206 16554 5212 16556
rect 4724 16552 4955 16554
rect 4724 16496 4894 16552
rect 4950 16496 4955 16552
rect 4724 16494 4955 16496
rect 5166 16494 5212 16554
rect 5276 16552 5323 16556
rect 5318 16496 5323 16552
rect 4724 16492 4730 16494
rect 4889 16491 4955 16494
rect 5206 16492 5212 16494
rect 5276 16492 5323 16496
rect 5257 16491 5323 16492
rect 8201 16554 8267 16557
rect 11145 16554 11211 16557
rect 8201 16552 11211 16554
rect 8201 16496 8206 16552
rect 8262 16496 11150 16552
rect 11206 16496 11211 16552
rect 8201 16494 11211 16496
rect 8201 16491 8267 16494
rect 11145 16491 11211 16494
rect 16941 16554 17007 16557
rect 20897 16554 20963 16557
rect 16941 16552 20963 16554
rect 16941 16496 16946 16552
rect 17002 16496 20902 16552
rect 20958 16496 20963 16552
rect 16941 16494 20963 16496
rect 16941 16491 17007 16494
rect 20897 16491 20963 16494
rect 9397 16418 9463 16421
rect 9857 16418 9923 16421
rect 9397 16416 9923 16418
rect 9397 16360 9402 16416
rect 9458 16360 9862 16416
rect 9918 16360 9923 16416
rect 9397 16358 9923 16360
rect 9397 16355 9463 16358
rect 9857 16355 9923 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 7373 16282 7439 16285
rect 11094 16282 11100 16284
rect 7373 16280 11100 16282
rect 7373 16224 7378 16280
rect 7434 16224 11100 16280
rect 7373 16222 11100 16224
rect 7373 16219 7439 16222
rect 11094 16220 11100 16222
rect 11164 16220 11170 16284
rect 1577 16146 1643 16149
rect 18045 16146 18111 16149
rect 1577 16144 18111 16146
rect 1577 16088 1582 16144
rect 1638 16088 18050 16144
rect 18106 16088 18111 16144
rect 1577 16086 18111 16088
rect 1577 16083 1643 16086
rect 18045 16083 18111 16086
rect 9489 15876 9555 15877
rect 9438 15874 9444 15876
rect 9398 15814 9444 15874
rect 9508 15872 9555 15876
rect 9550 15816 9555 15872
rect 9438 15812 9444 15814
rect 9508 15812 9555 15816
rect 9489 15811 9555 15812
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 8569 15738 8635 15741
rect 10317 15738 10383 15741
rect 8569 15736 10383 15738
rect 8569 15680 8574 15736
rect 8630 15680 10322 15736
rect 10378 15680 10383 15736
rect 8569 15678 10383 15680
rect 8569 15675 8635 15678
rect 10317 15675 10383 15678
rect 38285 15738 38351 15741
rect 39200 15738 39800 15768
rect 38285 15736 39800 15738
rect 38285 15680 38290 15736
rect 38346 15680 39800 15736
rect 38285 15678 39800 15680
rect 38285 15675 38351 15678
rect 39200 15648 39800 15678
rect 3918 15540 3924 15604
rect 3988 15602 3994 15604
rect 8477 15602 8543 15605
rect 3988 15600 8543 15602
rect 3988 15544 8482 15600
rect 8538 15544 8543 15600
rect 3988 15542 8543 15544
rect 3988 15540 3994 15542
rect 8477 15539 8543 15542
rect 7833 15466 7899 15469
rect 12750 15466 12756 15468
rect 7833 15464 12756 15466
rect 7833 15408 7838 15464
rect 7894 15408 12756 15464
rect 7833 15406 12756 15408
rect 7833 15403 7899 15406
rect 12750 15404 12756 15406
rect 12820 15404 12826 15468
rect 20713 15466 20779 15469
rect 23841 15466 23907 15469
rect 20713 15464 23907 15466
rect 20713 15408 20718 15464
rect 20774 15408 23846 15464
rect 23902 15408 23907 15464
rect 20713 15406 23907 15408
rect 20713 15403 20779 15406
rect 23841 15403 23907 15406
rect 2129 15332 2195 15333
rect 2078 15330 2084 15332
rect 2038 15270 2084 15330
rect 2148 15328 2195 15332
rect 2190 15272 2195 15328
rect 2078 15268 2084 15270
rect 2148 15268 2195 15272
rect 2129 15267 2195 15268
rect 4337 15330 4403 15333
rect 5574 15330 5580 15332
rect 4337 15328 5580 15330
rect 4337 15272 4342 15328
rect 4398 15272 5580 15328
rect 4337 15270 5580 15272
rect 4337 15267 4403 15270
rect 5574 15268 5580 15270
rect 5644 15268 5650 15332
rect 6913 15330 6979 15333
rect 8201 15332 8267 15333
rect 7046 15330 7052 15332
rect 6913 15328 7052 15330
rect 6913 15272 6918 15328
rect 6974 15272 7052 15328
rect 6913 15270 7052 15272
rect 6913 15267 6979 15270
rect 7046 15268 7052 15270
rect 7116 15268 7122 15332
rect 8150 15330 8156 15332
rect 8110 15270 8156 15330
rect 8220 15328 8267 15332
rect 8262 15272 8267 15328
rect 8150 15268 8156 15270
rect 8220 15268 8267 15272
rect 9070 15268 9076 15332
rect 9140 15330 9146 15332
rect 9213 15330 9279 15333
rect 9140 15328 9279 15330
rect 9140 15272 9218 15328
rect 9274 15272 9279 15328
rect 9140 15270 9279 15272
rect 9140 15268 9146 15270
rect 8201 15267 8267 15268
rect 9213 15267 9279 15270
rect 11421 15330 11487 15333
rect 13261 15330 13327 15333
rect 17953 15332 18019 15333
rect 17902 15330 17908 15332
rect 11421 15328 13327 15330
rect 11421 15272 11426 15328
rect 11482 15272 13266 15328
rect 13322 15272 13327 15328
rect 11421 15270 13327 15272
rect 17862 15270 17908 15330
rect 17972 15328 18019 15332
rect 18014 15272 18019 15328
rect 11421 15267 11487 15270
rect 13261 15267 13327 15270
rect 17902 15268 17908 15270
rect 17972 15268 18019 15272
rect 18086 15268 18092 15332
rect 18156 15330 18162 15332
rect 18229 15330 18295 15333
rect 18156 15328 18295 15330
rect 18156 15272 18234 15328
rect 18290 15272 18295 15328
rect 18156 15270 18295 15272
rect 18156 15268 18162 15270
rect 17953 15267 18019 15268
rect 18229 15267 18295 15270
rect 20294 15268 20300 15332
rect 20364 15330 20370 15332
rect 23933 15330 23999 15333
rect 20364 15328 23999 15330
rect 20364 15272 23938 15328
rect 23994 15272 23999 15328
rect 20364 15270 23999 15272
rect 20364 15268 20370 15270
rect 23933 15267 23999 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 9765 15194 9831 15197
rect 14549 15194 14615 15197
rect 9765 15192 14615 15194
rect 9765 15136 9770 15192
rect 9826 15136 14554 15192
rect 14610 15136 14615 15192
rect 9765 15134 14615 15136
rect 9765 15131 9831 15134
rect 14549 15131 14615 15134
rect 9213 15058 9279 15061
rect 10869 15058 10935 15061
rect 9213 15056 10935 15058
rect 9213 15000 9218 15056
rect 9274 15000 10874 15056
rect 10930 15000 10935 15056
rect 9213 14998 10935 15000
rect 9213 14995 9279 14998
rect 10869 14995 10935 14998
rect 14641 15058 14707 15061
rect 17493 15058 17559 15061
rect 22185 15058 22251 15061
rect 14641 15056 22251 15058
rect 14641 15000 14646 15056
rect 14702 15000 17498 15056
rect 17554 15000 22190 15056
rect 22246 15000 22251 15056
rect 14641 14998 22251 15000
rect 14641 14995 14707 14998
rect 17493 14995 17559 14998
rect 22185 14995 22251 14998
rect 37181 15058 37247 15061
rect 39200 15058 39800 15088
rect 37181 15056 39800 15058
rect 37181 15000 37186 15056
rect 37242 15000 39800 15056
rect 37181 14998 39800 15000
rect 37181 14995 37247 14998
rect 39200 14968 39800 14998
rect 8477 14922 8543 14925
rect 12985 14922 13051 14925
rect 8477 14920 13051 14922
rect 8477 14864 8482 14920
rect 8538 14864 12990 14920
rect 13046 14864 13051 14920
rect 8477 14862 13051 14864
rect 8477 14859 8543 14862
rect 12985 14859 13051 14862
rect 21909 14922 21975 14925
rect 24209 14922 24275 14925
rect 21909 14920 24275 14922
rect 21909 14864 21914 14920
rect 21970 14864 24214 14920
rect 24270 14864 24275 14920
rect 21909 14862 24275 14864
rect 21909 14859 21975 14862
rect 24209 14859 24275 14862
rect 8293 14786 8359 14789
rect 12566 14786 12572 14788
rect 8293 14784 12572 14786
rect 8293 14728 8298 14784
rect 8354 14728 12572 14784
rect 8293 14726 12572 14728
rect 8293 14723 8359 14726
rect 12566 14724 12572 14726
rect 12636 14724 12642 14788
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4613 14650 4679 14653
rect 4838 14650 4844 14652
rect 4613 14648 4844 14650
rect 4613 14592 4618 14648
rect 4674 14592 4844 14648
rect 4613 14590 4844 14592
rect 4613 14587 4679 14590
rect 4838 14588 4844 14590
rect 4908 14588 4914 14652
rect 8385 14650 8451 14653
rect 9213 14650 9279 14653
rect 8385 14648 9279 14650
rect 8385 14592 8390 14648
rect 8446 14592 9218 14648
rect 9274 14592 9279 14648
rect 8385 14590 9279 14592
rect 8385 14587 8451 14590
rect 9213 14587 9279 14590
rect 10133 14650 10199 14653
rect 13721 14652 13787 14653
rect 10910 14650 10916 14652
rect 10133 14648 10916 14650
rect 10133 14592 10138 14648
rect 10194 14592 10916 14648
rect 10133 14590 10916 14592
rect 10133 14587 10199 14590
rect 10910 14588 10916 14590
rect 10980 14588 10986 14652
rect 13670 14588 13676 14652
rect 13740 14650 13787 14652
rect 13740 14648 13832 14650
rect 13782 14592 13832 14648
rect 13740 14590 13832 14592
rect 13740 14588 13787 14590
rect 13721 14587 13787 14588
rect 8201 14514 8267 14517
rect 11421 14514 11487 14517
rect 8201 14512 11487 14514
rect 8201 14456 8206 14512
rect 8262 14456 11426 14512
rect 11482 14456 11487 14512
rect 8201 14454 11487 14456
rect 8201 14451 8267 14454
rect 11421 14451 11487 14454
rect 20345 14514 20411 14517
rect 23381 14514 23447 14517
rect 20345 14512 23447 14514
rect 20345 14456 20350 14512
rect 20406 14456 23386 14512
rect 23442 14456 23447 14512
rect 20345 14454 23447 14456
rect 20345 14451 20411 14454
rect 23381 14451 23447 14454
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 10225 14378 10291 14381
rect 10358 14378 10364 14380
rect 10225 14376 10364 14378
rect 10225 14320 10230 14376
rect 10286 14320 10364 14376
rect 10225 14318 10364 14320
rect 10225 14315 10291 14318
rect 10358 14316 10364 14318
rect 10428 14316 10434 14380
rect 10501 14378 10567 14381
rect 10685 14378 10751 14381
rect 10501 14376 10751 14378
rect 10501 14320 10506 14376
rect 10562 14320 10690 14376
rect 10746 14320 10751 14376
rect 10501 14318 10751 14320
rect 10501 14315 10567 14318
rect 10685 14315 10751 14318
rect 12709 14378 12775 14381
rect 13721 14378 13787 14381
rect 25957 14378 26023 14381
rect 12709 14376 26023 14378
rect 12709 14320 12714 14376
rect 12770 14320 13726 14376
rect 13782 14320 25962 14376
rect 26018 14320 26023 14376
rect 12709 14318 26023 14320
rect 12709 14315 12775 14318
rect 13721 14315 13787 14318
rect 25957 14315 26023 14318
rect 5809 14242 5875 14245
rect 8334 14242 8340 14244
rect 5809 14240 8340 14242
rect 5809 14184 5814 14240
rect 5870 14184 8340 14240
rect 5809 14182 8340 14184
rect 5809 14179 5875 14182
rect 8334 14180 8340 14182
rect 8404 14180 8410 14244
rect 8477 14242 8543 14245
rect 14457 14242 14523 14245
rect 8477 14240 14523 14242
rect 8477 14184 8482 14240
rect 8538 14184 14462 14240
rect 14518 14184 14523 14240
rect 8477 14182 14523 14184
rect 8477 14179 8543 14182
rect 14457 14179 14523 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 5441 14106 5507 14109
rect 10041 14106 10107 14109
rect 5441 14104 10107 14106
rect 5441 14048 5446 14104
rect 5502 14048 10046 14104
rect 10102 14048 10107 14104
rect 5441 14046 10107 14048
rect 5441 14043 5507 14046
rect 10041 14043 10107 14046
rect 12525 14106 12591 14109
rect 13670 14106 13676 14108
rect 12525 14104 13676 14106
rect 12525 14048 12530 14104
rect 12586 14048 13676 14104
rect 12525 14046 13676 14048
rect 12525 14043 12591 14046
rect 13670 14044 13676 14046
rect 13740 14044 13746 14108
rect 20805 14106 20871 14109
rect 24301 14106 24367 14109
rect 20805 14104 24367 14106
rect 20805 14048 20810 14104
rect 20866 14048 24306 14104
rect 24362 14048 24367 14104
rect 20805 14046 24367 14048
rect 20805 14043 20871 14046
rect 24301 14043 24367 14046
rect 7281 13970 7347 13973
rect 10133 13970 10199 13973
rect 14089 13970 14155 13973
rect 14641 13970 14707 13973
rect 7281 13968 9920 13970
rect 7281 13912 7286 13968
rect 7342 13912 9920 13968
rect 7281 13910 9920 13912
rect 7281 13907 7347 13910
rect 2630 13772 2636 13836
rect 2700 13834 2706 13836
rect 2700 13774 5642 13834
rect 2700 13772 2706 13774
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 5582 13698 5642 13774
rect 6126 13772 6132 13836
rect 6196 13834 6202 13836
rect 8385 13834 8451 13837
rect 6196 13832 8451 13834
rect 6196 13776 8390 13832
rect 8446 13776 8451 13832
rect 6196 13774 8451 13776
rect 6196 13772 6202 13774
rect 8385 13771 8451 13774
rect 9489 13834 9555 13837
rect 9622 13834 9628 13836
rect 9489 13832 9628 13834
rect 9489 13776 9494 13832
rect 9550 13776 9628 13832
rect 9489 13774 9628 13776
rect 9489 13771 9555 13774
rect 9622 13772 9628 13774
rect 9692 13772 9698 13836
rect 9860 13834 9920 13910
rect 10133 13968 14707 13970
rect 10133 13912 10138 13968
rect 10194 13912 14094 13968
rect 14150 13912 14646 13968
rect 14702 13912 14707 13968
rect 10133 13910 14707 13912
rect 10133 13907 10199 13910
rect 14089 13907 14155 13910
rect 14641 13907 14707 13910
rect 17718 13908 17724 13972
rect 17788 13970 17794 13972
rect 21541 13970 21607 13973
rect 17788 13968 21607 13970
rect 17788 13912 21546 13968
rect 21602 13912 21607 13968
rect 17788 13910 21607 13912
rect 17788 13908 17794 13910
rect 21541 13907 21607 13910
rect 21909 13970 21975 13973
rect 27153 13970 27219 13973
rect 21909 13968 27219 13970
rect 21909 13912 21914 13968
rect 21970 13912 27158 13968
rect 27214 13912 27219 13968
rect 21909 13910 27219 13912
rect 21909 13907 21975 13910
rect 27153 13907 27219 13910
rect 18270 13834 18276 13836
rect 9860 13774 18276 13834
rect 18270 13772 18276 13774
rect 18340 13772 18346 13836
rect 19241 13834 19307 13837
rect 23422 13834 23428 13836
rect 19241 13832 23428 13834
rect 19241 13776 19246 13832
rect 19302 13776 23428 13832
rect 19241 13774 23428 13776
rect 19241 13771 19307 13774
rect 23422 13772 23428 13774
rect 23492 13772 23498 13836
rect 6085 13698 6151 13701
rect 5582 13696 6151 13698
rect 5582 13640 6090 13696
rect 6146 13640 6151 13696
rect 5582 13638 6151 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 6085 13635 6151 13638
rect 6545 13698 6611 13701
rect 6862 13698 6868 13700
rect 6545 13696 6868 13698
rect 6545 13640 6550 13696
rect 6606 13640 6868 13696
rect 6545 13638 6868 13640
rect 6545 13635 6611 13638
rect 6862 13636 6868 13638
rect 6932 13636 6938 13700
rect 9121 13698 9187 13701
rect 9254 13698 9260 13700
rect 9121 13696 9260 13698
rect 9121 13640 9126 13696
rect 9182 13640 9260 13696
rect 9121 13638 9260 13640
rect 9121 13635 9187 13638
rect 9254 13636 9260 13638
rect 9324 13636 9330 13700
rect 10174 13636 10180 13700
rect 10244 13698 10250 13700
rect 12198 13698 12204 13700
rect 10244 13638 12204 13698
rect 10244 13636 10250 13638
rect 12198 13636 12204 13638
rect 12268 13636 12274 13700
rect 15377 13698 15443 13701
rect 16757 13698 16823 13701
rect 25957 13698 26023 13701
rect 15377 13696 26023 13698
rect 15377 13640 15382 13696
rect 15438 13640 16762 13696
rect 16818 13640 25962 13696
rect 26018 13640 26023 13696
rect 15377 13638 26023 13640
rect 15377 13635 15443 13638
rect 16757 13635 16823 13638
rect 25957 13635 26023 13638
rect 37181 13698 37247 13701
rect 39200 13698 39800 13728
rect 37181 13696 39800 13698
rect 37181 13640 37186 13696
rect 37242 13640 39800 13696
rect 37181 13638 39800 13640
rect 37181 13635 37247 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 5625 13562 5691 13565
rect 9029 13562 9095 13565
rect 5625 13560 9095 13562
rect 5625 13504 5630 13560
rect 5686 13504 9034 13560
rect 9090 13504 9095 13560
rect 5625 13502 9095 13504
rect 5625 13499 5691 13502
rect 9029 13499 9095 13502
rect 9397 13562 9463 13565
rect 9581 13562 9647 13565
rect 14089 13562 14155 13565
rect 9397 13560 14155 13562
rect 9397 13504 9402 13560
rect 9458 13504 9586 13560
rect 9642 13504 14094 13560
rect 14150 13504 14155 13560
rect 9397 13502 14155 13504
rect 9397 13499 9463 13502
rect 9581 13499 9647 13502
rect 14089 13499 14155 13502
rect 20345 13562 20411 13565
rect 24025 13562 24091 13565
rect 20345 13560 24091 13562
rect 20345 13504 20350 13560
rect 20406 13504 24030 13560
rect 24086 13504 24091 13560
rect 20345 13502 24091 13504
rect 20345 13499 20411 13502
rect 24025 13499 24091 13502
rect 7925 13426 7991 13429
rect 8753 13426 8819 13429
rect 7925 13424 8819 13426
rect 7925 13368 7930 13424
rect 7986 13368 8758 13424
rect 8814 13368 8819 13424
rect 7925 13366 8819 13368
rect 7925 13363 7991 13366
rect 8753 13363 8819 13366
rect 19793 13426 19859 13429
rect 22093 13426 22159 13429
rect 19793 13424 22159 13426
rect 19793 13368 19798 13424
rect 19854 13368 22098 13424
rect 22154 13368 22159 13424
rect 19793 13366 22159 13368
rect 19793 13363 19859 13366
rect 22093 13363 22159 13366
rect 6085 13290 6151 13293
rect 10726 13290 10732 13292
rect 6085 13288 10732 13290
rect 6085 13232 6090 13288
rect 6146 13232 10732 13288
rect 6085 13230 10732 13232
rect 6085 13227 6151 13230
rect 10726 13228 10732 13230
rect 10796 13228 10802 13292
rect 20345 13290 20411 13293
rect 24853 13290 24919 13293
rect 20345 13288 24919 13290
rect 20345 13232 20350 13288
rect 20406 13232 24858 13288
rect 24914 13232 24919 13288
rect 20345 13230 24919 13232
rect 20345 13227 20411 13230
rect 24853 13227 24919 13230
rect 11697 13154 11763 13157
rect 13353 13154 13419 13157
rect 2730 13152 13419 13154
rect 2730 13096 11702 13152
rect 11758 13096 13358 13152
rect 13414 13096 13419 13152
rect 2730 13094 13419 13096
rect 2730 13021 2790 13094
rect 11697 13091 11763 13094
rect 13353 13091 13419 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 2681 13016 2790 13021
rect 2681 12960 2686 13016
rect 2742 12960 2790 13016
rect 2681 12958 2790 12960
rect 10041 13018 10107 13021
rect 12433 13018 12499 13021
rect 17033 13018 17099 13021
rect 10041 13016 12499 13018
rect 10041 12960 10046 13016
rect 10102 12960 12438 13016
rect 12494 12960 12499 13016
rect 10041 12958 12499 12960
rect 2681 12955 2747 12958
rect 10041 12955 10107 12958
rect 12433 12955 12499 12958
rect 13126 13016 17099 13018
rect 13126 12960 17038 13016
rect 17094 12960 17099 13016
rect 13126 12958 17099 12960
rect 9765 12882 9831 12885
rect 13126 12882 13186 12958
rect 17033 12955 17099 12958
rect 9765 12880 13186 12882
rect 9765 12824 9770 12880
rect 9826 12824 13186 12880
rect 9765 12822 13186 12824
rect 13261 12882 13327 12885
rect 20713 12882 20779 12885
rect 13261 12880 20779 12882
rect 13261 12824 13266 12880
rect 13322 12824 20718 12880
rect 20774 12824 20779 12880
rect 13261 12822 20779 12824
rect 9765 12819 9831 12822
rect 13261 12819 13327 12822
rect 20713 12819 20779 12822
rect 4705 12746 4771 12749
rect 5625 12746 5691 12749
rect 4705 12744 5691 12746
rect 4705 12688 4710 12744
rect 4766 12688 5630 12744
rect 5686 12688 5691 12744
rect 4705 12686 5691 12688
rect 4705 12683 4771 12686
rect 5625 12683 5691 12686
rect 11513 12746 11579 12749
rect 17033 12746 17099 12749
rect 11513 12744 17099 12746
rect 11513 12688 11518 12744
rect 11574 12688 17038 12744
rect 17094 12688 17099 12744
rect 11513 12686 17099 12688
rect 11513 12683 11579 12686
rect 17033 12683 17099 12686
rect 4705 12610 4771 12613
rect 6177 12610 6243 12613
rect 4705 12608 6243 12610
rect 4705 12552 4710 12608
rect 4766 12552 6182 12608
rect 6238 12552 6243 12608
rect 4705 12550 6243 12552
rect 4705 12547 4771 12550
rect 6177 12547 6243 12550
rect 10542 12548 10548 12612
rect 10612 12610 10618 12612
rect 10961 12610 11027 12613
rect 10612 12608 11027 12610
rect 10612 12552 10966 12608
rect 11022 12552 11027 12608
rect 10612 12550 11027 12552
rect 10612 12548 10618 12550
rect 10961 12547 11027 12550
rect 11421 12610 11487 12613
rect 12249 12610 12315 12613
rect 11421 12608 12315 12610
rect 11421 12552 11426 12608
rect 11482 12552 12254 12608
rect 12310 12552 12315 12608
rect 11421 12550 12315 12552
rect 11421 12547 11487 12550
rect 12249 12547 12315 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 8385 12474 8451 12477
rect 12157 12474 12223 12477
rect 8385 12472 12223 12474
rect 8385 12416 8390 12472
rect 8446 12416 12162 12472
rect 12218 12416 12223 12472
rect 8385 12414 12223 12416
rect 8385 12411 8451 12414
rect 12157 12411 12223 12414
rect 12382 12412 12388 12476
rect 12452 12474 12458 12476
rect 12750 12474 12756 12476
rect 12452 12414 12756 12474
rect 12452 12412 12458 12414
rect 12750 12412 12756 12414
rect 12820 12412 12826 12476
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 9673 12338 9739 12341
rect 11789 12338 11855 12341
rect 9673 12336 11855 12338
rect 9673 12280 9678 12336
rect 9734 12280 11794 12336
rect 11850 12280 11855 12336
rect 9673 12278 11855 12280
rect 9673 12275 9739 12278
rect 11789 12275 11855 12278
rect 12382 12276 12388 12340
rect 12452 12338 12458 12340
rect 12750 12338 12756 12340
rect 12452 12278 12756 12338
rect 12452 12276 12458 12278
rect 12750 12276 12756 12278
rect 12820 12276 12826 12340
rect 14641 12338 14707 12341
rect 18229 12338 18295 12341
rect 14641 12336 18295 12338
rect 14641 12280 14646 12336
rect 14702 12280 18234 12336
rect 18290 12280 18295 12336
rect 14641 12278 18295 12280
rect 14641 12275 14707 12278
rect 18229 12275 18295 12278
rect 19425 12338 19491 12341
rect 21817 12338 21883 12341
rect 19425 12336 21883 12338
rect 19425 12280 19430 12336
rect 19486 12280 21822 12336
rect 21878 12280 21883 12336
rect 19425 12278 21883 12280
rect 19425 12275 19491 12278
rect 21817 12275 21883 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 5349 12202 5415 12205
rect 6453 12202 6519 12205
rect 5349 12200 6519 12202
rect 5349 12144 5354 12200
rect 5410 12144 6458 12200
rect 6514 12144 6519 12200
rect 5349 12142 6519 12144
rect 5349 12139 5415 12142
rect 6453 12139 6519 12142
rect 7833 12202 7899 12205
rect 11329 12204 11395 12205
rect 7966 12202 7972 12204
rect 7833 12200 7972 12202
rect 7833 12144 7838 12200
rect 7894 12144 7972 12200
rect 7833 12142 7972 12144
rect 7833 12139 7899 12142
rect 7966 12140 7972 12142
rect 8036 12140 8042 12204
rect 11278 12202 11284 12204
rect 11238 12142 11284 12202
rect 11348 12200 11395 12204
rect 15285 12202 15351 12205
rect 21265 12202 21331 12205
rect 11390 12144 11395 12200
rect 11278 12140 11284 12142
rect 11348 12140 11395 12144
rect 11329 12139 11395 12140
rect 12390 12200 15351 12202
rect 12390 12144 15290 12200
rect 15346 12144 15351 12200
rect 12390 12142 15351 12144
rect 11053 12066 11119 12069
rect 12390 12066 12450 12142
rect 15285 12139 15351 12142
rect 16070 12200 21331 12202
rect 16070 12144 21270 12200
rect 21326 12144 21331 12200
rect 16070 12142 21331 12144
rect 11053 12064 12450 12066
rect 11053 12008 11058 12064
rect 11114 12008 12450 12064
rect 11053 12006 12450 12008
rect 14457 12066 14523 12069
rect 16070 12066 16130 12142
rect 21265 12139 21331 12142
rect 14457 12064 16130 12066
rect 14457 12008 14462 12064
rect 14518 12008 16130 12064
rect 14457 12006 16130 12008
rect 11053 12003 11119 12006
rect 14457 12003 14523 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 5257 11930 5323 11933
rect 8109 11930 8175 11933
rect 5257 11928 8175 11930
rect 5257 11872 5262 11928
rect 5318 11872 8114 11928
rect 8170 11872 8175 11928
rect 5257 11870 8175 11872
rect 5257 11867 5323 11870
rect 8109 11867 8175 11870
rect 10409 11930 10475 11933
rect 16389 11930 16455 11933
rect 10409 11928 16455 11930
rect 10409 11872 10414 11928
rect 10470 11872 16394 11928
rect 16450 11872 16455 11928
rect 10409 11870 16455 11872
rect 10409 11867 10475 11870
rect 16389 11867 16455 11870
rect 21081 11930 21147 11933
rect 24393 11930 24459 11933
rect 26969 11930 27035 11933
rect 21081 11928 27035 11930
rect 21081 11872 21086 11928
rect 21142 11872 24398 11928
rect 24454 11872 26974 11928
rect 27030 11872 27035 11928
rect 21081 11870 27035 11872
rect 21081 11867 21147 11870
rect 24393 11867 24459 11870
rect 26969 11867 27035 11870
rect 10726 11732 10732 11796
rect 10796 11794 10802 11796
rect 21081 11794 21147 11797
rect 10796 11792 21147 11794
rect 10796 11736 21086 11792
rect 21142 11736 21147 11792
rect 10796 11734 21147 11736
rect 10796 11732 10802 11734
rect 21081 11731 21147 11734
rect 21265 11794 21331 11797
rect 27429 11794 27495 11797
rect 21265 11792 27495 11794
rect 21265 11736 21270 11792
rect 21326 11736 27434 11792
rect 27490 11736 27495 11792
rect 21265 11734 27495 11736
rect 21265 11731 21331 11734
rect 27429 11731 27495 11734
rect 9029 11658 9095 11661
rect 25221 11658 25287 11661
rect 9029 11656 25287 11658
rect 9029 11600 9034 11656
rect 9090 11600 25226 11656
rect 25282 11600 25287 11656
rect 9029 11598 25287 11600
rect 9029 11595 9095 11598
rect 25221 11595 25287 11598
rect 7782 11460 7788 11524
rect 7852 11522 7858 11524
rect 8017 11522 8083 11525
rect 7852 11520 8083 11522
rect 7852 11464 8022 11520
rect 8078 11464 8083 11520
rect 7852 11462 8083 11464
rect 7852 11460 7858 11462
rect 8017 11459 8083 11462
rect 18873 11522 18939 11525
rect 22093 11522 22159 11525
rect 18873 11520 22159 11522
rect 18873 11464 18878 11520
rect 18934 11464 22098 11520
rect 22154 11464 22159 11520
rect 18873 11462 22159 11464
rect 18873 11459 18939 11462
rect 22093 11459 22159 11462
rect 23105 11522 23171 11525
rect 23473 11522 23539 11525
rect 23105 11520 23539 11522
rect 23105 11464 23110 11520
rect 23166 11464 23478 11520
rect 23534 11464 23539 11520
rect 23105 11462 23539 11464
rect 23105 11459 23171 11462
rect 23473 11459 23539 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 14549 11386 14615 11389
rect 18321 11386 18387 11389
rect 18454 11386 18460 11388
rect 14549 11384 18460 11386
rect 14549 11328 14554 11384
rect 14610 11328 18326 11384
rect 18382 11328 18460 11384
rect 14549 11326 18460 11328
rect 14549 11323 14615 11326
rect 18321 11323 18387 11326
rect 18454 11324 18460 11326
rect 18524 11324 18530 11388
rect 7557 11250 7623 11253
rect 9029 11250 9095 11253
rect 7557 11248 9095 11250
rect 7557 11192 7562 11248
rect 7618 11192 9034 11248
rect 9090 11192 9095 11248
rect 7557 11190 9095 11192
rect 7557 11187 7623 11190
rect 9029 11187 9095 11190
rect 21081 11250 21147 11253
rect 24209 11250 24275 11253
rect 21081 11248 24275 11250
rect 21081 11192 21086 11248
rect 21142 11192 24214 11248
rect 24270 11192 24275 11248
rect 21081 11190 24275 11192
rect 21081 11187 21147 11190
rect 24209 11187 24275 11190
rect 4153 11114 4219 11117
rect 10358 11114 10364 11116
rect 4153 11112 10364 11114
rect 4153 11056 4158 11112
rect 4214 11056 10364 11112
rect 4153 11054 10364 11056
rect 4153 11051 4219 11054
rect 10358 11052 10364 11054
rect 10428 11052 10434 11116
rect 14825 11114 14891 11117
rect 12390 11112 14891 11114
rect 12390 11056 14830 11112
rect 14886 11056 14891 11112
rect 12390 11054 14891 11056
rect 200 10978 800 11008
rect 1577 10978 1643 10981
rect 200 10976 1643 10978
rect 200 10920 1582 10976
rect 1638 10920 1643 10976
rect 200 10918 1643 10920
rect 200 10888 800 10918
rect 1577 10915 1643 10918
rect 4981 10978 5047 10981
rect 5441 10978 5507 10981
rect 9489 10978 9555 10981
rect 12390 10978 12450 11054
rect 14825 11051 14891 11054
rect 21265 11114 21331 11117
rect 22369 11114 22435 11117
rect 21265 11112 22435 11114
rect 21265 11056 21270 11112
rect 21326 11056 22374 11112
rect 22430 11056 22435 11112
rect 21265 11054 22435 11056
rect 21265 11051 21331 11054
rect 22369 11051 22435 11054
rect 23422 11052 23428 11116
rect 23492 11114 23498 11116
rect 27797 11114 27863 11117
rect 23492 11112 27863 11114
rect 23492 11056 27802 11112
rect 27858 11056 27863 11112
rect 23492 11054 27863 11056
rect 23492 11052 23498 11054
rect 27797 11051 27863 11054
rect 4981 10976 12450 10978
rect 4981 10920 4986 10976
rect 5042 10920 5446 10976
rect 5502 10920 9494 10976
rect 9550 10920 12450 10976
rect 4981 10918 12450 10920
rect 13445 10978 13511 10981
rect 14733 10978 14799 10981
rect 13445 10976 14799 10978
rect 13445 10920 13450 10976
rect 13506 10920 14738 10976
rect 14794 10920 14799 10976
rect 13445 10918 14799 10920
rect 4981 10915 5047 10918
rect 5441 10915 5507 10918
rect 9489 10915 9555 10918
rect 13445 10915 13511 10918
rect 14733 10915 14799 10918
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 1577 10842 1643 10845
rect 2630 10842 2636 10844
rect 1577 10840 2636 10842
rect 1577 10784 1582 10840
rect 1638 10784 2636 10840
rect 1577 10782 2636 10784
rect 1577 10779 1643 10782
rect 2630 10780 2636 10782
rect 2700 10780 2706 10844
rect 6729 10842 6795 10845
rect 7465 10842 7531 10845
rect 6729 10840 7531 10842
rect 6729 10784 6734 10840
rect 6790 10784 7470 10840
rect 7526 10784 7531 10840
rect 6729 10782 7531 10784
rect 6729 10779 6795 10782
rect 7465 10779 7531 10782
rect 8661 10842 8727 10845
rect 15009 10842 15075 10845
rect 15929 10842 15995 10845
rect 8661 10840 15995 10842
rect 8661 10784 8666 10840
rect 8722 10784 15014 10840
rect 15070 10784 15934 10840
rect 15990 10784 15995 10840
rect 8661 10782 15995 10784
rect 8661 10779 8727 10782
rect 15009 10779 15075 10782
rect 15929 10779 15995 10782
rect 21173 10706 21239 10709
rect 21398 10706 21404 10708
rect 21173 10704 21404 10706
rect 21173 10648 21178 10704
rect 21234 10648 21404 10704
rect 21173 10646 21404 10648
rect 21173 10643 21239 10646
rect 21398 10644 21404 10646
rect 21468 10644 21474 10708
rect 12985 10570 13051 10573
rect 15193 10570 15259 10573
rect 12985 10568 15259 10570
rect 12985 10512 12990 10568
rect 13046 10512 15198 10568
rect 15254 10512 15259 10568
rect 12985 10510 15259 10512
rect 12985 10507 13051 10510
rect 15193 10507 15259 10510
rect 4705 10436 4771 10437
rect 4654 10372 4660 10436
rect 4724 10434 4771 10436
rect 6729 10434 6795 10437
rect 8201 10434 8267 10437
rect 4724 10432 4816 10434
rect 4766 10376 4816 10432
rect 4724 10374 4816 10376
rect 6729 10432 8267 10434
rect 6729 10376 6734 10432
rect 6790 10376 8206 10432
rect 8262 10376 8267 10432
rect 6729 10374 8267 10376
rect 4724 10372 4771 10374
rect 4705 10371 4771 10372
rect 6729 10371 6795 10374
rect 8201 10371 8267 10374
rect 11697 10434 11763 10437
rect 18086 10434 18092 10436
rect 11697 10432 18092 10434
rect 11697 10376 11702 10432
rect 11758 10376 18092 10432
rect 11697 10374 18092 10376
rect 11697 10371 11763 10374
rect 18086 10372 18092 10374
rect 18156 10372 18162 10436
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1761 10298 1827 10301
rect 200 10296 1827 10298
rect 200 10240 1766 10296
rect 1822 10240 1827 10296
rect 200 10238 1827 10240
rect 200 10208 800 10238
rect 1761 10235 1827 10238
rect 7782 10236 7788 10300
rect 7852 10298 7858 10300
rect 8201 10298 8267 10301
rect 7852 10296 8267 10298
rect 7852 10240 8206 10296
rect 8262 10240 8267 10296
rect 7852 10238 8267 10240
rect 7852 10236 7858 10238
rect 8201 10235 8267 10238
rect 11278 10236 11284 10300
rect 11348 10298 11354 10300
rect 22185 10298 22251 10301
rect 11348 10296 22251 10298
rect 11348 10240 22190 10296
rect 22246 10240 22251 10296
rect 11348 10238 22251 10240
rect 11348 10236 11354 10238
rect 22185 10235 22251 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 4889 10162 4955 10165
rect 8017 10162 8083 10165
rect 4889 10160 8083 10162
rect 4889 10104 4894 10160
rect 4950 10104 8022 10160
rect 8078 10104 8083 10160
rect 4889 10102 8083 10104
rect 4889 10099 4955 10102
rect 8017 10099 8083 10102
rect 10225 10162 10291 10165
rect 15009 10162 15075 10165
rect 10225 10160 15075 10162
rect 10225 10104 10230 10160
rect 10286 10104 15014 10160
rect 15070 10104 15075 10160
rect 10225 10102 15075 10104
rect 10225 10099 10291 10102
rect 15009 10099 15075 10102
rect 13445 10026 13511 10029
rect 20294 10026 20300 10028
rect 13445 10024 20300 10026
rect 13445 9968 13450 10024
rect 13506 9968 20300 10024
rect 13445 9966 20300 9968
rect 13445 9963 13511 9966
rect 20294 9964 20300 9966
rect 20364 9964 20370 10028
rect 9213 9890 9279 9893
rect 10542 9890 10548 9892
rect 9213 9888 10548 9890
rect 9213 9832 9218 9888
rect 9274 9832 10548 9888
rect 9213 9830 10548 9832
rect 9213 9827 9279 9830
rect 10542 9828 10548 9830
rect 10612 9890 10618 9892
rect 15101 9890 15167 9893
rect 10612 9888 15167 9890
rect 10612 9832 15106 9888
rect 15162 9832 15167 9888
rect 10612 9830 15167 9832
rect 10612 9828 10618 9830
rect 15101 9827 15167 9830
rect 24577 9890 24643 9893
rect 29821 9890 29887 9893
rect 24577 9888 29887 9890
rect 24577 9832 24582 9888
rect 24638 9832 29826 9888
rect 29882 9832 29887 9888
rect 24577 9830 29887 9832
rect 24577 9827 24643 9830
rect 29821 9827 29887 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 3918 9692 3924 9756
rect 3988 9754 3994 9756
rect 5257 9754 5323 9757
rect 3988 9752 5323 9754
rect 3988 9696 5262 9752
rect 5318 9696 5323 9752
rect 3988 9694 5323 9696
rect 3988 9692 3994 9694
rect 5257 9691 5323 9694
rect 6913 9754 6979 9757
rect 9121 9756 9187 9757
rect 7598 9754 7604 9756
rect 6913 9752 7604 9754
rect 6913 9696 6918 9752
rect 6974 9696 7604 9752
rect 6913 9694 7604 9696
rect 6913 9691 6979 9694
rect 7598 9692 7604 9694
rect 7668 9692 7674 9756
rect 9070 9754 9076 9756
rect 9030 9694 9076 9754
rect 9140 9752 9187 9756
rect 9182 9696 9187 9752
rect 9070 9692 9076 9694
rect 9140 9692 9187 9696
rect 9121 9691 9187 9692
rect 17309 9754 17375 9757
rect 17902 9754 17908 9756
rect 17309 9752 17908 9754
rect 17309 9696 17314 9752
rect 17370 9696 17908 9752
rect 17309 9694 17908 9696
rect 17309 9691 17375 9694
rect 17902 9692 17908 9694
rect 17972 9692 17978 9756
rect 9305 9618 9371 9621
rect 10225 9618 10291 9621
rect 9305 9616 10291 9618
rect 9305 9560 9310 9616
rect 9366 9560 10230 9616
rect 10286 9560 10291 9616
rect 9305 9558 10291 9560
rect 9305 9555 9371 9558
rect 10225 9555 10291 9558
rect 12566 9556 12572 9620
rect 12636 9618 12642 9620
rect 13537 9618 13603 9621
rect 12636 9616 13603 9618
rect 12636 9560 13542 9616
rect 13598 9560 13603 9616
rect 12636 9558 13603 9560
rect 12636 9556 12642 9558
rect 13537 9555 13603 9558
rect 14958 9556 14964 9620
rect 15028 9618 15034 9620
rect 20713 9618 20779 9621
rect 28809 9618 28875 9621
rect 15028 9558 17418 9618
rect 15028 9556 15034 9558
rect 4981 9482 5047 9485
rect 9438 9482 9444 9484
rect 4981 9480 9444 9482
rect 4981 9424 4986 9480
rect 5042 9424 9444 9480
rect 4981 9422 9444 9424
rect 4981 9419 5047 9422
rect 9438 9420 9444 9422
rect 9508 9482 9514 9484
rect 10961 9482 11027 9485
rect 9508 9480 11027 9482
rect 9508 9424 10966 9480
rect 11022 9424 11027 9480
rect 9508 9422 11027 9424
rect 9508 9420 9514 9422
rect 10961 9419 11027 9422
rect 11973 9482 12039 9485
rect 13118 9482 13124 9484
rect 11973 9480 13124 9482
rect 11973 9424 11978 9480
rect 12034 9424 13124 9480
rect 11973 9422 13124 9424
rect 11973 9419 12039 9422
rect 13118 9420 13124 9422
rect 13188 9482 13194 9484
rect 17125 9482 17191 9485
rect 13188 9480 17191 9482
rect 13188 9424 17130 9480
rect 17186 9424 17191 9480
rect 13188 9422 17191 9424
rect 17358 9482 17418 9558
rect 20713 9616 28875 9618
rect 20713 9560 20718 9616
rect 20774 9560 28814 9616
rect 28870 9560 28875 9616
rect 20713 9558 28875 9560
rect 20713 9555 20779 9558
rect 28809 9555 28875 9558
rect 22553 9482 22619 9485
rect 17358 9480 22619 9482
rect 17358 9424 22558 9480
rect 22614 9424 22619 9480
rect 17358 9422 22619 9424
rect 13188 9420 13194 9422
rect 17125 9419 17191 9422
rect 22553 9419 22619 9422
rect 9397 9346 9463 9349
rect 9765 9346 9831 9349
rect 9397 9344 9831 9346
rect 9397 9288 9402 9344
rect 9458 9288 9770 9344
rect 9826 9288 9831 9344
rect 9397 9286 9831 9288
rect 9397 9283 9463 9286
rect 9765 9283 9831 9286
rect 13261 9346 13327 9349
rect 13813 9346 13879 9349
rect 13261 9344 13879 9346
rect 13261 9288 13266 9344
rect 13322 9288 13818 9344
rect 13874 9288 13879 9344
rect 13261 9286 13879 9288
rect 13261 9283 13327 9286
rect 13813 9283 13879 9286
rect 14825 9346 14891 9349
rect 16297 9346 16363 9349
rect 21449 9346 21515 9349
rect 14825 9344 21515 9346
rect 14825 9288 14830 9344
rect 14886 9288 16302 9344
rect 16358 9288 21454 9344
rect 21510 9288 21515 9344
rect 14825 9286 21515 9288
rect 14825 9283 14891 9286
rect 16297 9283 16363 9286
rect 21449 9283 21515 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4981 9210 5047 9213
rect 5206 9210 5212 9212
rect 4981 9208 5212 9210
rect 4981 9152 4986 9208
rect 5042 9152 5212 9208
rect 4981 9150 5212 9152
rect 4981 9147 5047 9150
rect 5206 9148 5212 9150
rect 5276 9148 5282 9212
rect 16573 9210 16639 9213
rect 17769 9210 17835 9213
rect 25681 9210 25747 9213
rect 16573 9208 25747 9210
rect 16573 9152 16578 9208
rect 16634 9152 17774 9208
rect 17830 9152 25686 9208
rect 25742 9152 25747 9208
rect 16573 9150 25747 9152
rect 16573 9147 16639 9150
rect 17769 9147 17835 9150
rect 25681 9147 25747 9150
rect 9673 9074 9739 9077
rect 9630 9072 9739 9074
rect 9630 9016 9678 9072
rect 9734 9016 9739 9072
rect 9630 9011 9739 9016
rect 10041 9074 10107 9077
rect 18229 9074 18295 9077
rect 10041 9072 18295 9074
rect 10041 9016 10046 9072
rect 10102 9016 18234 9072
rect 18290 9016 18295 9072
rect 10041 9014 18295 9016
rect 10041 9011 10107 9014
rect 18229 9011 18295 9014
rect 19701 9074 19767 9077
rect 21173 9074 21239 9077
rect 19701 9072 21239 9074
rect 19701 9016 19706 9072
rect 19762 9016 21178 9072
rect 21234 9016 21239 9072
rect 19701 9014 21239 9016
rect 19701 9011 19767 9014
rect 21173 9011 21239 9014
rect 21817 9074 21883 9077
rect 23749 9074 23815 9077
rect 21817 9072 23815 9074
rect 21817 9016 21822 9072
rect 21878 9016 23754 9072
rect 23810 9016 23815 9072
rect 21817 9014 23815 9016
rect 21817 9011 21883 9014
rect 23749 9011 23815 9014
rect 200 8938 800 8968
rect 2865 8938 2931 8941
rect 200 8936 2931 8938
rect 200 8880 2870 8936
rect 2926 8880 2931 8936
rect 200 8878 2931 8880
rect 200 8848 800 8878
rect 2865 8875 2931 8878
rect 6494 8876 6500 8940
rect 6564 8938 6570 8940
rect 6821 8938 6887 8941
rect 6564 8936 6887 8938
rect 6564 8880 6826 8936
rect 6882 8880 6887 8936
rect 6564 8878 6887 8880
rect 6564 8876 6570 8878
rect 6821 8875 6887 8878
rect 9630 8938 9690 9011
rect 10409 8938 10475 8941
rect 11881 8938 11947 8941
rect 9630 8936 11947 8938
rect 9630 8880 10414 8936
rect 10470 8880 11886 8936
rect 11942 8880 11947 8936
rect 9630 8878 11947 8880
rect 9630 8669 9690 8878
rect 10409 8875 10475 8878
rect 11881 8875 11947 8878
rect 21817 8938 21883 8941
rect 21950 8938 21956 8940
rect 21817 8936 21956 8938
rect 21817 8880 21822 8936
rect 21878 8880 21956 8936
rect 21817 8878 21956 8880
rect 21817 8875 21883 8878
rect 21950 8876 21956 8878
rect 22020 8938 22026 8940
rect 24894 8938 24900 8940
rect 22020 8878 24900 8938
rect 22020 8876 22026 8878
rect 24894 8876 24900 8878
rect 24964 8876 24970 8940
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 20161 8802 20227 8805
rect 21357 8802 21423 8805
rect 20161 8800 21423 8802
rect 20161 8744 20166 8800
rect 20222 8744 21362 8800
rect 21418 8744 21423 8800
rect 20161 8742 21423 8744
rect 20161 8739 20227 8742
rect 21357 8739 21423 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 9630 8664 9739 8669
rect 20529 8668 20595 8669
rect 9630 8608 9678 8664
rect 9734 8608 9739 8664
rect 9630 8606 9739 8608
rect 9673 8603 9739 8606
rect 20478 8604 20484 8668
rect 20548 8666 20595 8668
rect 23381 8666 23447 8669
rect 25313 8666 25379 8669
rect 20548 8664 20640 8666
rect 20590 8608 20640 8664
rect 20548 8606 20640 8608
rect 23381 8664 25379 8666
rect 23381 8608 23386 8664
rect 23442 8608 25318 8664
rect 25374 8608 25379 8664
rect 23381 8606 25379 8608
rect 20548 8604 20595 8606
rect 20529 8603 20595 8604
rect 23381 8603 23447 8606
rect 25313 8603 25379 8606
rect 8150 8468 8156 8532
rect 8220 8530 8226 8532
rect 8569 8530 8635 8533
rect 8220 8528 8635 8530
rect 8220 8472 8574 8528
rect 8630 8472 8635 8528
rect 8220 8470 8635 8472
rect 8220 8468 8226 8470
rect 8569 8467 8635 8470
rect 15377 8530 15443 8533
rect 26049 8530 26115 8533
rect 15377 8528 26115 8530
rect 15377 8472 15382 8528
rect 15438 8472 26054 8528
rect 26110 8472 26115 8528
rect 15377 8470 26115 8472
rect 15377 8467 15443 8470
rect 26049 8467 26115 8470
rect 2681 8394 2747 8397
rect 24761 8394 24827 8397
rect 2681 8392 24827 8394
rect 2681 8336 2686 8392
rect 2742 8336 24766 8392
rect 24822 8336 24827 8392
rect 2681 8334 24827 8336
rect 2681 8331 2747 8334
rect 24761 8331 24827 8334
rect 1853 8260 1919 8261
rect 1853 8256 1900 8260
rect 1964 8258 1970 8260
rect 1853 8200 1858 8256
rect 1853 8196 1900 8200
rect 1964 8198 2010 8258
rect 1964 8196 1970 8198
rect 5574 8196 5580 8260
rect 5644 8258 5650 8260
rect 9489 8258 9555 8261
rect 11145 8260 11211 8261
rect 11094 8258 11100 8260
rect 5644 8256 9555 8258
rect 5644 8200 9494 8256
rect 9550 8200 9555 8256
rect 5644 8198 9555 8200
rect 11054 8198 11100 8258
rect 11164 8256 11211 8260
rect 11206 8200 11211 8256
rect 5644 8196 5650 8198
rect 1853 8195 1919 8196
rect 9489 8195 9555 8198
rect 11094 8196 11100 8198
rect 11164 8196 11211 8200
rect 11145 8195 11211 8196
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 10685 7986 10751 7989
rect 16481 7986 16547 7989
rect 10685 7984 16547 7986
rect 10685 7928 10690 7984
rect 10746 7928 16486 7984
rect 16542 7928 16547 7984
rect 10685 7926 16547 7928
rect 10685 7923 10751 7926
rect 16481 7923 16547 7926
rect 19885 7850 19951 7853
rect 24485 7850 24551 7853
rect 19885 7848 24551 7850
rect 19885 7792 19890 7848
rect 19946 7792 24490 7848
rect 24546 7792 24551 7848
rect 19885 7790 24551 7792
rect 19885 7787 19951 7790
rect 24485 7787 24551 7790
rect 13261 7714 13327 7717
rect 19149 7714 19215 7717
rect 13261 7712 19215 7714
rect 13261 7656 13266 7712
rect 13322 7656 19154 7712
rect 19210 7656 19215 7712
rect 13261 7654 19215 7656
rect 13261 7651 13327 7654
rect 19149 7651 19215 7654
rect 24761 7714 24827 7717
rect 27061 7714 27127 7717
rect 24761 7712 27127 7714
rect 24761 7656 24766 7712
rect 24822 7656 27066 7712
rect 27122 7656 27127 7712
rect 24761 7654 27127 7656
rect 24761 7651 24827 7654
rect 27061 7651 27127 7654
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 2773 7578 2839 7581
rect 200 7576 2839 7578
rect 200 7520 2778 7576
rect 2834 7520 2839 7576
rect 200 7518 2839 7520
rect 200 7488 800 7518
rect 2773 7515 2839 7518
rect 21081 7578 21147 7581
rect 25865 7578 25931 7581
rect 21081 7576 25931 7578
rect 21081 7520 21086 7576
rect 21142 7520 25870 7576
rect 25926 7520 25931 7576
rect 21081 7518 25931 7520
rect 21081 7515 21147 7518
rect 25865 7515 25931 7518
rect 38193 7578 38259 7581
rect 39200 7578 39800 7608
rect 38193 7576 39800 7578
rect 38193 7520 38198 7576
rect 38254 7520 39800 7576
rect 38193 7518 39800 7520
rect 38193 7515 38259 7518
rect 39200 7488 39800 7518
rect 15009 7442 15075 7445
rect 17718 7442 17724 7444
rect 15009 7440 17724 7442
rect 15009 7384 15014 7440
rect 15070 7384 17724 7440
rect 15009 7382 17724 7384
rect 15009 7379 15075 7382
rect 17718 7380 17724 7382
rect 17788 7380 17794 7444
rect 27153 7442 27219 7445
rect 17910 7440 27219 7442
rect 17910 7384 27158 7440
rect 27214 7384 27219 7440
rect 17910 7382 27219 7384
rect 13261 7306 13327 7309
rect 17910 7306 17970 7382
rect 27153 7379 27219 7382
rect 13261 7304 17970 7306
rect 13261 7248 13266 7304
rect 13322 7248 17970 7304
rect 13261 7246 17970 7248
rect 18689 7306 18755 7309
rect 26693 7306 26759 7309
rect 18689 7304 26759 7306
rect 18689 7248 18694 7304
rect 18750 7248 26698 7304
rect 26754 7248 26759 7304
rect 18689 7246 26759 7248
rect 13261 7243 13327 7246
rect 18689 7243 18755 7246
rect 26693 7243 26759 7246
rect 16481 7170 16547 7173
rect 28809 7170 28875 7173
rect 16481 7168 28875 7170
rect 16481 7112 16486 7168
rect 16542 7112 28814 7168
rect 28870 7112 28875 7168
rect 16481 7110 28875 7112
rect 16481 7107 16547 7110
rect 28809 7107 28875 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 9622 6972 9628 7036
rect 9692 7034 9698 7036
rect 11421 7034 11487 7037
rect 12801 7036 12867 7037
rect 9692 7032 11487 7034
rect 9692 6976 11426 7032
rect 11482 6976 11487 7032
rect 9692 6974 11487 6976
rect 9692 6972 9698 6974
rect 11421 6971 11487 6974
rect 12750 6972 12756 7036
rect 12820 7034 12867 7036
rect 21633 7034 21699 7037
rect 26325 7034 26391 7037
rect 12820 7032 12912 7034
rect 12862 6976 12912 7032
rect 12820 6974 12912 6976
rect 21633 7032 26391 7034
rect 21633 6976 21638 7032
rect 21694 6976 26330 7032
rect 26386 6976 26391 7032
rect 21633 6974 26391 6976
rect 12820 6972 12867 6974
rect 12801 6971 12867 6972
rect 21633 6971 21699 6974
rect 26325 6971 26391 6974
rect 200 6898 800 6928
rect 1577 6898 1643 6901
rect 200 6896 1643 6898
rect 200 6840 1582 6896
rect 1638 6840 1643 6896
rect 200 6838 1643 6840
rect 200 6808 800 6838
rect 1577 6835 1643 6838
rect 4838 6836 4844 6900
rect 4908 6898 4914 6900
rect 8661 6898 8727 6901
rect 4908 6896 8727 6898
rect 4908 6840 8666 6896
rect 8722 6840 8727 6896
rect 4908 6838 8727 6840
rect 4908 6836 4914 6838
rect 8661 6835 8727 6838
rect 10910 6836 10916 6900
rect 10980 6898 10986 6900
rect 11145 6898 11211 6901
rect 10980 6896 11211 6898
rect 10980 6840 11150 6896
rect 11206 6840 11211 6896
rect 10980 6838 11211 6840
rect 10980 6836 10986 6838
rect 11145 6835 11211 6838
rect 11830 6836 11836 6900
rect 11900 6898 11906 6900
rect 12065 6898 12131 6901
rect 11900 6896 12131 6898
rect 11900 6840 12070 6896
rect 12126 6840 12131 6896
rect 11900 6838 12131 6840
rect 11900 6836 11906 6838
rect 12065 6835 12131 6838
rect 18229 6900 18295 6901
rect 18229 6896 18276 6900
rect 18340 6898 18346 6900
rect 19517 6898 19583 6901
rect 20621 6898 20687 6901
rect 22277 6898 22343 6901
rect 18229 6840 18234 6896
rect 18229 6836 18276 6840
rect 18340 6838 18386 6898
rect 19517 6896 22343 6898
rect 19517 6840 19522 6896
rect 19578 6840 20626 6896
rect 20682 6840 22282 6896
rect 22338 6840 22343 6896
rect 19517 6838 22343 6840
rect 18340 6836 18346 6838
rect 18229 6835 18295 6836
rect 19517 6835 19583 6838
rect 20621 6835 20687 6838
rect 22277 6835 22343 6838
rect 24894 6836 24900 6900
rect 24964 6898 24970 6900
rect 25037 6898 25103 6901
rect 24964 6896 25103 6898
rect 24964 6840 25042 6896
rect 25098 6840 25103 6896
rect 24964 6838 25103 6840
rect 24964 6836 24970 6838
rect 25037 6835 25103 6838
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 3877 6762 3943 6765
rect 10174 6762 10180 6764
rect 3877 6760 10180 6762
rect 3877 6704 3882 6760
rect 3938 6704 10180 6760
rect 3877 6702 10180 6704
rect 3877 6699 3943 6702
rect 10174 6700 10180 6702
rect 10244 6700 10250 6764
rect 16665 6762 16731 6765
rect 28993 6762 29059 6765
rect 16665 6760 29059 6762
rect 16665 6704 16670 6760
rect 16726 6704 28998 6760
rect 29054 6704 29059 6760
rect 16665 6702 29059 6704
rect 16665 6699 16731 6702
rect 28993 6699 29059 6702
rect 4521 6626 4587 6629
rect 7373 6626 7439 6629
rect 4521 6624 7439 6626
rect 4521 6568 4526 6624
rect 4582 6568 7378 6624
rect 7434 6568 7439 6624
rect 4521 6566 7439 6568
rect 4521 6563 4587 6566
rect 7373 6563 7439 6566
rect 20345 6626 20411 6629
rect 20478 6626 20484 6628
rect 20345 6624 20484 6626
rect 20345 6568 20350 6624
rect 20406 6568 20484 6624
rect 20345 6566 20484 6568
rect 20345 6563 20411 6566
rect 20478 6564 20484 6566
rect 20548 6626 20554 6628
rect 22185 6626 22251 6629
rect 24945 6626 25011 6629
rect 20548 6624 22251 6626
rect 20548 6568 22190 6624
rect 22246 6568 22251 6624
rect 20548 6566 22251 6568
rect 20548 6564 20554 6566
rect 22185 6563 22251 6566
rect 23062 6624 25011 6626
rect 23062 6568 24950 6624
rect 25006 6568 25011 6624
rect 23062 6566 25011 6568
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 12157 6490 12223 6493
rect 12433 6490 12499 6493
rect 12157 6488 12499 6490
rect 12157 6432 12162 6488
rect 12218 6432 12438 6488
rect 12494 6432 12499 6488
rect 12157 6430 12499 6432
rect 12157 6427 12223 6430
rect 12433 6427 12499 6430
rect 20989 6490 21055 6493
rect 23062 6490 23122 6566
rect 24945 6563 25011 6566
rect 20989 6488 23122 6490
rect 20989 6432 20994 6488
rect 21050 6432 23122 6488
rect 20989 6430 23122 6432
rect 24761 6490 24827 6493
rect 25405 6490 25471 6493
rect 24761 6488 25471 6490
rect 24761 6432 24766 6488
rect 24822 6432 25410 6488
rect 25466 6432 25471 6488
rect 24761 6430 25471 6432
rect 20989 6427 21055 6430
rect 24761 6427 24827 6430
rect 25405 6427 25471 6430
rect 26049 6490 26115 6493
rect 38009 6490 38075 6493
rect 26049 6488 38075 6490
rect 26049 6432 26054 6488
rect 26110 6432 38014 6488
rect 38070 6432 38075 6488
rect 26049 6430 38075 6432
rect 26049 6427 26115 6430
rect 38009 6427 38075 6430
rect 3601 6354 3667 6357
rect 17534 6354 17540 6356
rect 3601 6352 17540 6354
rect 3601 6296 3606 6352
rect 3662 6296 17540 6352
rect 3601 6294 17540 6296
rect 3601 6291 3667 6294
rect 17534 6292 17540 6294
rect 17604 6292 17610 6356
rect 18781 6354 18847 6357
rect 28901 6354 28967 6357
rect 18781 6352 28967 6354
rect 18781 6296 18786 6352
rect 18842 6296 28906 6352
rect 28962 6296 28967 6352
rect 18781 6294 28967 6296
rect 18781 6291 18847 6294
rect 28901 6291 28967 6294
rect 6821 6218 6887 6221
rect 8293 6218 8359 6221
rect 6821 6216 8359 6218
rect 6821 6160 6826 6216
rect 6882 6160 8298 6216
rect 8354 6160 8359 6216
rect 6821 6158 8359 6160
rect 6821 6155 6887 6158
rect 8293 6155 8359 6158
rect 16113 6218 16179 6221
rect 30465 6218 30531 6221
rect 16113 6216 30531 6218
rect 16113 6160 16118 6216
rect 16174 6160 30470 6216
rect 30526 6160 30531 6216
rect 16113 6158 30531 6160
rect 16113 6155 16179 6158
rect 30465 6155 30531 6158
rect 18965 6082 19031 6085
rect 21817 6082 21883 6085
rect 18965 6080 21883 6082
rect 18965 6024 18970 6080
rect 19026 6024 21822 6080
rect 21878 6024 21883 6080
rect 18965 6022 21883 6024
rect 18965 6019 19031 6022
rect 21817 6019 21883 6022
rect 23013 6082 23079 6085
rect 30649 6082 30715 6085
rect 23013 6080 30715 6082
rect 23013 6024 23018 6080
rect 23074 6024 30654 6080
rect 30710 6024 30715 6080
rect 23013 6022 30715 6024
rect 23013 6019 23079 6022
rect 30649 6019 30715 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 6729 5946 6795 5949
rect 8845 5946 8911 5949
rect 6729 5944 8911 5946
rect 6729 5888 6734 5944
rect 6790 5888 8850 5944
rect 8906 5888 8911 5944
rect 6729 5886 8911 5888
rect 6729 5883 6795 5886
rect 8845 5883 8911 5886
rect 15837 5946 15903 5949
rect 21081 5946 21147 5949
rect 15837 5944 21147 5946
rect 15837 5888 15842 5944
rect 15898 5888 21086 5944
rect 21142 5888 21147 5944
rect 15837 5886 21147 5888
rect 15837 5883 15903 5886
rect 21081 5883 21147 5886
rect 23841 5946 23907 5949
rect 25681 5946 25747 5949
rect 26785 5946 26851 5949
rect 23841 5944 26851 5946
rect 23841 5888 23846 5944
rect 23902 5888 25686 5944
rect 25742 5888 26790 5944
rect 26846 5888 26851 5944
rect 23841 5886 26851 5888
rect 23841 5883 23907 5886
rect 25681 5883 25747 5886
rect 26785 5883 26851 5886
rect 6269 5810 6335 5813
rect 7281 5810 7347 5813
rect 6269 5808 7347 5810
rect 6269 5752 6274 5808
rect 6330 5752 7286 5808
rect 7342 5752 7347 5808
rect 6269 5750 7347 5752
rect 6269 5747 6335 5750
rect 7281 5747 7347 5750
rect 17493 5810 17559 5813
rect 30649 5810 30715 5813
rect 17493 5808 30715 5810
rect 17493 5752 17498 5808
rect 17554 5752 30654 5808
rect 30710 5752 30715 5808
rect 17493 5750 30715 5752
rect 17493 5747 17559 5750
rect 30649 5747 30715 5750
rect 6821 5674 6887 5677
rect 7046 5674 7052 5676
rect 6821 5672 7052 5674
rect 6821 5616 6826 5672
rect 6882 5616 7052 5672
rect 6821 5614 7052 5616
rect 6821 5611 6887 5614
rect 7046 5612 7052 5614
rect 7116 5674 7122 5676
rect 8201 5674 8267 5677
rect 7116 5672 8267 5674
rect 7116 5616 8206 5672
rect 8262 5616 8267 5672
rect 7116 5614 8267 5616
rect 7116 5612 7122 5614
rect 8201 5611 8267 5614
rect 9254 5612 9260 5676
rect 9324 5674 9330 5676
rect 13721 5674 13787 5677
rect 9324 5672 13787 5674
rect 9324 5616 13726 5672
rect 13782 5616 13787 5672
rect 9324 5614 13787 5616
rect 9324 5612 9330 5614
rect 13721 5611 13787 5614
rect 20069 5674 20135 5677
rect 23749 5674 23815 5677
rect 20069 5672 23815 5674
rect 20069 5616 20074 5672
rect 20130 5616 23754 5672
rect 23810 5616 23815 5672
rect 20069 5614 23815 5616
rect 20069 5611 20135 5614
rect 23749 5611 23815 5614
rect 24393 5674 24459 5677
rect 27797 5674 27863 5677
rect 24393 5672 27863 5674
rect 24393 5616 24398 5672
rect 24454 5616 27802 5672
rect 27858 5616 27863 5672
rect 24393 5614 27863 5616
rect 24393 5611 24459 5614
rect 27797 5611 27863 5614
rect 200 5538 800 5568
rect 2957 5538 3023 5541
rect 200 5536 3023 5538
rect 200 5480 2962 5536
rect 3018 5480 3023 5536
rect 200 5478 3023 5480
rect 200 5448 800 5478
rect 2957 5475 3023 5478
rect 8569 5538 8635 5541
rect 14406 5538 14412 5540
rect 8569 5536 14412 5538
rect 8569 5480 8574 5536
rect 8630 5480 14412 5536
rect 8569 5478 14412 5480
rect 8569 5475 8635 5478
rect 14406 5476 14412 5478
rect 14476 5476 14482 5540
rect 19977 5538 20043 5541
rect 27245 5538 27311 5541
rect 19977 5536 27311 5538
rect 19977 5480 19982 5536
rect 20038 5480 27250 5536
rect 27306 5480 27311 5536
rect 19977 5478 27311 5480
rect 19977 5475 20043 5478
rect 27245 5475 27311 5478
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 14641 5402 14707 5405
rect 18137 5402 18203 5405
rect 14641 5400 18203 5402
rect 14641 5344 14646 5400
rect 14702 5344 18142 5400
rect 18198 5344 18203 5400
rect 14641 5342 18203 5344
rect 14641 5339 14707 5342
rect 18137 5339 18203 5342
rect 22093 5402 22159 5405
rect 22553 5402 22619 5405
rect 22093 5400 22619 5402
rect 22093 5344 22098 5400
rect 22154 5344 22558 5400
rect 22614 5344 22619 5400
rect 22093 5342 22619 5344
rect 22093 5339 22159 5342
rect 22553 5339 22619 5342
rect 24669 5402 24735 5405
rect 35617 5402 35683 5405
rect 24669 5400 35683 5402
rect 24669 5344 24674 5400
rect 24730 5344 35622 5400
rect 35678 5344 35683 5400
rect 24669 5342 35683 5344
rect 24669 5339 24735 5342
rect 35617 5339 35683 5342
rect 13997 5266 14063 5269
rect 20345 5266 20411 5269
rect 13997 5264 20411 5266
rect 13997 5208 14002 5264
rect 14058 5208 20350 5264
rect 20406 5208 20411 5264
rect 13997 5206 20411 5208
rect 13997 5203 14063 5206
rect 20345 5203 20411 5206
rect 17861 5130 17927 5133
rect 21357 5130 21423 5133
rect 17861 5128 21423 5130
rect 17861 5072 17866 5128
rect 17922 5072 21362 5128
rect 21418 5072 21423 5128
rect 17861 5070 21423 5072
rect 17861 5067 17927 5070
rect 21357 5067 21423 5070
rect 25037 5130 25103 5133
rect 28809 5130 28875 5133
rect 25037 5128 28875 5130
rect 25037 5072 25042 5128
rect 25098 5072 28814 5128
rect 28870 5072 28875 5128
rect 25037 5070 28875 5072
rect 25037 5067 25103 5070
rect 28809 5067 28875 5070
rect 19425 4994 19491 4997
rect 21449 4994 21515 4997
rect 19425 4992 21515 4994
rect 19425 4936 19430 4992
rect 19486 4936 21454 4992
rect 21510 4936 21515 4992
rect 19425 4934 21515 4936
rect 19425 4931 19491 4934
rect 21449 4931 21515 4934
rect 22645 4994 22711 4997
rect 23749 4994 23815 4997
rect 31293 4994 31359 4997
rect 22645 4992 31359 4994
rect 22645 4936 22650 4992
rect 22706 4936 23754 4992
rect 23810 4936 31298 4992
rect 31354 4936 31359 4992
rect 22645 4934 31359 4936
rect 22645 4931 22711 4934
rect 23749 4931 23815 4934
rect 31293 4931 31359 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 5533 4858 5599 4861
rect 15694 4858 15700 4860
rect 5533 4856 15700 4858
rect 5533 4800 5538 4856
rect 5594 4800 15700 4856
rect 5533 4798 15700 4800
rect 5533 4795 5599 4798
rect 15694 4796 15700 4798
rect 15764 4796 15770 4860
rect 26325 4858 26391 4861
rect 29729 4858 29795 4861
rect 26325 4856 29795 4858
rect 26325 4800 26330 4856
rect 26386 4800 29734 4856
rect 29790 4800 29795 4856
rect 26325 4798 29795 4800
rect 26325 4795 26391 4798
rect 29729 4795 29795 4798
rect 4521 4722 4587 4725
rect 6085 4722 6151 4725
rect 4521 4720 6151 4722
rect 4521 4664 4526 4720
rect 4582 4664 6090 4720
rect 6146 4664 6151 4720
rect 4521 4662 6151 4664
rect 4521 4659 4587 4662
rect 6085 4659 6151 4662
rect 11881 4722 11947 4725
rect 13813 4722 13879 4725
rect 11881 4720 13879 4722
rect 11881 4664 11886 4720
rect 11942 4664 13818 4720
rect 13874 4664 13879 4720
rect 11881 4662 13879 4664
rect 11881 4659 11947 4662
rect 13813 4659 13879 4662
rect 14273 4722 14339 4725
rect 33593 4722 33659 4725
rect 14273 4720 33659 4722
rect 14273 4664 14278 4720
rect 14334 4664 33598 4720
rect 33654 4664 33659 4720
rect 14273 4662 33659 4664
rect 14273 4659 14339 4662
rect 33593 4659 33659 4662
rect 10041 4586 10107 4589
rect 12934 4586 12940 4588
rect 10041 4584 12940 4586
rect 10041 4528 10046 4584
rect 10102 4528 12940 4584
rect 10041 4526 12940 4528
rect 10041 4523 10107 4526
rect 12934 4524 12940 4526
rect 13004 4524 13010 4588
rect 21081 4586 21147 4589
rect 31109 4586 31175 4589
rect 21081 4584 31175 4586
rect 21081 4528 21086 4584
rect 21142 4528 31114 4584
rect 31170 4528 31175 4584
rect 21081 4526 31175 4528
rect 21081 4523 21147 4526
rect 31109 4523 31175 4526
rect 23289 4450 23355 4453
rect 26233 4450 26299 4453
rect 23289 4448 26299 4450
rect 23289 4392 23294 4448
rect 23350 4392 26238 4448
rect 26294 4392 26299 4448
rect 23289 4390 26299 4392
rect 23289 4387 23355 4390
rect 26233 4387 26299 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4521 4314 4587 4317
rect 8753 4314 8819 4317
rect 4521 4312 8819 4314
rect 4521 4256 4526 4312
rect 4582 4256 8758 4312
rect 8814 4256 8819 4312
rect 4521 4254 8819 4256
rect 4521 4251 4587 4254
rect 8753 4251 8819 4254
rect 24761 4314 24827 4317
rect 30373 4314 30439 4317
rect 24761 4312 30439 4314
rect 24761 4256 24766 4312
rect 24822 4256 30378 4312
rect 30434 4256 30439 4312
rect 24761 4254 30439 4256
rect 24761 4251 24827 4254
rect 30373 4251 30439 4254
rect 200 4178 800 4208
rect 2773 4178 2839 4181
rect 200 4176 2839 4178
rect 200 4120 2778 4176
rect 2834 4120 2839 4176
rect 200 4118 2839 4120
rect 200 4088 800 4118
rect 2773 4115 2839 4118
rect 10961 4178 11027 4181
rect 32857 4178 32923 4181
rect 10961 4176 32923 4178
rect 10961 4120 10966 4176
rect 11022 4120 32862 4176
rect 32918 4120 32923 4176
rect 10961 4118 32923 4120
rect 10961 4115 11027 4118
rect 32857 4115 32923 4118
rect 38193 4178 38259 4181
rect 39200 4178 39800 4208
rect 38193 4176 39800 4178
rect 38193 4120 38198 4176
rect 38254 4120 39800 4176
rect 38193 4118 39800 4120
rect 38193 4115 38259 4118
rect 39200 4088 39800 4118
rect 3785 4042 3851 4045
rect 8293 4044 8359 4045
rect 6126 4042 6132 4044
rect 3785 4040 6132 4042
rect 3785 3984 3790 4040
rect 3846 3984 6132 4040
rect 3785 3982 6132 3984
rect 3785 3979 3851 3982
rect 6126 3980 6132 3982
rect 6196 3980 6202 4044
rect 8293 4042 8340 4044
rect 8248 4040 8340 4042
rect 8404 4042 8410 4044
rect 11053 4042 11119 4045
rect 8404 4040 11119 4042
rect 8248 3984 8298 4040
rect 8404 3984 11058 4040
rect 11114 3984 11119 4040
rect 8248 3982 8340 3984
rect 8293 3980 8340 3982
rect 8404 3982 11119 3984
rect 8404 3980 8410 3982
rect 8293 3979 8359 3980
rect 11053 3979 11119 3982
rect 25589 4042 25655 4045
rect 30741 4042 30807 4045
rect 25589 4040 30807 4042
rect 25589 3984 25594 4040
rect 25650 3984 30746 4040
rect 30802 3984 30807 4040
rect 25589 3982 30807 3984
rect 25589 3979 25655 3982
rect 30741 3979 30807 3982
rect 12801 3906 12867 3909
rect 16573 3906 16639 3909
rect 12801 3904 16639 3906
rect 12801 3848 12806 3904
rect 12862 3848 16578 3904
rect 16634 3848 16639 3904
rect 12801 3846 16639 3848
rect 12801 3843 12867 3846
rect 16573 3843 16639 3846
rect 22277 3906 22343 3909
rect 32949 3906 33015 3909
rect 22277 3904 33015 3906
rect 22277 3848 22282 3904
rect 22338 3848 32954 3904
rect 33010 3848 33015 3904
rect 22277 3846 33015 3848
rect 22277 3843 22343 3846
rect 32949 3843 33015 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 10685 3770 10751 3773
rect 12709 3770 12775 3773
rect 10685 3768 12775 3770
rect 10685 3712 10690 3768
rect 10746 3712 12714 3768
rect 12770 3712 12775 3768
rect 10685 3710 12775 3712
rect 10685 3707 10751 3710
rect 12709 3707 12775 3710
rect 24485 3770 24551 3773
rect 28809 3770 28875 3773
rect 24485 3768 28875 3770
rect 24485 3712 24490 3768
rect 24546 3712 28814 3768
rect 28870 3712 28875 3768
rect 24485 3710 28875 3712
rect 24485 3707 24551 3710
rect 28809 3707 28875 3710
rect 2037 3636 2103 3637
rect 2037 3634 2084 3636
rect 1992 3632 2084 3634
rect 1992 3576 2042 3632
rect 1992 3574 2084 3576
rect 2037 3572 2084 3574
rect 2148 3572 2154 3636
rect 11053 3634 11119 3637
rect 5030 3632 11119 3634
rect 5030 3576 11058 3632
rect 11114 3576 11119 3632
rect 5030 3574 11119 3576
rect 2037 3571 2103 3572
rect 200 3498 800 3528
rect 2865 3498 2931 3501
rect 200 3496 2931 3498
rect 200 3440 2870 3496
rect 2926 3440 2931 3496
rect 200 3438 2931 3440
rect 200 3408 800 3438
rect 2865 3435 2931 3438
rect 4889 3498 4955 3501
rect 5030 3500 5090 3574
rect 11053 3571 11119 3574
rect 12525 3634 12591 3637
rect 13077 3634 13143 3637
rect 12525 3632 13143 3634
rect 12525 3576 12530 3632
rect 12586 3576 13082 3632
rect 13138 3576 13143 3632
rect 12525 3574 13143 3576
rect 12525 3571 12591 3574
rect 13077 3571 13143 3574
rect 16573 3634 16639 3637
rect 20621 3634 20687 3637
rect 16573 3632 20687 3634
rect 16573 3576 16578 3632
rect 16634 3576 20626 3632
rect 20682 3576 20687 3632
rect 16573 3574 20687 3576
rect 16573 3571 16639 3574
rect 20621 3571 20687 3574
rect 24669 3634 24735 3637
rect 32489 3634 32555 3637
rect 24669 3632 32555 3634
rect 24669 3576 24674 3632
rect 24730 3576 32494 3632
rect 32550 3576 32555 3632
rect 24669 3574 32555 3576
rect 24669 3571 24735 3574
rect 32489 3571 32555 3574
rect 5022 3498 5028 3500
rect 4889 3496 5028 3498
rect 4889 3440 4894 3496
rect 4950 3440 5028 3496
rect 4889 3438 5028 3440
rect 4889 3435 4955 3438
rect 5022 3436 5028 3438
rect 5092 3436 5098 3500
rect 9121 3498 9187 3501
rect 25405 3498 25471 3501
rect 9121 3496 25471 3498
rect 9121 3440 9126 3496
rect 9182 3440 25410 3496
rect 25466 3440 25471 3496
rect 9121 3438 25471 3440
rect 9121 3435 9187 3438
rect 25405 3435 25471 3438
rect 25957 3498 26023 3501
rect 26877 3498 26943 3501
rect 25957 3496 26943 3498
rect 25957 3440 25962 3496
rect 26018 3440 26882 3496
rect 26938 3440 26943 3496
rect 25957 3438 26943 3440
rect 25957 3435 26023 3438
rect 26877 3435 26943 3438
rect 38285 3498 38351 3501
rect 39200 3498 39800 3528
rect 38285 3496 39800 3498
rect 38285 3440 38290 3496
rect 38346 3440 39800 3496
rect 38285 3438 39800 3440
rect 38285 3435 38351 3438
rect 39200 3408 39800 3438
rect 2037 3362 2103 3365
rect 21541 3362 21607 3365
rect 24853 3362 24919 3365
rect 27613 3362 27679 3365
rect 2037 3360 2790 3362
rect 2037 3304 2042 3360
rect 2098 3304 2790 3360
rect 2037 3302 2790 3304
rect 2037 3299 2103 3302
rect 2730 3226 2790 3302
rect 21541 3360 24594 3362
rect 21541 3304 21546 3360
rect 21602 3304 24594 3360
rect 21541 3302 24594 3304
rect 21541 3299 21607 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 8569 3226 8635 3229
rect 23933 3228 23999 3229
rect 11278 3226 11284 3228
rect 2730 3224 11284 3226
rect 2730 3168 8574 3224
rect 8630 3168 11284 3224
rect 2730 3166 11284 3168
rect 8569 3163 8635 3166
rect 11278 3164 11284 3166
rect 11348 3164 11354 3228
rect 23933 3226 23980 3228
rect 23888 3224 23980 3226
rect 23888 3168 23938 3224
rect 23888 3166 23980 3168
rect 23933 3164 23980 3166
rect 24044 3164 24050 3228
rect 23933 3163 23999 3164
rect 6821 3090 6887 3093
rect 24393 3090 24459 3093
rect 6821 3088 24459 3090
rect 6821 3032 6826 3088
rect 6882 3032 24398 3088
rect 24454 3032 24459 3088
rect 6821 3030 24459 3032
rect 24534 3090 24594 3302
rect 24853 3360 27679 3362
rect 24853 3304 24858 3360
rect 24914 3304 27618 3360
rect 27674 3304 27679 3360
rect 24853 3302 27679 3304
rect 24853 3299 24919 3302
rect 27613 3299 27679 3302
rect 25497 3226 25563 3229
rect 26325 3226 26391 3229
rect 25497 3224 26391 3226
rect 25497 3168 25502 3224
rect 25558 3168 26330 3224
rect 26386 3168 26391 3224
rect 25497 3166 26391 3168
rect 25497 3163 25563 3166
rect 26325 3163 26391 3166
rect 27245 3226 27311 3229
rect 33593 3226 33659 3229
rect 27245 3224 33659 3226
rect 27245 3168 27250 3224
rect 27306 3168 33598 3224
rect 33654 3168 33659 3224
rect 27245 3166 33659 3168
rect 27245 3163 27311 3166
rect 33593 3163 33659 3166
rect 28901 3090 28967 3093
rect 24534 3088 28967 3090
rect 24534 3032 28906 3088
rect 28962 3032 28967 3088
rect 24534 3030 28967 3032
rect 6821 3027 6887 3030
rect 24393 3027 24459 3030
rect 28901 3027 28967 3030
rect 5257 2954 5323 2957
rect 7465 2954 7531 2957
rect 5257 2952 7531 2954
rect 5257 2896 5262 2952
rect 5318 2896 7470 2952
rect 7526 2896 7531 2952
rect 5257 2894 7531 2896
rect 5257 2891 5323 2894
rect 7465 2891 7531 2894
rect 22369 2954 22435 2957
rect 29729 2954 29795 2957
rect 22369 2952 29795 2954
rect 22369 2896 22374 2952
rect 22430 2896 29734 2952
rect 29790 2896 29795 2952
rect 22369 2894 29795 2896
rect 22369 2891 22435 2894
rect 29729 2891 29795 2894
rect 11605 2818 11671 2821
rect 12617 2818 12683 2821
rect 11605 2816 12683 2818
rect 11605 2760 11610 2816
rect 11666 2760 12622 2816
rect 12678 2760 12683 2816
rect 11605 2758 12683 2760
rect 11605 2755 11671 2758
rect 12617 2755 12683 2758
rect 16481 2818 16547 2821
rect 26693 2818 26759 2821
rect 16481 2816 26759 2818
rect 16481 2760 16486 2816
rect 16542 2760 26698 2816
rect 26754 2760 26759 2816
rect 16481 2758 26759 2760
rect 16481 2755 16547 2758
rect 26693 2755 26759 2758
rect 27061 2818 27127 2821
rect 34697 2818 34763 2821
rect 27061 2816 34763 2818
rect 27061 2760 27066 2816
rect 27122 2760 34702 2816
rect 34758 2760 34763 2816
rect 27061 2758 34763 2760
rect 27061 2755 27127 2758
rect 34697 2755 34763 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19885 2682 19951 2685
rect 24853 2682 24919 2685
rect 19885 2680 24919 2682
rect 19885 2624 19890 2680
rect 19946 2624 24858 2680
rect 24914 2624 24919 2680
rect 19885 2622 24919 2624
rect 19885 2619 19951 2622
rect 24853 2619 24919 2622
rect 25037 2682 25103 2685
rect 28993 2682 29059 2685
rect 25037 2680 29059 2682
rect 25037 2624 25042 2680
rect 25098 2624 28998 2680
rect 29054 2624 29059 2680
rect 25037 2622 29059 2624
rect 25037 2619 25103 2622
rect 28993 2619 29059 2622
rect 13721 2546 13787 2549
rect 30465 2546 30531 2549
rect 13721 2544 30531 2546
rect 13721 2488 13726 2544
rect 13782 2488 30470 2544
rect 30526 2488 30531 2544
rect 13721 2486 30531 2488
rect 13721 2483 13787 2486
rect 30465 2483 30531 2486
rect 5901 2410 5967 2413
rect 27245 2410 27311 2413
rect 5901 2408 27311 2410
rect 5901 2352 5906 2408
rect 5962 2352 27250 2408
rect 27306 2352 27311 2408
rect 5901 2350 27311 2352
rect 5901 2347 5967 2350
rect 27245 2347 27311 2350
rect 25313 2274 25379 2277
rect 35525 2274 35591 2277
rect 25313 2272 35591 2274
rect 25313 2216 25318 2272
rect 25374 2216 35530 2272
rect 35586 2216 35591 2272
rect 25313 2214 35591 2216
rect 25313 2211 25379 2214
rect 35525 2211 35591 2214
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 2773 2138 2839 2141
rect 200 2136 2839 2138
rect 200 2080 2778 2136
rect 2834 2080 2839 2136
rect 200 2078 2839 2080
rect 200 2048 800 2078
rect 2773 2075 2839 2078
rect 38193 2138 38259 2141
rect 39200 2138 39800 2168
rect 38193 2136 39800 2138
rect 38193 2080 38198 2136
rect 38254 2080 39800 2136
rect 38193 2078 39800 2080
rect 38193 2075 38259 2078
rect 39200 2048 39800 2078
rect 13537 2002 13603 2005
rect 30557 2002 30623 2005
rect 13537 2000 30623 2002
rect 13537 1944 13542 2000
rect 13598 1944 30562 2000
rect 30618 1944 30623 2000
rect 13537 1942 30623 1944
rect 13537 1939 13603 1942
rect 30557 1939 30623 1942
rect 13721 1866 13787 1869
rect 28073 1866 28139 1869
rect 13721 1864 28139 1866
rect 13721 1808 13726 1864
rect 13782 1808 28078 1864
rect 28134 1808 28139 1864
rect 13721 1806 28139 1808
rect 13721 1803 13787 1806
rect 28073 1803 28139 1806
rect 3969 1730 4035 1733
rect 26509 1730 26575 1733
rect 3969 1728 26575 1730
rect 3969 1672 3974 1728
rect 4030 1672 26514 1728
rect 26570 1672 26575 1728
rect 3969 1670 26575 1672
rect 3969 1667 4035 1670
rect 26509 1667 26575 1670
rect 37457 1458 37523 1461
rect 37457 1456 39314 1458
rect 37457 1400 37462 1456
rect 37518 1400 39314 1456
rect 37457 1398 39314 1400
rect 37457 1395 37523 1398
rect 39254 1050 39314 1398
rect 39070 990 39314 1050
rect 3325 914 3391 917
rect 1902 912 3391 914
rect 1902 856 3330 912
rect 3386 856 3391 912
rect 1902 854 3391 856
rect 200 778 800 808
rect 1902 778 1962 854
rect 3325 851 3391 854
rect 200 718 1962 778
rect 39070 778 39130 990
rect 39200 778 39800 808
rect 39070 718 39800 778
rect 200 688 800 718
rect 39200 688 39800 718
rect 37181 98 37247 101
rect 39200 98 39800 128
rect 37181 96 39800 98
rect 37181 40 37186 96
rect 37242 40 39800 96
rect 37181 38 39800 40
rect 37181 35 37247 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 14964 37224 15028 37228
rect 14964 37168 14978 37224
rect 14978 37168 15028 37224
rect 14964 37164 15028 37168
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 21404 23020 21468 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 1900 22476 1964 22540
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 7972 19756 8036 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 13676 19408 13740 19412
rect 13676 19352 13726 19408
rect 13726 19352 13740 19408
rect 13676 19348 13740 19352
rect 17540 19408 17604 19412
rect 17540 19352 17554 19408
rect 17554 19352 17604 19408
rect 17540 19348 17604 19352
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 7604 18804 7668 18868
rect 21956 18668 22020 18732
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 6868 17988 6932 18052
rect 11836 17988 11900 18052
rect 12940 17988 13004 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 12204 17580 12268 17644
rect 18460 17580 18524 17644
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 13124 17172 13188 17236
rect 5028 17036 5092 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 6500 16688 6564 16692
rect 6500 16632 6550 16688
rect 6550 16632 6564 16688
rect 6500 16628 6564 16632
rect 11284 16628 11348 16692
rect 14412 16688 14476 16692
rect 14412 16632 14462 16688
rect 14462 16632 14476 16688
rect 14412 16628 14476 16632
rect 15700 16688 15764 16692
rect 15700 16632 15714 16688
rect 15714 16632 15764 16688
rect 15700 16628 15764 16632
rect 23980 16628 24044 16692
rect 4660 16492 4724 16556
rect 5212 16552 5276 16556
rect 5212 16496 5262 16552
rect 5262 16496 5276 16552
rect 5212 16492 5276 16496
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 11100 16220 11164 16284
rect 9444 15872 9508 15876
rect 9444 15816 9494 15872
rect 9494 15816 9508 15872
rect 9444 15812 9508 15816
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 3924 15540 3988 15604
rect 12756 15404 12820 15468
rect 2084 15328 2148 15332
rect 2084 15272 2134 15328
rect 2134 15272 2148 15328
rect 2084 15268 2148 15272
rect 5580 15268 5644 15332
rect 7052 15268 7116 15332
rect 8156 15328 8220 15332
rect 8156 15272 8206 15328
rect 8206 15272 8220 15328
rect 8156 15268 8220 15272
rect 9076 15268 9140 15332
rect 17908 15328 17972 15332
rect 17908 15272 17958 15328
rect 17958 15272 17972 15328
rect 17908 15268 17972 15272
rect 18092 15268 18156 15332
rect 20300 15268 20364 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 12572 14724 12636 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4844 14588 4908 14652
rect 10916 14588 10980 14652
rect 13676 14648 13740 14652
rect 13676 14592 13726 14648
rect 13726 14592 13740 14648
rect 13676 14588 13740 14592
rect 10364 14316 10428 14380
rect 8340 14180 8404 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 13676 14044 13740 14108
rect 2636 13772 2700 13836
rect 6132 13772 6196 13836
rect 9628 13772 9692 13836
rect 17724 13908 17788 13972
rect 18276 13772 18340 13836
rect 23428 13772 23492 13836
rect 6868 13636 6932 13700
rect 9260 13636 9324 13700
rect 10180 13636 10244 13700
rect 12204 13636 12268 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 10732 13228 10796 13292
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 10548 12548 10612 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 12388 12412 12452 12476
rect 12756 12412 12820 12476
rect 12388 12276 12452 12340
rect 12756 12276 12820 12340
rect 7972 12140 8036 12204
rect 11284 12200 11348 12204
rect 11284 12144 11334 12200
rect 11334 12144 11348 12200
rect 11284 12140 11348 12144
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 10732 11732 10796 11796
rect 7788 11460 7852 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 18460 11324 18524 11388
rect 10364 11052 10428 11116
rect 23428 11052 23492 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 2636 10780 2700 10844
rect 21404 10644 21468 10708
rect 4660 10432 4724 10436
rect 4660 10376 4710 10432
rect 4710 10376 4724 10432
rect 4660 10372 4724 10376
rect 18092 10372 18156 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 7788 10236 7852 10300
rect 11284 10236 11348 10300
rect 20300 9964 20364 10028
rect 10548 9828 10612 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 3924 9692 3988 9756
rect 7604 9692 7668 9756
rect 9076 9752 9140 9756
rect 9076 9696 9126 9752
rect 9126 9696 9140 9752
rect 9076 9692 9140 9696
rect 17908 9692 17972 9756
rect 12572 9556 12636 9620
rect 14964 9556 15028 9620
rect 9444 9420 9508 9484
rect 13124 9420 13188 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 5212 9148 5276 9212
rect 6500 8876 6564 8940
rect 21956 8876 22020 8940
rect 24900 8876 24964 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 20484 8664 20548 8668
rect 20484 8608 20534 8664
rect 20534 8608 20548 8664
rect 20484 8604 20548 8608
rect 8156 8468 8220 8532
rect 1900 8256 1964 8260
rect 1900 8200 1914 8256
rect 1914 8200 1964 8256
rect 1900 8196 1964 8200
rect 5580 8196 5644 8260
rect 11100 8256 11164 8260
rect 11100 8200 11150 8256
rect 11150 8200 11164 8256
rect 11100 8196 11164 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 17724 7380 17788 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 9628 6972 9692 7036
rect 12756 7032 12820 7036
rect 12756 6976 12806 7032
rect 12806 6976 12820 7032
rect 12756 6972 12820 6976
rect 4844 6836 4908 6900
rect 10916 6836 10980 6900
rect 11836 6836 11900 6900
rect 18276 6896 18340 6900
rect 18276 6840 18290 6896
rect 18290 6840 18340 6896
rect 18276 6836 18340 6840
rect 24900 6836 24964 6900
rect 10180 6700 10244 6764
rect 20484 6564 20548 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 17540 6292 17604 6356
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 7052 5612 7116 5676
rect 9260 5612 9324 5676
rect 14412 5476 14476 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 15700 4796 15764 4860
rect 12940 4524 13004 4588
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 6132 3980 6196 4044
rect 8340 4040 8404 4044
rect 8340 3984 8354 4040
rect 8354 3984 8404 4040
rect 8340 3980 8404 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 2084 3632 2148 3636
rect 2084 3576 2098 3632
rect 2098 3576 2148 3632
rect 2084 3572 2148 3576
rect 5028 3436 5092 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 11284 3164 11348 3228
rect 23980 3224 24044 3228
rect 23980 3168 23994 3224
rect 23994 3168 24044 3224
rect 23980 3164 24044 3168
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 14963 37228 15029 37229
rect 14963 37164 14964 37228
rect 15028 37164 15029 37228
rect 14963 37163 15029 37164
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 1899 22540 1965 22541
rect 1899 22476 1900 22540
rect 1964 22476 1965 22540
rect 1899 22475 1965 22476
rect 1902 8261 1962 22475
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 7971 19820 8037 19821
rect 7971 19756 7972 19820
rect 8036 19756 8037 19820
rect 7971 19755 8037 19756
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 7603 18868 7669 18869
rect 7603 18804 7604 18868
rect 7668 18804 7669 18868
rect 7603 18803 7669 18804
rect 6867 18052 6933 18053
rect 6867 17988 6868 18052
rect 6932 17988 6933 18052
rect 6867 17987 6933 17988
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 5027 17100 5093 17101
rect 5027 17036 5028 17100
rect 5092 17036 5093 17100
rect 5027 17035 5093 17036
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4659 16556 4725 16557
rect 4659 16492 4660 16556
rect 4724 16492 4725 16556
rect 4659 16491 4725 16492
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 3923 15604 3989 15605
rect 3923 15540 3924 15604
rect 3988 15540 3989 15604
rect 3923 15539 3989 15540
rect 2083 15332 2149 15333
rect 2083 15268 2084 15332
rect 2148 15268 2149 15332
rect 2083 15267 2149 15268
rect 1899 8260 1965 8261
rect 1899 8196 1900 8260
rect 1964 8196 1965 8260
rect 1899 8195 1965 8196
rect 2086 3637 2146 15267
rect 2635 13836 2701 13837
rect 2635 13772 2636 13836
rect 2700 13772 2701 13836
rect 2635 13771 2701 13772
rect 2638 10845 2698 13771
rect 2635 10844 2701 10845
rect 2635 10780 2636 10844
rect 2700 10780 2701 10844
rect 2635 10779 2701 10780
rect 3926 9757 3986 15539
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4662 10437 4722 16491
rect 4843 14652 4909 14653
rect 4843 14588 4844 14652
rect 4908 14588 4909 14652
rect 4843 14587 4909 14588
rect 4659 10436 4725 10437
rect 4659 10372 4660 10436
rect 4724 10372 4725 10436
rect 4659 10371 4725 10372
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3923 9756 3989 9757
rect 3923 9692 3924 9756
rect 3988 9692 3989 9756
rect 3923 9691 3989 9692
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4846 6901 4906 14587
rect 4843 6900 4909 6901
rect 4843 6836 4844 6900
rect 4908 6836 4909 6900
rect 4843 6835 4909 6836
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 2083 3636 2149 3637
rect 2083 3572 2084 3636
rect 2148 3572 2149 3636
rect 2083 3571 2149 3572
rect 4208 2752 4528 3776
rect 5030 3501 5090 17035
rect 6499 16692 6565 16693
rect 6499 16628 6500 16692
rect 6564 16628 6565 16692
rect 6499 16627 6565 16628
rect 5211 16556 5277 16557
rect 5211 16492 5212 16556
rect 5276 16492 5277 16556
rect 5211 16491 5277 16492
rect 5214 9213 5274 16491
rect 5579 15332 5645 15333
rect 5579 15268 5580 15332
rect 5644 15268 5645 15332
rect 5579 15267 5645 15268
rect 5211 9212 5277 9213
rect 5211 9148 5212 9212
rect 5276 9148 5277 9212
rect 5211 9147 5277 9148
rect 5582 8261 5642 15267
rect 6131 13836 6197 13837
rect 6131 13772 6132 13836
rect 6196 13772 6197 13836
rect 6131 13771 6197 13772
rect 5579 8260 5645 8261
rect 5579 8196 5580 8260
rect 5644 8196 5645 8260
rect 5579 8195 5645 8196
rect 6134 4045 6194 13771
rect 6502 8941 6562 16627
rect 6870 13701 6930 17987
rect 7051 15332 7117 15333
rect 7051 15268 7052 15332
rect 7116 15268 7117 15332
rect 7051 15267 7117 15268
rect 6867 13700 6933 13701
rect 6867 13636 6868 13700
rect 6932 13636 6933 13700
rect 6867 13635 6933 13636
rect 6499 8940 6565 8941
rect 6499 8876 6500 8940
rect 6564 8876 6565 8940
rect 6499 8875 6565 8876
rect 7054 5677 7114 15267
rect 7606 9757 7666 18803
rect 7974 12205 8034 19755
rect 13675 19412 13741 19413
rect 13675 19348 13676 19412
rect 13740 19348 13741 19412
rect 13675 19347 13741 19348
rect 11835 18052 11901 18053
rect 11835 17988 11836 18052
rect 11900 17988 11901 18052
rect 11835 17987 11901 17988
rect 12939 18052 13005 18053
rect 12939 17988 12940 18052
rect 13004 17988 13005 18052
rect 12939 17987 13005 17988
rect 11283 16692 11349 16693
rect 11283 16628 11284 16692
rect 11348 16628 11349 16692
rect 11283 16627 11349 16628
rect 11099 16284 11165 16285
rect 11099 16220 11100 16284
rect 11164 16220 11165 16284
rect 11099 16219 11165 16220
rect 9443 15876 9509 15877
rect 9443 15812 9444 15876
rect 9508 15812 9509 15876
rect 9443 15811 9509 15812
rect 8155 15332 8221 15333
rect 8155 15268 8156 15332
rect 8220 15268 8221 15332
rect 8155 15267 8221 15268
rect 9075 15332 9141 15333
rect 9075 15268 9076 15332
rect 9140 15268 9141 15332
rect 9075 15267 9141 15268
rect 7971 12204 8037 12205
rect 7971 12140 7972 12204
rect 8036 12140 8037 12204
rect 7971 12139 8037 12140
rect 7787 11524 7853 11525
rect 7787 11460 7788 11524
rect 7852 11460 7853 11524
rect 7787 11459 7853 11460
rect 7790 10301 7850 11459
rect 7787 10300 7853 10301
rect 7787 10236 7788 10300
rect 7852 10236 7853 10300
rect 7787 10235 7853 10236
rect 7603 9756 7669 9757
rect 7603 9692 7604 9756
rect 7668 9692 7669 9756
rect 7603 9691 7669 9692
rect 8158 8533 8218 15267
rect 8339 14244 8405 14245
rect 8339 14180 8340 14244
rect 8404 14180 8405 14244
rect 8339 14179 8405 14180
rect 8155 8532 8221 8533
rect 8155 8468 8156 8532
rect 8220 8468 8221 8532
rect 8155 8467 8221 8468
rect 7051 5676 7117 5677
rect 7051 5612 7052 5676
rect 7116 5612 7117 5676
rect 7051 5611 7117 5612
rect 8342 4045 8402 14179
rect 9078 9757 9138 15267
rect 9259 13700 9325 13701
rect 9259 13636 9260 13700
rect 9324 13636 9325 13700
rect 9259 13635 9325 13636
rect 9075 9756 9141 9757
rect 9075 9692 9076 9756
rect 9140 9692 9141 9756
rect 9075 9691 9141 9692
rect 9262 5677 9322 13635
rect 9446 9485 9506 15811
rect 10915 14652 10981 14653
rect 10915 14588 10916 14652
rect 10980 14588 10981 14652
rect 10915 14587 10981 14588
rect 10363 14380 10429 14381
rect 10363 14316 10364 14380
rect 10428 14316 10429 14380
rect 10363 14315 10429 14316
rect 9627 13836 9693 13837
rect 9627 13772 9628 13836
rect 9692 13772 9693 13836
rect 9627 13771 9693 13772
rect 9443 9484 9509 9485
rect 9443 9420 9444 9484
rect 9508 9420 9509 9484
rect 9443 9419 9509 9420
rect 9630 7037 9690 13771
rect 10179 13700 10245 13701
rect 10179 13636 10180 13700
rect 10244 13636 10245 13700
rect 10179 13635 10245 13636
rect 9627 7036 9693 7037
rect 9627 6972 9628 7036
rect 9692 6972 9693 7036
rect 9627 6971 9693 6972
rect 10182 6765 10242 13635
rect 10366 11117 10426 14315
rect 10731 13292 10797 13293
rect 10731 13228 10732 13292
rect 10796 13228 10797 13292
rect 10731 13227 10797 13228
rect 10547 12612 10613 12613
rect 10547 12548 10548 12612
rect 10612 12548 10613 12612
rect 10547 12547 10613 12548
rect 10363 11116 10429 11117
rect 10363 11052 10364 11116
rect 10428 11052 10429 11116
rect 10363 11051 10429 11052
rect 10550 9893 10610 12547
rect 10734 11797 10794 13227
rect 10731 11796 10797 11797
rect 10731 11732 10732 11796
rect 10796 11732 10797 11796
rect 10731 11731 10797 11732
rect 10547 9892 10613 9893
rect 10547 9828 10548 9892
rect 10612 9828 10613 9892
rect 10547 9827 10613 9828
rect 10918 6901 10978 14587
rect 11102 8261 11162 16219
rect 11286 12205 11346 16627
rect 11283 12204 11349 12205
rect 11283 12140 11284 12204
rect 11348 12140 11349 12204
rect 11283 12139 11349 12140
rect 11283 10300 11349 10301
rect 11283 10236 11284 10300
rect 11348 10236 11349 10300
rect 11283 10235 11349 10236
rect 11099 8260 11165 8261
rect 11099 8196 11100 8260
rect 11164 8196 11165 8260
rect 11099 8195 11165 8196
rect 10915 6900 10981 6901
rect 10915 6836 10916 6900
rect 10980 6836 10981 6900
rect 10915 6835 10981 6836
rect 10179 6764 10245 6765
rect 10179 6700 10180 6764
rect 10244 6700 10245 6764
rect 10179 6699 10245 6700
rect 9259 5676 9325 5677
rect 9259 5612 9260 5676
rect 9324 5612 9325 5676
rect 9259 5611 9325 5612
rect 6131 4044 6197 4045
rect 6131 3980 6132 4044
rect 6196 3980 6197 4044
rect 6131 3979 6197 3980
rect 8339 4044 8405 4045
rect 8339 3980 8340 4044
rect 8404 3980 8405 4044
rect 8339 3979 8405 3980
rect 5027 3500 5093 3501
rect 5027 3436 5028 3500
rect 5092 3436 5093 3500
rect 5027 3435 5093 3436
rect 11286 3229 11346 10235
rect 11838 6901 11898 17987
rect 12203 17644 12269 17645
rect 12203 17580 12204 17644
rect 12268 17580 12269 17644
rect 12203 17579 12269 17580
rect 12206 13701 12266 17579
rect 12755 15468 12821 15469
rect 12755 15404 12756 15468
rect 12820 15404 12821 15468
rect 12755 15403 12821 15404
rect 12571 14788 12637 14789
rect 12571 14724 12572 14788
rect 12636 14724 12637 14788
rect 12571 14723 12637 14724
rect 12203 13700 12269 13701
rect 12203 13636 12204 13700
rect 12268 13636 12269 13700
rect 12203 13635 12269 13636
rect 12387 12476 12453 12477
rect 12387 12412 12388 12476
rect 12452 12412 12453 12476
rect 12387 12411 12453 12412
rect 12390 12341 12450 12411
rect 12387 12340 12453 12341
rect 12387 12276 12388 12340
rect 12452 12276 12453 12340
rect 12387 12275 12453 12276
rect 12574 9621 12634 14723
rect 12758 12477 12818 15403
rect 12755 12476 12821 12477
rect 12755 12412 12756 12476
rect 12820 12412 12821 12476
rect 12755 12411 12821 12412
rect 12755 12340 12821 12341
rect 12755 12276 12756 12340
rect 12820 12276 12821 12340
rect 12755 12275 12821 12276
rect 12571 9620 12637 9621
rect 12571 9556 12572 9620
rect 12636 9556 12637 9620
rect 12571 9555 12637 9556
rect 12758 7037 12818 12275
rect 12755 7036 12821 7037
rect 12755 6972 12756 7036
rect 12820 6972 12821 7036
rect 12755 6971 12821 6972
rect 11835 6900 11901 6901
rect 11835 6836 11836 6900
rect 11900 6836 11901 6900
rect 11835 6835 11901 6836
rect 12942 4589 13002 17987
rect 13123 17236 13189 17237
rect 13123 17172 13124 17236
rect 13188 17172 13189 17236
rect 13123 17171 13189 17172
rect 13126 9485 13186 17171
rect 13678 14653 13738 19347
rect 14411 16692 14477 16693
rect 14411 16628 14412 16692
rect 14476 16628 14477 16692
rect 14411 16627 14477 16628
rect 13675 14652 13741 14653
rect 13675 14588 13676 14652
rect 13740 14588 13741 14652
rect 13675 14587 13741 14588
rect 13678 14109 13738 14587
rect 13675 14108 13741 14109
rect 13675 14044 13676 14108
rect 13740 14044 13741 14108
rect 13675 14043 13741 14044
rect 13123 9484 13189 9485
rect 13123 9420 13124 9484
rect 13188 9420 13189 9484
rect 13123 9419 13189 9420
rect 14414 5541 14474 16627
rect 14966 9621 15026 37163
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 21403 23084 21469 23085
rect 21403 23020 21404 23084
rect 21468 23020 21469 23084
rect 21403 23019 21469 23020
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 15699 16692 15765 16693
rect 15699 16628 15700 16692
rect 15764 16628 15765 16692
rect 15699 16627 15765 16628
rect 14963 9620 15029 9621
rect 14963 9556 14964 9620
rect 15028 9556 15029 9620
rect 14963 9555 15029 9556
rect 14411 5540 14477 5541
rect 14411 5476 14412 5540
rect 14476 5476 14477 5540
rect 14411 5475 14477 5476
rect 15702 4861 15762 16627
rect 17542 6357 17602 19347
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 18459 17644 18525 17645
rect 18459 17580 18460 17644
rect 18524 17580 18525 17644
rect 18459 17579 18525 17580
rect 17907 15332 17973 15333
rect 17907 15268 17908 15332
rect 17972 15268 17973 15332
rect 17907 15267 17973 15268
rect 18091 15332 18157 15333
rect 18091 15268 18092 15332
rect 18156 15268 18157 15332
rect 18091 15267 18157 15268
rect 17723 13972 17789 13973
rect 17723 13908 17724 13972
rect 17788 13908 17789 13972
rect 17723 13907 17789 13908
rect 17726 7445 17786 13907
rect 17910 9757 17970 15267
rect 18094 10437 18154 15267
rect 18275 13836 18341 13837
rect 18275 13772 18276 13836
rect 18340 13772 18341 13836
rect 18275 13771 18341 13772
rect 18091 10436 18157 10437
rect 18091 10372 18092 10436
rect 18156 10372 18157 10436
rect 18091 10371 18157 10372
rect 17907 9756 17973 9757
rect 17907 9692 17908 9756
rect 17972 9692 17973 9756
rect 17907 9691 17973 9692
rect 17723 7444 17789 7445
rect 17723 7380 17724 7444
rect 17788 7380 17789 7444
rect 17723 7379 17789 7380
rect 18278 6901 18338 13771
rect 18462 11389 18522 17579
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 20299 15332 20365 15333
rect 20299 15268 20300 15332
rect 20364 15268 20365 15332
rect 20299 15267 20365 15268
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 18459 11388 18525 11389
rect 18459 11324 18460 11388
rect 18524 11324 18525 11388
rect 18459 11323 18525 11324
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 20302 10029 20362 15267
rect 21406 10709 21466 23019
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 21955 18732 22021 18733
rect 21955 18668 21956 18732
rect 22020 18668 22021 18732
rect 21955 18667 22021 18668
rect 21403 10708 21469 10709
rect 21403 10644 21404 10708
rect 21468 10644 21469 10708
rect 21403 10643 21469 10644
rect 20299 10028 20365 10029
rect 20299 9964 20300 10028
rect 20364 9964 20365 10028
rect 20299 9963 20365 9964
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 21958 8941 22018 18667
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 23979 16692 24045 16693
rect 23979 16628 23980 16692
rect 24044 16628 24045 16692
rect 23979 16627 24045 16628
rect 23427 13836 23493 13837
rect 23427 13772 23428 13836
rect 23492 13772 23493 13836
rect 23427 13771 23493 13772
rect 23430 11117 23490 13771
rect 23427 11116 23493 11117
rect 23427 11052 23428 11116
rect 23492 11052 23493 11116
rect 23427 11051 23493 11052
rect 21955 8940 22021 8941
rect 21955 8876 21956 8940
rect 22020 8876 22021 8940
rect 21955 8875 22021 8876
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 20483 8668 20549 8669
rect 20483 8604 20484 8668
rect 20548 8604 20549 8668
rect 20483 8603 20549 8604
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 18275 6900 18341 6901
rect 18275 6836 18276 6900
rect 18340 6836 18341 6900
rect 18275 6835 18341 6836
rect 19568 6560 19888 7584
rect 20486 6629 20546 8603
rect 20483 6628 20549 6629
rect 20483 6564 20484 6628
rect 20548 6564 20549 6628
rect 20483 6563 20549 6564
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 17539 6356 17605 6357
rect 17539 6292 17540 6356
rect 17604 6292 17605 6356
rect 17539 6291 17605 6292
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 15699 4860 15765 4861
rect 15699 4796 15700 4860
rect 15764 4796 15765 4860
rect 15699 4795 15765 4796
rect 12939 4588 13005 4589
rect 12939 4524 12940 4588
rect 13004 4524 13005 4588
rect 12939 4523 13005 4524
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 11283 3228 11349 3229
rect 11283 3164 11284 3228
rect 11348 3164 11349 3228
rect 11283 3163 11349 3164
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 23982 3229 24042 16627
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 24899 8940 24965 8941
rect 24899 8876 24900 8940
rect 24964 8876 24965 8940
rect 24899 8875 24965 8876
rect 24902 6901 24962 8875
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 24899 6900 24965 6901
rect 24899 6836 24900 6900
rect 24964 6836 24965 6900
rect 24899 6835 24965 6836
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 23979 3228 24045 3229
rect 23979 3164 23980 3228
rect 24044 3164 24045 3228
rect 23979 3163 24045 3164
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1667941163
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1667941163
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1667941163
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1667941163
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1667941163
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1667941163
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1667941163
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1667941163
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1667941163
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1667941163
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1667941163
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1667941163
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1667941163
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1667941163
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1667941163
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_82
timestamp 1667941163
transform 1 0 8648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1667941163
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1667941163
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1667941163
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_194
timestamp 1667941163
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1667941163
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_229
timestamp 1667941163
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1667941163
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1667941163
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_257
timestamp 1667941163
transform 1 0 24748 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1667941163
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1667941163
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1667941163
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_313
timestamp 1667941163
transform 1 0 29900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_320
timestamp 1667941163
transform 1 0 30544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_327
timestamp 1667941163
transform 1 0 31188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1667941163
transform 1 0 32568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1667941163
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1667941163
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1667941163
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1667941163
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_384
timestamp 1667941163
transform 1 0 36432 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1667941163
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1667941163
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1667941163
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_156
timestamp 1667941163
transform 1 0 15456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1667941163
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_220
timestamp 1667941163
transform 1 0 21344 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_228
timestamp 1667941163
transform 1 0 22080 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_234
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1667941163
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_268
timestamp 1667941163
transform 1 0 25760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1667941163
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_282
timestamp 1667941163
transform 1 0 27048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_290
timestamp 1667941163
transform 1 0 27784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1667941163
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1667941163
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_314
timestamp 1667941163
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1667941163
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1667941163
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_342
timestamp 1667941163
transform 1 0 32568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_349
timestamp 1667941163
transform 1 0 33212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1667941163
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_370
timestamp 1667941163
transform 1 0 35144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_385
timestamp 1667941163
transform 1 0 36524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_390
timestamp 1667941163
transform 1 0 36984 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_398
timestamp 1667941163
transform 1 0 37720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_26
timestamp 1667941163
transform 1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1667941163
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_80
timestamp 1667941163
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1667941163
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_138
timestamp 1667941163
transform 1 0 13800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1667941163
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1667941163
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1667941163
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1667941163
transform 1 0 24656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1667941163
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_267
timestamp 1667941163
transform 1 0 25668 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_271
timestamp 1667941163
transform 1 0 26036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1667941163
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1667941163
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1667941163
transform 1 0 28704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1667941163
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_314
timestamp 1667941163
transform 1 0 29992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_321
timestamp 1667941163
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1667941163
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1667941163
transform 1 0 32568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_356
timestamp 1667941163
transform 1 0 33856 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_363 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_375
timestamp 1667941163
transform 1 0 35604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1667941163
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_401
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1667941163
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1667941163
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1667941163
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_114
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1667941163
transform 1 0 14628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_174
timestamp 1667941163
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_182
timestamp 1667941163
transform 1 0 17848 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1667941163
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1667941163
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_243
timestamp 1667941163
transform 1 0 23460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1667941163
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_264
timestamp 1667941163
transform 1 0 25392 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_270
timestamp 1667941163
transform 1 0 25944 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_274
timestamp 1667941163
transform 1 0 26312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_281
timestamp 1667941163
transform 1 0 26956 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_288
timestamp 1667941163
transform 1 0 27600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_295
timestamp 1667941163
transform 1 0 28244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1667941163
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1667941163
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_328
timestamp 1667941163
transform 1 0 31280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1667941163
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_342
timestamp 1667941163
transform 1 0 32568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_349
timestamp 1667941163
transform 1 0 33212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1667941163
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1667941163
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1667941163
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_70
timestamp 1667941163
transform 1 0 7544 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_78
timestamp 1667941163
transform 1 0 8280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_102
timestamp 1667941163
transform 1 0 10488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_106
timestamp 1667941163
transform 1 0 10856 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1667941163
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1667941163
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_247
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_258
timestamp 1667941163
transform 1 0 24840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_265
timestamp 1667941163
transform 1 0 25484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_272
timestamp 1667941163
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_292
timestamp 1667941163
transform 1 0 27968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1667941163
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_319
timestamp 1667941163
transform 1 0 30452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_326
timestamp 1667941163
transform 1 0 31096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1667941163
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_342
timestamp 1667941163
transform 1 0 32568 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_354
timestamp 1667941163
transform 1 0 33672 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_366
timestamp 1667941163
transform 1 0 34776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_378
timestamp 1667941163
transform 1 0 35880 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1667941163
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1667941163
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1667941163
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1667941163
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1667941163
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_108
timestamp 1667941163
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1667941163
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1667941163
transform 1 0 14720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1667941163
transform 1 0 17020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_182
timestamp 1667941163
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1667941163
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1667941163
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_238
timestamp 1667941163
transform 1 0 23000 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 1667941163
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_264
timestamp 1667941163
transform 1 0 25392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1667941163
transform 1 0 26036 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_278
timestamp 1667941163
transform 1 0 26680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_285
timestamp 1667941163
transform 1 0 27324 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_292
timestamp 1667941163
transform 1 0 27968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_299
timestamp 1667941163
transform 1 0 28612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1667941163
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_314
timestamp 1667941163
transform 1 0 29992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_328
timestamp 1667941163
transform 1 0 31280 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_335
timestamp 1667941163
transform 1 0 31924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_347
timestamp 1667941163
transform 1 0 33028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1667941163
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_371
timestamp 1667941163
transform 1 0 35236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_375
timestamp 1667941163
transform 1 0 35604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_387
timestamp 1667941163
transform 1 0 36708 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_399
timestamp 1667941163
transform 1 0 37812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1667941163
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_21
timestamp 1667941163
transform 1 0 3036 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1667941163
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1667941163
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1667941163
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_82
timestamp 1667941163
transform 1 0 8648 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1667941163
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_144
timestamp 1667941163
transform 1 0 14352 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_156
timestamp 1667941163
transform 1 0 15456 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_162
timestamp 1667941163
transform 1 0 16008 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1667941163
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_192
timestamp 1667941163
transform 1 0 18768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_198
timestamp 1667941163
transform 1 0 19320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1667941163
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1667941163
transform 1 0 22540 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_250
timestamp 1667941163
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_257
timestamp 1667941163
transform 1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_264
timestamp 1667941163
transform 1 0 25392 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_271
timestamp 1667941163
transform 1 0 26036 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1667941163
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_300
timestamp 1667941163
transform 1 0 28704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_307
timestamp 1667941163
transform 1 0 29348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_314
timestamp 1667941163
transform 1 0 29992 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_321
timestamp 1667941163
transform 1 0 30636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_333
timestamp 1667941163
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1667941163
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1667941163
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1667941163
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1667941163
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_91
timestamp 1667941163
transform 1 0 9476 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_120
timestamp 1667941163
transform 1 0 12144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1667941163
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_149
timestamp 1667941163
transform 1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_173
timestamp 1667941163
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_181
timestamp 1667941163
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1667941163
transform 1 0 19596 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_222
timestamp 1667941163
transform 1 0 21528 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1667941163
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_272
timestamp 1667941163
transform 1 0 26128 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_279
timestamp 1667941163
transform 1 0 26772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1667941163
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_298
timestamp 1667941163
transform 1 0 28520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_302
timestamp 1667941163
transform 1 0 28888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1667941163
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_314
timestamp 1667941163
transform 1 0 29992 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_326
timestamp 1667941163
transform 1 0 31096 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_338
timestamp 1667941163
transform 1 0 32200 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_346
timestamp 1667941163
transform 1 0 32936 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_352
timestamp 1667941163
transform 1 0 33488 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_22
timestamp 1667941163
transform 1 0 3128 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp 1667941163
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1667941163
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1667941163
transform 1 0 6808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_70
timestamp 1667941163
transform 1 0 7544 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_95
timestamp 1667941163
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_152
timestamp 1667941163
transform 1 0 15088 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1667941163
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_191
timestamp 1667941163
transform 1 0 18676 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1667941163
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_247
timestamp 1667941163
transform 1 0 23828 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_254
timestamp 1667941163
transform 1 0 24472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_268
timestamp 1667941163
transform 1 0 25760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1667941163
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_286
timestamp 1667941163
transform 1 0 27416 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_298
timestamp 1667941163
transform 1 0 28520 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_310
timestamp 1667941163
transform 1 0 29624 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_322
timestamp 1667941163
transform 1 0 30728 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1667941163
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1667941163
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1667941163
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1667941163
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1667941163
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_58
timestamp 1667941163
transform 1 0 6440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_105
timestamp 1667941163
transform 1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1667941163
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1667941163
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_147
timestamp 1667941163
transform 1 0 14628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_159
timestamp 1667941163
transform 1 0 15732 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_163
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_185
timestamp 1667941163
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1667941163
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_223
timestamp 1667941163
transform 1 0 21620 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_235
timestamp 1667941163
transform 1 0 22724 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_241
timestamp 1667941163
transform 1 0 23276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_268
timestamp 1667941163
transform 1 0 25760 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_283
timestamp 1667941163
transform 1 0 27140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_290
timestamp 1667941163
transform 1 0 27784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_296
timestamp 1667941163
transform 1 0 28336 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1667941163
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1667941163
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1667941163
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_28
timestamp 1667941163
transform 1 0 3680 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_65
timestamp 1667941163
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1667941163
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_126
timestamp 1667941163
transform 1 0 12696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_130
timestamp 1667941163
transform 1 0 13064 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_152
timestamp 1667941163
transform 1 0 15088 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1667941163
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1667941163
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1667941163
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1667941163
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_291
timestamp 1667941163
transform 1 0 27876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_298
timestamp 1667941163
transform 1 0 28520 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_312
timestamp 1667941163
transform 1 0 29808 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_324
timestamp 1667941163
transform 1 0 30912 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_379
timestamp 1667941163
transform 1 0 35972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_383
timestamp 1667941163
transform 1 0 36340 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_13
timestamp 1667941163
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1667941163
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_34
timestamp 1667941163
transform 1 0 4232 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1667941163
transform 1 0 4784 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1667941163
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1667941163
transform 1 0 5796 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1667941163
transform 1 0 6532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1667941163
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_113
timestamp 1667941163
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1667941163
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1667941163
transform 1 0 14536 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_173
timestamp 1667941163
transform 1 0 17020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_185
timestamp 1667941163
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1667941163
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1667941163
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1667941163
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_284
timestamp 1667941163
transform 1 0 27232 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_296
timestamp 1667941163
transform 1 0 28336 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_370
timestamp 1667941163
transform 1 0 35144 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_382
timestamp 1667941163
transform 1 0 36248 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_394
timestamp 1667941163
transform 1 0 37352 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_400
timestamp 1667941163
transform 1 0 37904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1667941163
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1667941163
transform 1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_18
timestamp 1667941163
transform 1 0 2760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_25
timestamp 1667941163
transform 1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1667941163
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1667941163
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1667941163
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_118
timestamp 1667941163
transform 1 0 11960 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 1667941163
transform 1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_152
timestamp 1667941163
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1667941163
transform 1 0 15732 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_191
timestamp 1667941163
transform 1 0 18676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_199
timestamp 1667941163
transform 1 0 19412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1667941163
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_242
timestamp 1667941163
transform 1 0 23368 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_248
timestamp 1667941163
transform 1 0 23920 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_252
timestamp 1667941163
transform 1 0 24288 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_265
timestamp 1667941163
transform 1 0 25484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_272
timestamp 1667941163
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_298
timestamp 1667941163
transform 1 0 28520 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_311
timestamp 1667941163
transform 1 0 29716 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_315
timestamp 1667941163
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_327
timestamp 1667941163
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1667941163
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1667941163
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_18
timestamp 1667941163
transform 1 0 2760 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1667941163
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp 1667941163
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1667941163
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1667941163
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_154
timestamp 1667941163
transform 1 0 15272 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_160
timestamp 1667941163
transform 1 0 15824 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1667941163
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1667941163
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1667941163
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_285
timestamp 1667941163
transform 1 0 27324 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_320
timestamp 1667941163
transform 1 0 30544 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_332
timestamp 1667941163
transform 1 0 31648 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_344
timestamp 1667941163
transform 1 0 32752 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_356
timestamp 1667941163
transform 1 0 33856 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_397
timestamp 1667941163
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_402
timestamp 1667941163
transform 1 0 38088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1667941163
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1667941163
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_25
timestamp 1667941163
transform 1 0 3404 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_36
timestamp 1667941163
transform 1 0 4416 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1667941163
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1667941163
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_94
timestamp 1667941163
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1667941163
transform 1 0 10396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1667941163
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_119
timestamp 1667941163
transform 1 0 12052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_128
timestamp 1667941163
transform 1 0 12880 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_153
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1667941163
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1667941163
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_247
timestamp 1667941163
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_259
timestamp 1667941163
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_271
timestamp 1667941163
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_299
timestamp 1667941163
transform 1 0 28612 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_311
timestamp 1667941163
transform 1 0 29716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_323
timestamp 1667941163
transform 1 0 30820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1667941163
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_36
timestamp 1667941163
transform 1 0 4416 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_43
timestamp 1667941163
transform 1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_58
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_92
timestamp 1667941163
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1667941163
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_126
timestamp 1667941163
transform 1 0 12696 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 1667941163
transform 1 0 13248 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1667941163
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1667941163
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1667941163
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_282
timestamp 1667941163
transform 1 0 27048 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_294
timestamp 1667941163
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1667941163
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_351
timestamp 1667941163
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1667941163
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_20
timestamp 1667941163
transform 1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1667941163
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_33
timestamp 1667941163
transform 1 0 4140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1667941163
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_47
timestamp 1667941163
transform 1 0 5428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1667941163
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_89
timestamp 1667941163
transform 1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1667941163
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_177
timestamp 1667941163
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1667941163
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1667941163
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1667941163
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_232
timestamp 1667941163
transform 1 0 22448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_256
timestamp 1667941163
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1667941163
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_270
timestamp 1667941163
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_296
timestamp 1667941163
transform 1 0 28336 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_308
timestamp 1667941163
transform 1 0 29440 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_320
timestamp 1667941163
transform 1 0 30544 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1667941163
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_379
timestamp 1667941163
transform 1 0 35972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1667941163
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_16
timestamp 1667941163
transform 1 0 2576 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_50
timestamp 1667941163
transform 1 0 5704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1667941163
transform 1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1667941163
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_111
timestamp 1667941163
transform 1 0 11316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1667941163
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_147
timestamp 1667941163
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1667941163
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_178
timestamp 1667941163
transform 1 0 17480 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1667941163
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_220
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_228
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_238
timestamp 1667941163
transform 1 0 23000 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_258
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_270
timestamp 1667941163
transform 1 0 25944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_275
timestamp 1667941163
transform 1 0 26404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_284
timestamp 1667941163
transform 1 0 27232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1667941163
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1667941163
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1667941163
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_324
timestamp 1667941163
transform 1 0 30912 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_336
timestamp 1667941163
transform 1 0 32016 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_348
timestamp 1667941163
transform 1 0 33120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1667941163
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_17
timestamp 1667941163
transform 1 0 2668 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1667941163
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_35
timestamp 1667941163
transform 1 0 4324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_42
timestamp 1667941163
transform 1 0 4968 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1667941163
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_86
timestamp 1667941163
transform 1 0 9016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1667941163
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1667941163
transform 1 0 17388 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_204
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_213
timestamp 1667941163
transform 1 0 20700 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1667941163
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1667941163
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1667941163
transform 1 0 23092 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1667941163
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 1667941163
transform 1 0 24380 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_260
timestamp 1667941163
transform 1 0 25024 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1667941163
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_309
timestamp 1667941163
transform 1 0 29532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_321
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1667941163
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_40
timestamp 1667941163
transform 1 0 4784 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_49
timestamp 1667941163
transform 1 0 5612 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_56
timestamp 1667941163
transform 1 0 6256 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_73
timestamp 1667941163
transform 1 0 7820 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1667941163
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1667941163
transform 1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_134
timestamp 1667941163
transform 1 0 13432 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1667941163
transform 1 0 16008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_176
timestamp 1667941163
transform 1 0 17296 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1667941163
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_214
timestamp 1667941163
transform 1 0 20792 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1667941163
transform 1 0 22080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1667941163
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1667941163
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1667941163
transform 1 0 25760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_285
timestamp 1667941163
transform 1 0 27324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_291
timestamp 1667941163
transform 1 0 27876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1667941163
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1667941163
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_31
timestamp 1667941163
transform 1 0 3956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_40
timestamp 1667941163
transform 1 0 4784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_47
timestamp 1667941163
transform 1 0 5428 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1667941163
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_76
timestamp 1667941163
transform 1 0 8096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1667941163
transform 1 0 8740 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1667941163
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_119
timestamp 1667941163
transform 1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1667941163
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1667941163
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1667941163
transform 1 0 18032 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_230
timestamp 1667941163
transform 1 0 22264 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_238
timestamp 1667941163
transform 1 0 23000 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_253
timestamp 1667941163
transform 1 0 24380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_260
timestamp 1667941163
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_267
timestamp 1667941163
transform 1 0 25668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1667941163
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_292
timestamp 1667941163
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_304
timestamp 1667941163
transform 1 0 29072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_315
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_327
timestamp 1667941163
transform 1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_9
timestamp 1667941163
transform 1 0 1932 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_48
timestamp 1667941163
transform 1 0 5520 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1667941163
transform 1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_61
timestamp 1667941163
transform 1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_68
timestamp 1667941163
transform 1 0 7360 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_75
timestamp 1667941163
transform 1 0 8004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1667941163
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1667941163
transform 1 0 9660 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_100
timestamp 1667941163
transform 1 0 10304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_117
timestamp 1667941163
transform 1 0 11868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1667941163
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1667941163
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_169
timestamp 1667941163
transform 1 0 16652 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_184
timestamp 1667941163
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_212
timestamp 1667941163
transform 1 0 20608 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_220
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_225
timestamp 1667941163
transform 1 0 21804 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_233
timestamp 1667941163
transform 1 0 22540 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1667941163
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_265
timestamp 1667941163
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_271
timestamp 1667941163
transform 1 0 26036 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_275
timestamp 1667941163
transform 1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_281
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_285
timestamp 1667941163
transform 1 0 27324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_292
timestamp 1667941163
transform 1 0 27968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1667941163
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1667941163
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_313
timestamp 1667941163
transform 1 0 29900 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_322
timestamp 1667941163
transform 1 0 30728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_334
timestamp 1667941163
transform 1 0 31832 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_346
timestamp 1667941163
transform 1 0 32936 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1667941163
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1667941163
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_19
timestamp 1667941163
transform 1 0 2852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1667941163
transform 1 0 3496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp 1667941163
transform 1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_40
timestamp 1667941163
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1667941163
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1667941163
transform 1 0 7176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_73
timestamp 1667941163
transform 1 0 7820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_80
timestamp 1667941163
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_87
timestamp 1667941163
transform 1 0 9108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1667941163
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1667941163
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1667941163
transform 1 0 12788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1667941163
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_148
timestamp 1667941163
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1667941163
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_204
timestamp 1667941163
transform 1 0 19872 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_211
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1667941163
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_253
timestamp 1667941163
transform 1 0 24380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_265
timestamp 1667941163
transform 1 0 25484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1667941163
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_285
timestamp 1667941163
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1667941163
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1667941163
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_303
timestamp 1667941163
transform 1 0 28980 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_318
timestamp 1667941163
transform 1 0 30360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_330
timestamp 1667941163
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_402
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1667941163
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1667941163
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_19
timestamp 1667941163
transform 1 0 2852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1667941163
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_37
timestamp 1667941163
transform 1 0 4508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_50
timestamp 1667941163
transform 1 0 5704 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_64
timestamp 1667941163
transform 1 0 6992 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_75
timestamp 1667941163
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_102
timestamp 1667941163
transform 1 0 10488 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1667941163
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1667941163
transform 1 0 13156 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_174
timestamp 1667941163
transform 1 0 17112 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_216
timestamp 1667941163
transform 1 0 20976 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_225
timestamp 1667941163
transform 1 0 21804 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_233
timestamp 1667941163
transform 1 0 22540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_243
timestamp 1667941163
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1667941163
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1667941163
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_301
timestamp 1667941163
transform 1 0 28796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1667941163
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_324
timestamp 1667941163
transform 1 0 30912 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_336
timestamp 1667941163
transform 1 0 32016 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_348
timestamp 1667941163
transform 1 0 33120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1667941163
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1667941163
transform 1 0 2944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1667941163
transform 1 0 4232 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1667941163
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1667941163
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_73
timestamp 1667941163
transform 1 0 7820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1667941163
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1667941163
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1667941163
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1667941163
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 1667941163
transform 1 0 12696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1667941163
transform 1 0 14260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_159
timestamp 1667941163
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 1667941163
transform 1 0 17388 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_186
timestamp 1667941163
transform 1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_194
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_198
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_206
timestamp 1667941163
transform 1 0 20056 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1667941163
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1667941163
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_234
timestamp 1667941163
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_248
timestamp 1667941163
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_265
timestamp 1667941163
transform 1 0 25484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1667941163
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1667941163
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1667941163
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_401
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1667941163
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_17
timestamp 1667941163
transform 1 0 2668 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1667941163
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_40
timestamp 1667941163
transform 1 0 4784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1667941163
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_54
timestamp 1667941163
transform 1 0 6072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1667941163
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1667941163
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1667941163
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1667941163
transform 1 0 9476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1667941163
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_108
timestamp 1667941163
transform 1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1667941163
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_147
timestamp 1667941163
transform 1 0 14628 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_164
timestamp 1667941163
transform 1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_173
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1667941163
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1667941163
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1667941163
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1667941163
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1667941163
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1667941163
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_258
timestamp 1667941163
transform 1 0 24840 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_270
timestamp 1667941163
transform 1 0 25944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_274
timestamp 1667941163
transform 1 0 26312 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_282
timestamp 1667941163
transform 1 0 27048 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_286
timestamp 1667941163
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_298
timestamp 1667941163
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_314
timestamp 1667941163
transform 1 0 29992 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_326
timestamp 1667941163
transform 1 0 31096 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_338
timestamp 1667941163
transform 1 0 32200 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_350
timestamp 1667941163
transform 1 0 33304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_23
timestamp 1667941163
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_29
timestamp 1667941163
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1667941163
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_43
timestamp 1667941163
transform 1 0 5060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_63
timestamp 1667941163
transform 1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_76
timestamp 1667941163
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_92
timestamp 1667941163
transform 1 0 9568 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_100
timestamp 1667941163
transform 1 0 10304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1667941163
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_121
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_128
timestamp 1667941163
transform 1 0 12880 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_138
timestamp 1667941163
transform 1 0 13800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_151
timestamp 1667941163
transform 1 0 14996 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1667941163
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_191
timestamp 1667941163
transform 1 0 18676 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_204
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1667941163
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1667941163
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_257
timestamp 1667941163
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_264
timestamp 1667941163
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_268
timestamp 1667941163
transform 1 0 25760 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_312
timestamp 1667941163
transform 1 0 29808 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_324
timestamp 1667941163
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_401
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_38
timestamp 1667941163
transform 1 0 4600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_50
timestamp 1667941163
transform 1 0 5704 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_55
timestamp 1667941163
transform 1 0 6164 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1667941163
transform 1 0 6808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_74
timestamp 1667941163
transform 1 0 7912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_78
timestamp 1667941163
transform 1 0 8280 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1667941163
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1667941163
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_101
timestamp 1667941163
transform 1 0 10396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_111
timestamp 1667941163
transform 1 0 11316 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_118
timestamp 1667941163
transform 1 0 11960 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_125
timestamp 1667941163
transform 1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1667941163
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_160
timestamp 1667941163
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_167
timestamp 1667941163
transform 1 0 16468 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_175
timestamp 1667941163
transform 1 0 17204 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_185
timestamp 1667941163
transform 1 0 18124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1667941163
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1667941163
transform 1 0 19780 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_214
timestamp 1667941163
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_226
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_234
timestamp 1667941163
transform 1 0 22632 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_238
timestamp 1667941163
transform 1 0 23000 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1667941163
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_261
timestamp 1667941163
transform 1 0 25116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_268
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_281
timestamp 1667941163
transform 1 0 26956 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_290
timestamp 1667941163
transform 1 0 27784 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1667941163
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_314
timestamp 1667941163
transform 1 0 29992 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_326
timestamp 1667941163
transform 1 0 31096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_334
timestamp 1667941163
transform 1 0 31832 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_340
timestamp 1667941163
transform 1 0 32384 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_352
timestamp 1667941163
transform 1 0 33488 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1667941163
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1667941163
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1667941163
transform 1 0 4048 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_42
timestamp 1667941163
transform 1 0 4968 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_50
timestamp 1667941163
transform 1 0 5704 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_68
timestamp 1667941163
transform 1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1667941163
transform 1 0 8004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1667941163
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_103
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1667941163
transform 1 0 11960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_147
timestamp 1667941163
transform 1 0 14628 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_155
timestamp 1667941163
transform 1 0 15364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1667941163
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_191
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1667941163
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_204
timestamp 1667941163
transform 1 0 19872 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1667941163
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_240
timestamp 1667941163
transform 1 0 23184 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1667941163
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1667941163
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_304
timestamp 1667941163
transform 1 0 29072 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_316
timestamp 1667941163
transform 1 0 30176 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1667941163
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_40
timestamp 1667941163
transform 1 0 4784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_48
timestamp 1667941163
transform 1 0 5520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1667941163
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1667941163
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_68
timestamp 1667941163
transform 1 0 7360 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1667941163
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_96
timestamp 1667941163
transform 1 0 9936 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_102
timestamp 1667941163
transform 1 0 10488 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_112
timestamp 1667941163
transform 1 0 11408 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1667941163
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_161
timestamp 1667941163
transform 1 0 15916 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_172
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_181
timestamp 1667941163
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_212
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_221
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_229
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_240
timestamp 1667941163
transform 1 0 23184 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_260
timestamp 1667941163
transform 1 0 25024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_267
timestamp 1667941163
transform 1 0 25668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_271
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_275
timestamp 1667941163
transform 1 0 26404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_281
timestamp 1667941163
transform 1 0 26956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_285
timestamp 1667941163
transform 1 0 27324 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_296
timestamp 1667941163
transform 1 0 28336 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_8
timestamp 1667941163
transform 1 0 1840 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_20
timestamp 1667941163
transform 1 0 2944 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_32
timestamp 1667941163
transform 1 0 4048 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1667941163
transform 1 0 4876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1667941163
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1667941163
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1667941163
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_89
timestamp 1667941163
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_100
timestamp 1667941163
transform 1 0 10304 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1667941163
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_117
timestamp 1667941163
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_131
timestamp 1667941163
transform 1 0 13156 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_148
timestamp 1667941163
transform 1 0 14720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1667941163
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_175
timestamp 1667941163
transform 1 0 17204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_190
timestamp 1667941163
transform 1 0 18584 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_198
timestamp 1667941163
transform 1 0 19320 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_202
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_242
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_266
timestamp 1667941163
transform 1 0 25576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_297
timestamp 1667941163
transform 1 0 28428 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_301
timestamp 1667941163
transform 1 0 28796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_313
timestamp 1667941163
transform 1 0 29900 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_318
timestamp 1667941163
transform 1 0 30360 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_330
timestamp 1667941163
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_70
timestamp 1667941163
transform 1 0 7544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_101
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_108
timestamp 1667941163
transform 1 0 11040 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1667941163
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_171
timestamp 1667941163
transform 1 0 16836 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_179
timestamp 1667941163
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_202
timestamp 1667941163
transform 1 0 19688 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_206
timestamp 1667941163
transform 1 0 20056 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1667941163
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_222
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_230
timestamp 1667941163
transform 1 0 22264 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_235
timestamp 1667941163
transform 1 0 22724 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1667941163
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1667941163
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_293
timestamp 1667941163
transform 1 0 28060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1667941163
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_326
timestamp 1667941163
transform 1 0 31096 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_338
timestamp 1667941163
transform 1 0 32200 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_350
timestamp 1667941163
transform 1 0 33304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1667941163
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_76
timestamp 1667941163
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_97
timestamp 1667941163
transform 1 0 10028 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 1667941163
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_129
timestamp 1667941163
transform 1 0 12972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_133
timestamp 1667941163
transform 1 0 13340 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_145
timestamp 1667941163
transform 1 0 14444 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1667941163
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1667941163
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_175
timestamp 1667941163
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_182
timestamp 1667941163
transform 1 0 17848 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1667941163
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1667941163
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_203
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1667941163
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1667941163
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_245
timestamp 1667941163
transform 1 0 23644 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_252
timestamp 1667941163
transform 1 0 24288 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_264
timestamp 1667941163
transform 1 0 25392 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1667941163
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_301
timestamp 1667941163
transform 1 0 28796 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_306
timestamp 1667941163
transform 1 0 29256 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_318
timestamp 1667941163
transform 1 0 30360 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_330
timestamp 1667941163
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_358
timestamp 1667941163
transform 1 0 34040 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_370
timestamp 1667941163
transform 1 0 35144 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_382
timestamp 1667941163
transform 1 0 36248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1667941163
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_62
timestamp 1667941163
transform 1 0 6808 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_69
timestamp 1667941163
transform 1 0 7452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1667941163
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_113
timestamp 1667941163
transform 1 0 11500 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_125
timestamp 1667941163
transform 1 0 12604 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_129
timestamp 1667941163
transform 1 0 12972 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1667941163
transform 1 0 15272 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_158
timestamp 1667941163
transform 1 0 15640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1667941163
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_212
timestamp 1667941163
transform 1 0 20608 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_233
timestamp 1667941163
transform 1 0 22540 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1667941163
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1667941163
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_258
timestamp 1667941163
transform 1 0 24840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_270
timestamp 1667941163
transform 1 0 25944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_278
timestamp 1667941163
transform 1 0 26680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_282
timestamp 1667941163
transform 1 0 27048 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_290
timestamp 1667941163
transform 1 0 27784 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1667941163
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_353
timestamp 1667941163
transform 1 0 33580 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1667941163
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1667941163
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1667941163
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1667941163
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_65
timestamp 1667941163
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_77
timestamp 1667941163
transform 1 0 8188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1667941163
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_90
timestamp 1667941163
transform 1 0 9384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_129
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_135
timestamp 1667941163
transform 1 0 13524 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_145
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_151
timestamp 1667941163
transform 1 0 14996 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1667941163
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_174
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1667941163
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1667941163
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_200
timestamp 1667941163
transform 1 0 19504 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_213
timestamp 1667941163
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1667941163
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_241
timestamp 1667941163
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_250
timestamp 1667941163
transform 1 0 24104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_258
timestamp 1667941163
transform 1 0 24840 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_264
timestamp 1667941163
transform 1 0 25392 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_268
timestamp 1667941163
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1667941163
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_299
timestamp 1667941163
transform 1 0 28612 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_311
timestamp 1667941163
transform 1 0 29716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_323
timestamp 1667941163
transform 1 0 30820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_330
timestamp 1667941163
transform 1 0 31464 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_10
timestamp 1667941163
transform 1 0 2024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_22
timestamp 1667941163
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_68
timestamp 1667941163
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1667941163
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1667941163
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1667941163
transform 1 0 12420 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1667941163
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_173
timestamp 1667941163
transform 1 0 17020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1667941163
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1667941163
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1667941163
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_329
timestamp 1667941163
transform 1 0 31372 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_9
timestamp 1667941163
transform 1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_16
timestamp 1667941163
transform 1 0 2576 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_28
timestamp 1667941163
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_40
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1667941163
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_63
timestamp 1667941163
transform 1 0 6900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_67
timestamp 1667941163
transform 1 0 7268 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_75
timestamp 1667941163
transform 1 0 8004 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1667941163
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_97
timestamp 1667941163
transform 1 0 10028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_127
timestamp 1667941163
transform 1 0 12788 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_135
timestamp 1667941163
transform 1 0 13524 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_139
timestamp 1667941163
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1667941163
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_153
timestamp 1667941163
transform 1 0 15180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1667941163
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_193
timestamp 1667941163
transform 1 0 18860 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_209
timestamp 1667941163
transform 1 0 20332 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_230
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_238
timestamp 1667941163
transform 1 0 23000 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_254
timestamp 1667941163
transform 1 0 24472 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1667941163
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1667941163
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_301
timestamp 1667941163
transform 1 0 28796 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_307
timestamp 1667941163
transform 1 0 29348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_319
timestamp 1667941163
transform 1 0 30452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1667941163
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_71
timestamp 1667941163
transform 1 0 7636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1667941163
transform 1 0 8004 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_90
timestamp 1667941163
transform 1 0 9384 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_102
timestamp 1667941163
transform 1 0 10488 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_107
timestamp 1667941163
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_127
timestamp 1667941163
transform 1 0 12788 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1667941163
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_147
timestamp 1667941163
transform 1 0 14628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_151
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_163
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_175
timestamp 1667941163
transform 1 0 17204 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_183
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_205
timestamp 1667941163
transform 1 0 19964 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1667941163
transform 1 0 20424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_214
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_218
timestamp 1667941163
transform 1 0 21160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_226
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1667941163
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1667941163
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1667941163
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_73
timestamp 1667941163
transform 1 0 7820 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_80
timestamp 1667941163
transform 1 0 8464 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_92
timestamp 1667941163
transform 1 0 9568 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_98
timestamp 1667941163
transform 1 0 10120 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1667941163
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_134
timestamp 1667941163
transform 1 0 13432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_159
timestamp 1667941163
transform 1 0 15732 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_176
timestamp 1667941163
transform 1 0 17296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_189
timestamp 1667941163
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_196
timestamp 1667941163
transform 1 0 19136 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_208
timestamp 1667941163
transform 1 0 20240 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1667941163
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_242
timestamp 1667941163
transform 1 0 23368 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_254
timestamp 1667941163
transform 1 0 24472 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1667941163
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1667941163
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_324
timestamp 1667941163
transform 1 0 30912 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_21
timestamp 1667941163
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_92
timestamp 1667941163
transform 1 0 9568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1667941163
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1667941163
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_113
timestamp 1667941163
transform 1 0 11500 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_119
timestamp 1667941163
transform 1 0 12052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1667941163
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_164
timestamp 1667941163
transform 1 0 16192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_178
timestamp 1667941163
transform 1 0 17480 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1667941163
transform 1 0 18216 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1667941163
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_212
timestamp 1667941163
transform 1 0 20608 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_224
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_232
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_237
timestamp 1667941163
transform 1 0 22908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1667941163
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1667941163
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_65
timestamp 1667941163
transform 1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_71
timestamp 1667941163
transform 1 0 7636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_83
timestamp 1667941163
transform 1 0 8740 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_89
timestamp 1667941163
transform 1 0 9292 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_101
timestamp 1667941163
transform 1 0 10396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 1667941163
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_133
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_138
timestamp 1667941163
transform 1 0 13800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1667941163
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_155
timestamp 1667941163
transform 1 0 15364 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_159
timestamp 1667941163
transform 1 0 15732 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_180
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_192
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_204
timestamp 1667941163
transform 1 0 19872 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1667941163
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_243
timestamp 1667941163
transform 1 0 23460 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_255
timestamp 1667941163
transform 1 0 24564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_267
timestamp 1667941163
transform 1 0 25668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1667941163
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_146
timestamp 1667941163
transform 1 0 14536 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_154
timestamp 1667941163
transform 1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_166
timestamp 1667941163
transform 1 0 16376 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_172
timestamp 1667941163
transform 1 0 16928 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_176
timestamp 1667941163
transform 1 0 17296 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_184
timestamp 1667941163
transform 1 0 18032 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1667941163
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_295
timestamp 1667941163
transform 1 0 28244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_133
timestamp 1667941163
transform 1 0 13340 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_150
timestamp 1667941163
transform 1 0 14904 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_162
timestamp 1667941163
transform 1 0 16008 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_185
timestamp 1667941163
transform 1 0 18124 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_196
timestamp 1667941163
transform 1 0 19136 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_208
timestamp 1667941163
transform 1 0 20240 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1667941163
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1667941163
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1667941163
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1667941163
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1667941163
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_289
timestamp 1667941163
transform 1 0 27692 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_295
timestamp 1667941163
transform 1 0 28244 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_307
timestamp 1667941163
transform 1 0 29348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_319
timestamp 1667941163
transform 1 0 30452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1667941163
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_123
timestamp 1667941163
transform 1 0 12420 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_146
timestamp 1667941163
transform 1 0 14536 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_150
timestamp 1667941163
transform 1 0 14904 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_154
timestamp 1667941163
transform 1 0 15272 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_161
timestamp 1667941163
transform 1 0 15916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_173
timestamp 1667941163
transform 1 0 17020 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1667941163
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1667941163
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1667941163
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1667941163
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_370
timestamp 1667941163
transform 1 0 35144 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_382
timestamp 1667941163
transform 1 0 36248 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_394
timestamp 1667941163
transform 1 0 37352 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_64
timestamp 1667941163
transform 1 0 6992 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_76
timestamp 1667941163
transform 1 0 8096 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_88
timestamp 1667941163
transform 1 0 9200 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_100
timestamp 1667941163
transform 1 0 10304 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_130
timestamp 1667941163
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1667941163
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1667941163
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_231
timestamp 1667941163
transform 1 0 22356 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_243
timestamp 1667941163
transform 1 0 23460 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_255
timestamp 1667941163
transform 1 0 24564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_267
timestamp 1667941163
transform 1 0 25668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1667941163
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_369
timestamp 1667941163
transform 1 0 35052 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_374
timestamp 1667941163
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_386
timestamp 1667941163
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_8
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1667941163
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1667941163
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_401
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_156
timestamp 1667941163
transform 1 0 15456 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_248
timestamp 1667941163
transform 1 0 23920 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_260
timestamp 1667941163
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1667941163
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1667941163
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_372
timestamp 1667941163
transform 1 0 35328 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1667941163
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_120
timestamp 1667941163
transform 1 0 12144 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1667941163
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_183
timestamp 1667941163
transform 1 0 17940 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 1667941163
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1667941163
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_9
timestamp 1667941163
transform 1 0 1932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_21
timestamp 1667941163
transform 1 0 3036 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_33
timestamp 1667941163
transform 1 0 4140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_45
timestamp 1667941163
transform 1 0 5244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_145
timestamp 1667941163
transform 1 0 14444 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_155
timestamp 1667941163
transform 1 0 15364 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1667941163
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1667941163
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1667941163
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1667941163
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1667941163
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_8
timestamp 1667941163
transform 1 0 1840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1667941163
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_76
timestamp 1667941163
transform 1 0 8096 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_106
timestamp 1667941163
transform 1 0 10856 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_118
timestamp 1667941163
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_130
timestamp 1667941163
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1667941163
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1667941163
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1667941163
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1667941163
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_353
timestamp 1667941163
transform 1 0 33580 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_358
timestamp 1667941163
transform 1 0 34040 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_31
timestamp 1667941163
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_43
timestamp 1667941163
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_62
timestamp 1667941163
transform 1 0 6808 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_74
timestamp 1667941163
transform 1 0 7912 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_86
timestamp 1667941163
transform 1 0 9016 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_98
timestamp 1667941163
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_129
timestamp 1667941163
transform 1 0 12972 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_133
timestamp 1667941163
transform 1 0 13340 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_145
timestamp 1667941163
transform 1 0 14444 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_157
timestamp 1667941163
transform 1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1667941163
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_265
timestamp 1667941163
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1667941163
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_286
timestamp 1667941163
transform 1 0 27416 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_298
timestamp 1667941163
transform 1 0 28520 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_310
timestamp 1667941163
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_322
timestamp 1667941163
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1667941163
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_61
timestamp 1667941163
transform 1 0 6716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_73
timestamp 1667941163
transform 1 0 7820 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1667941163
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_105
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_111
timestamp 1667941163
transform 1 0 11316 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_123
timestamp 1667941163
transform 1 0 12420 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1667941163
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_314
timestamp 1667941163
transform 1 0 29992 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_318
timestamp 1667941163
transform 1 0 30360 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_322
timestamp 1667941163
transform 1 0 30728 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_334
timestamp 1667941163
transform 1 0 31832 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_346
timestamp 1667941163
transform 1 0 32936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1667941163
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_47
timestamp 1667941163
transform 1 0 5428 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1667941163
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1667941163
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1667941163
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_353
timestamp 1667941163
transform 1 0 33580 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_365
timestamp 1667941163
transform 1 0 34684 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_377
timestamp 1667941163
transform 1 0 35788 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1667941163
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_49
timestamp 1667941163
transform 1 0 5612 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_54
timestamp 1667941163
transform 1 0 6072 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_66
timestamp 1667941163
transform 1 0 7176 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_78
timestamp 1667941163
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_203
timestamp 1667941163
transform 1 0 19780 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_215
timestamp 1667941163
transform 1 0 20884 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_226
timestamp 1667941163
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_234
timestamp 1667941163
transform 1 0 22632 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_240
timestamp 1667941163
transform 1 0 23184 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_273
timestamp 1667941163
transform 1 0 26220 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_279
timestamp 1667941163
transform 1 0 26772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_291
timestamp 1667941163
transform 1 0 27876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1667941163
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_141
timestamp 1667941163
transform 1 0 14076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_153
timestamp 1667941163
transform 1 0 15180 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_157
timestamp 1667941163
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_165
timestamp 1667941163
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1667941163
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1667941163
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_34
timestamp 1667941163
transform 1 0 4232 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_46
timestamp 1667941163
transform 1 0 5336 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_58
timestamp 1667941163
transform 1 0 6440 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_70
timestamp 1667941163
transform 1 0 7544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1667941163
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_293
timestamp 1667941163
transform 1 0 28060 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_297
timestamp 1667941163
transform 1 0 28428 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_305
timestamp 1667941163
transform 1 0 29164 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_393
timestamp 1667941163
transform 1 0 37260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_397
timestamp 1667941163
transform 1 0 37628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_35
timestamp 1667941163
transform 1 0 4324 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_40
timestamp 1667941163
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1667941163
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1667941163
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1667941163
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1667941163
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1667941163
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1667941163
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1667941163
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1667941163
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_8
timestamp 1667941163
transform 1 0 1840 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_20
timestamp 1667941163
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_32
timestamp 1667941163
transform 1 0 4048 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_44
timestamp 1667941163
transform 1 0 5152 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_121
timestamp 1667941163
transform 1 0 12236 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_127
timestamp 1667941163
transform 1 0 12788 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_139
timestamp 1667941163
transform 1 0 13892 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_151
timestamp 1667941163
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1667941163
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_8
timestamp 1667941163
transform 1 0 1840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_20
timestamp 1667941163
transform 1 0 2944 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1667941163
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_16
timestamp 1667941163
transform 1 0 2576 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_23
timestamp 1667941163
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1667941163
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_90
timestamp 1667941163
transform 1 0 9384 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_102
timestamp 1667941163
transform 1 0 10488 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1667941163
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_132
timestamp 1667941163
transform 1 0 13248 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_144
timestamp 1667941163
transform 1 0 14352 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_156
timestamp 1667941163
transform 1 0 15456 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_174
timestamp 1667941163
transform 1 0 17112 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_183
timestamp 1667941163
transform 1 0 17940 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_195
timestamp 1667941163
transform 1 0 19044 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_203
timestamp 1667941163
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1667941163
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_244
timestamp 1667941163
transform 1 0 23552 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_256
timestamp 1667941163
transform 1 0 24656 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_268
timestamp 1667941163
transform 1 0 25760 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_301
timestamp 1667941163
transform 1 0 28796 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_308
timestamp 1667941163
transform 1 0 29440 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_320
timestamp 1667941163
transform 1 0 30544 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_328
timestamp 1667941163
transform 1 0 31280 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1667941163
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_377
timestamp 1667941163
transform 1 0 35788 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_386
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1667941163
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1667941163
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1667941163
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_144
timestamp 1667941163
transform 1 0 14352 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_148
timestamp 1667941163
transform 1 0 14720 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1667941163
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1667941163
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_270
timestamp 1667941163
transform 1 0 25944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_289
timestamp 1667941163
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1667941163
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1667941163
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_329
timestamp 1667941163
transform 1 0 31372 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1667941163
transform 1 0 31924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0384_
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0385_
timestamp 1667941163
transform 1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0386_
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0387_
timestamp 1667941163
transform 1 0 25392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0388_
timestamp 1667941163
transform 1 0 29532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0389_
timestamp 1667941163
transform 1 0 32292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0390_
timestamp 1667941163
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0392_
timestamp 1667941163
transform 1 0 31464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0393_
timestamp 1667941163
transform 1 0 29808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0394_
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0395_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 24748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0397_
timestamp 1667941163
transform 1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0398_
timestamp 1667941163
transform 1 0 25208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0399_
timestamp 1667941163
transform 1 0 21160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0400_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0401_
timestamp 1667941163
transform 1 0 16652 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1667941163
transform 1 0 24748 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0403_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0406_
timestamp 1667941163
transform 1 0 24472 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0407_
timestamp 1667941163
transform 1 0 11960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0408_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0409_
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0410_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 17848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0413_
timestamp 1667941163
transform 1 0 27048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0414_
timestamp 1667941163
transform 1 0 28244 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0416_
timestamp 1667941163
transform 1 0 28704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0418_
timestamp 1667941163
transform 1 0 20884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 21068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 21252 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0422_
timestamp 1667941163
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 20148 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 22540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 23184 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0426_
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0427_
timestamp 1667941163
transform 1 0 28428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0428_
timestamp 1667941163
transform 1 0 22448 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1667941163
transform 1 0 23552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 27048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 27508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 28980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0436_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 15640 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 14996 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0440_
timestamp 1667941163
transform 1 0 13524 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 13432 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 13524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0444_
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1667941163
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0446_
timestamp 1667941163
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1667941163
transform 1 0 7176 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 20884 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1667941163
transform 1 0 30360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1667941163
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 28980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 30360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 32292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1667941163
transform 1 0 9292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1667941163
transform 1 0 10580 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 8188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1667941163
transform 1 0 9016 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1667941163
transform 1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0462_
timestamp 1667941163
transform 1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0463_
timestamp 1667941163
transform 1 0 22172 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 4784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0466_
timestamp 1667941163
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0467_
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1667941163
transform 1 0 3496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0469_
timestamp 1667941163
transform 1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0472_
timestamp 1667941163
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0473_
timestamp 1667941163
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0474_
timestamp 1667941163
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0475_
timestamp 1667941163
transform 1 0 11960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 11684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0478_
timestamp 1667941163
transform 1 0 4600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0479_
timestamp 1667941163
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 7176 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0484_
timestamp 1667941163
transform 1 0 6992 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0485_
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 8832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 14904 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 10120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 13616 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 27784 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 26772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 6900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 4140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 32936 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 26680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 17940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 16744 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 16100 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 18400 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 25024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 9752 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 20516 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 12052 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 10672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 14352 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 19596 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 12696 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 18400 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 14260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 15456 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 11224 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 17572 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 26956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 21528 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 21160 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 25668 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 27784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 28428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 2300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 27140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 26036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 23368 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 10764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 18400 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 9108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 5888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 28244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 10764 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 9108 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 27140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 16928 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 29072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 21528 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 25392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 21160 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 7728 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 28336 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 26128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 17204 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 17480 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 4140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 11040 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 31464 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 36340 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 29624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 34224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 2760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 25668 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 35512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 27140 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 36708 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 8280 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 28980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 25024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 33212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0627_
timestamp 1667941163
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 7820 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 15456 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 5796 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 6808 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 35236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 19504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 7544 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 14536 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 30452 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 21620 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 5704 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 32292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 10580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 19688 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 31188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 4600 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 23644 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 21068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 8004 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 31648 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 25208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 4140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 27692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 18032 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 27968 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 22908 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 6716 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 12328 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 19136 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 16192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 11868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 23092 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 4416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 6532 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 16100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 9108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 31004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 26128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 34224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 27968 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 13800 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 29072 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 27784 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 30084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 26772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 25484 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 12144 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 15272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 17848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 3772 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 6532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 29716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 33120 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 32936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 29072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 7360 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0710_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _0711_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 28612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 24104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 30360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 33580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0722_
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 27048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 25760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 26036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 27968 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 23736 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 28336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0733_
timestamp 1667941163
transform 1 0 12236 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 22448 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 32292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0744_
timestamp 1667941163
transform 1 0 18400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 30176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 34868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 27140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 31004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0755_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 3864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 9936 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 19596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 8464 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0766_
timestamp 1667941163
transform 1 0 12144 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 7820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 6532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 7544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 6900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0777_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 4508 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 4508 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 6440 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 3404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0788_
timestamp 1667941163
transform 1 0 14720 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 7728 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 24380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 30360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 12512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 27324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 28428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0799_
timestamp 1667941163
transform 1 0 13248 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 15456 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 3956 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 3220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0810_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 4784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 4232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 16100 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0821_
timestamp 1667941163
transform 1 0 10764 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 6164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 20424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 20240 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 25208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 24748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0832_
timestamp 1667941163
transform 1 0 11040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 26128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 26772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 29716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 25760 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 26496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0843_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1656 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0844_
timestamp 1667941163
transform 1 0 1656 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0845_
timestamp 1667941163
transform 1 0 2024 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0846_
timestamp 1667941163
transform 1 0 11960 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0847_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19504 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0848_
timestamp 1667941163
transform 1 0 13156 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0849_
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0850_
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0851_
timestamp 1667941163
transform 1 0 19780 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0852_
timestamp 1667941163
transform 1 0 19136 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0853_
timestamp 1667941163
transform 1 0 21896 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0854_
timestamp 1667941163
transform 1 0 12236 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0855_
timestamp 1667941163
transform 1 0 16192 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0856_
timestamp 1667941163
transform 1 0 19412 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0857_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11684 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0858_
timestamp 1667941163
transform 1 0 6532 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0862_
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0863_
timestamp 1667941163
transform 1 0 7360 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0864_
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0865_
timestamp 1667941163
transform 1 0 6808 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0866_
timestamp 1667941163
transform 1 0 19228 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 11960 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 14536 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 12328 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0870_
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0871_
timestamp 1667941163
transform 1 0 19780 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0872_
timestamp 1667941163
transform 1 0 22264 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0873_
timestamp 1667941163
transform 1 0 17204 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0874_
timestamp 1667941163
transform 1 0 15088 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 15824 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0878_
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0879_
timestamp 1667941163
transform 1 0 12972 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0880_
timestamp 1667941163
transform 1 0 19596 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0881_
timestamp 1667941163
transform 1 0 15088 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0882_
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 9476 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0885_
timestamp 1667941163
transform 1 0 6716 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 9384 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0887_
timestamp 1667941163
transform 1 0 7176 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0888_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0889_
timestamp 1667941163
transform 1 0 16560 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0890_
timestamp 1667941163
transform 1 0 15088 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 15640 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 9660 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0896_
timestamp 1667941163
transform 1 0 10948 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0897_
timestamp 1667941163
transform 1 0 13156 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0898_
timestamp 1667941163
transform 1 0 11868 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0899_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 6808 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 4232 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0902_
timestamp 1667941163
transform 1 0 7820 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 10580 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0904_
timestamp 1667941163
transform 1 0 8372 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 9752 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 4232 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0909_
timestamp 1667941163
transform 1 0 7176 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 12328 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0911_
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 4232 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0913_
timestamp 1667941163
transform 1 0 6808 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 3956 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 9384 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 19596 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 21988 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 9384 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 4600 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 14996 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0922_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 15916 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 11960 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 6624 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 6072 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0927_
timestamp 1667941163
transform 1 0 11868 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0928_
timestamp 1667941163
transform 1 0 14444 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0929_
timestamp 1667941163
transform 1 0 6808 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 6164 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 4600 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 9384 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0933_
timestamp 1667941163
transform 1 0 1656 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 1656 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0936_
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 4232 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0938_
timestamp 1667941163
transform 1 0 9108 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 11224 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform 1 0 9660 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0943_
timestamp 1667941163
transform 1 0 10212 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0944_
timestamp 1667941163
transform 1 0 7728 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 14536 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0946_
timestamp 1667941163
transform 1 0 12236 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 19504 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0948_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 21988 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0950_
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1667941163
transform 1 0 16928 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 19136 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0954_
timestamp 1667941163
transform 1 0 17940 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0955_
timestamp 1667941163
transform 1 0 12052 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0956_
timestamp 1667941163
transform 1 0 13248 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform 1 0 21620 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform 1 0 9752 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0960_
timestamp 1667941163
transform 1 0 11408 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0961_
timestamp 1667941163
transform 1 0 19504 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0962_
timestamp 1667941163
transform 1 0 19412 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 13064 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1667941163
transform 1 0 33764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 35696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0991_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 24472 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 32108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 35052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 25208 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0996_
timestamp 1667941163
transform 1 0 22356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 12972 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0999_
timestamp 1667941163
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 17480 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1001_
timestamp 1667941163
transform 1 0 23276 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 37352 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 17664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 37812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 36064 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 3956 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 28152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1010_
timestamp 1667941163
transform 1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 14444 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 32936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 2300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1015_
timestamp 1667941163
transform 1 0 2024 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 35512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1018_
timestamp 1667941163
transform 1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 36616 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1022_
timestamp 1667941163
transform 1 0 15732 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 26128 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 25576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 33764 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 26496 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 37812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1030_
timestamp 1667941163
transform 1 0 20516 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 29716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 33764 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 35328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 12512 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 4508 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 3680 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 3864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1667941163
transform 1 0 33304 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1667941163
transform 1 0 31648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1044_
timestamp 1667941163
transform 1 0 33580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1046_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1047_
timestamp 1667941163
transform 1 0 10028 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1047__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1048_
timestamp 1667941163
transform 1 0 14996 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1049_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1050_
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1051_
timestamp 1667941163
transform 1 0 12604 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1052_
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1053_
timestamp 1667941163
transform 1 0 29716 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1054_
timestamp 1667941163
transform 1 0 12420 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1055_
timestamp 1667941163
transform 1 0 27968 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1056_
timestamp 1667941163
transform 1 0 27416 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1057_
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1058_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1059__143
timestamp 1667941163
transform 1 0 22816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 11960 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1061_
timestamp 1667941163
transform 1 0 23460 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1062_
timestamp 1667941163
transform 1 0 9476 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1063_
timestamp 1667941163
transform 1 0 22264 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1064_
timestamp 1667941163
transform 1 0 24840 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1065_
timestamp 1667941163
transform 1 0 15732 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1066_
timestamp 1667941163
transform 1 0 19596 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 10672 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1068_
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1069_
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1070_
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1071_
timestamp 1667941163
transform 1 0 27324 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1071__144
timestamp 1667941163
transform 1 0 27416 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1072_
timestamp 1667941163
transform 1 0 6900 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1073_
timestamp 1667941163
transform 1 0 10580 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1074_
timestamp 1667941163
transform 1 0 7820 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1075_
timestamp 1667941163
transform 1 0 4508 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1076_
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1077_
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1078_
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1079_
timestamp 1667941163
transform 1 0 15088 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1080_
timestamp 1667941163
transform 1 0 23276 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 22816 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1082_
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1083_
timestamp 1667941163
transform 1 0 26036 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1083__145
timestamp 1667941163
transform 1 0 27508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1084_
timestamp 1667941163
transform 1 0 13064 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1085_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1086_
timestamp 1667941163
transform 1 0 11960 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1087_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1088_
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1089_
timestamp 1667941163
transform 1 0 24564 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1090_
timestamp 1667941163
transform 1 0 24932 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1091_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1092_
timestamp 1667941163
transform 1 0 25852 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1093_
timestamp 1667941163
transform 1 0 25024 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1094_
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1095_
timestamp 1667941163
transform 1 0 27232 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1095__146
timestamp 1667941163
transform 1 0 27600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1096_
timestamp 1667941163
transform 1 0 24288 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1097_
timestamp 1667941163
transform 1 0 12604 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1098_
timestamp 1667941163
transform 1 0 1748 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1100_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1101_
timestamp 1667941163
transform 1 0 25852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1102_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1103_
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1104_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1105_
timestamp 1667941163
transform 1 0 13524 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1106_
timestamp 1667941163
transform 1 0 12144 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1107__147
timestamp 1667941163
transform 1 0 14720 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1107_
timestamp 1667941163
transform 1 0 14628 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1108_
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1109_
timestamp 1667941163
transform 1 0 8464 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1110_
timestamp 1667941163
transform 1 0 6624 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1111_
timestamp 1667941163
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1112_
timestamp 1667941163
transform 1 0 19872 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1113_
timestamp 1667941163
transform 1 0 11408 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1114_
timestamp 1667941163
transform 1 0 12604 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1115_
timestamp 1667941163
transform 1 0 22724 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1116_
timestamp 1667941163
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1117_
timestamp 1667941163
transform 1 0 17296 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1118_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1119_
timestamp 1667941163
transform 1 0 20976 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1119__148
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1120_
timestamp 1667941163
transform 1 0 10120 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1121_
timestamp 1667941163
transform 1 0 10396 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1122_
timestamp 1667941163
transform 1 0 18124 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1123_
timestamp 1667941163
transform 1 0 14904 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1124_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1125_
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1126_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 15548 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 17664 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1129__149
timestamp 1667941163
transform 1 0 13156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1129_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12788 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1130_
timestamp 1667941163
transform 1 0 14996 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1131_
timestamp 1667941163
transform 1 0 13616 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 17848 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 7268 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 20424 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 9568 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 12052 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 9568 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1140_
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1141_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1141__150
timestamp 1667941163
transform 1 0 24196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 15548 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1144_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 19044 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1147__151
timestamp 1667941163
transform 1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 11408 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 17296 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1151_
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 17664 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 23828 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1154__152
timestamp 1667941163
transform 1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1154_
timestamp 1667941163
transform 1 0 27140 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1155_
timestamp 1667941163
transform 1 0 4324 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1156_
timestamp 1667941163
transform 1 0 9660 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 23000 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 26312 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1159_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 16192 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1162__153
timestamp 1667941163
transform 1 0 19228 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1162_
timestamp 1667941163
transform 1 0 19872 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1163_
timestamp 1667941163
transform 1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1164_
timestamp 1667941163
transform 1 0 12328 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1165_
timestamp 1667941163
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 14536 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1168__154
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 9108 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 7176 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1170_
timestamp 1667941163
transform 1 0 6716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1171_
timestamp 1667941163
transform 1 0 8832 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1172_
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1172__155
timestamp 1667941163
transform 1 0 4324 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 9660 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 14996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1176__156
timestamp 1667941163
transform 1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 2668 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 6256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform 1 0 3128 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 9108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1180__157
timestamp 1667941163
transform 1 0 2852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1180_
timestamp 1667941163
transform 1 0 2668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1182_
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1183_
timestamp 1667941163
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 12144 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1184__158
timestamp 1667941163
transform 1 0 12328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 10212 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 12052 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1188__159
timestamp 1667941163
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 22724 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 27784 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 28336 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 27140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 22540 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1192__160
timestamp 1667941163
transform 1 0 22632 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1193_
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1195_
timestamp 1667941163
transform 1 0 10580 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 14260 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1197__161
timestamp 1667941163
transform 1 0 13524 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 13800 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1198_
timestamp 1667941163
transform 1 0 15456 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1199_
timestamp 1667941163
transform 1 0 14168 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1200_
timestamp 1667941163
transform 1 0 12696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 16744 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 27692 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1203__162
timestamp 1667941163
transform 1 0 28060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 28336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1204_
timestamp 1667941163
transform 1 0 23552 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1205_
timestamp 1667941163
transform 1 0 26128 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1206_
timestamp 1667941163
transform 1 0 29072 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 26680 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1208_
timestamp 1667941163
transform 1 0 23368 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1209__163
timestamp 1667941163
transform 1 0 22632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 20148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 22908 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 29256 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1215__164
timestamp 1667941163
transform 1 0 30084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 16928 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1217_
timestamp 1667941163
transform 1 0 22632 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 28796 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1219_
timestamp 1667941163
transform 1 0 18124 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1220_
timestamp 1667941163
transform 1 0 22172 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1221_
timestamp 1667941163
transform 1 0 23184 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1222_
timestamp 1667941163
transform 1 0 22356 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1223_
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1223__165
timestamp 1667941163
transform 1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1224_
timestamp 1667941163
transform 1 0 12788 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1225_
timestamp 1667941163
transform 1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1226_
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1227_
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1228_
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1229_
timestamp 1667941163
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 13156 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1231_
timestamp 1667941163
transform 1 0 20240 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1232_
timestamp 1667941163
transform 1 0 28428 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1233_
timestamp 1667941163
transform 1 0 27140 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1234_
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1235__166
timestamp 1667941163
transform 1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1235_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1236_
timestamp 1667941163
transform 1 0 27784 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1237_
timestamp 1667941163
transform 1 0 17204 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1238_
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1239_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1240_
timestamp 1667941163
transform 1 0 24656 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1241_
timestamp 1667941163
transform 1 0 25484 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1242_
timestamp 1667941163
transform 1 0 29716 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1243_
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9384 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 2852 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 6532 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 12512 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 5060 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 5428 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 14444 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 14720 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 17940 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 21988 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 15640 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 17940 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 21804 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 36156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1667941163
transform 1 0 18032 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 32292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform 1 0 37444 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform 1 0 37444 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1667941163
transform 1 0 2576 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1667941163
transform 1 0 2852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1667941163
transform 1 0 37444 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 38088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 38088 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 38088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 2944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 36708 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 28980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 36708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1667941163
transform 1 0 33580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1667941163
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1667941163
transform 1 0 2668 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 16100 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 35512 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 30360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 34868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 1564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 31004 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 2 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 3 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 ccff_head
port 4 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 82 nsew signal input
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 83 nsew signal input
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 84 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 85 nsew signal input
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 86 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 87 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_bottom_in[15]
port 88 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 89 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 90 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_bottom_in[18]
port 91 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 92 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 93 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 94 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 95 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 96 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 97 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 98 nsew signal input
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 99 nsew signal input
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 100 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 101 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 102 nsew signal tristate
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 103 nsew signal tristate
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 104 nsew signal tristate
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 105 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 106 nsew signal tristate
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_bottom_out[15]
port 107 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_bottom_out[16]
port 108 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_bottom_out[17]
port 109 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 110 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 111 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_bottom_out[2]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 113 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 114 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 115 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 116 nsew signal tristate
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 117 nsew signal tristate
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 118 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 119 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 120 nsew signal input
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 121 nsew signal input
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 122 nsew signal input
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 123 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 124 nsew signal input
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 125 nsew signal input
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 126 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 pReset
port 130 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 prog_clk
port 131 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 132 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 133 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 138 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 139 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 140 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 141 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 vssd1
port 143 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 3174 14790 3174 14790 0 _0000_
rlabel metal1 8464 13158 8464 13158 0 _0001_
rlabel metal1 15502 13362 15502 13362 0 _0002_
rlabel metal1 18722 14790 18722 14790 0 _0003_
rlabel metal1 21988 13158 21988 13158 0 _0004_
rlabel metal1 8740 13838 8740 13838 0 _0005_
rlabel metal1 15962 11621 15962 11621 0 _0006_
rlabel metal1 8280 13702 8280 13702 0 _0007_
rlabel via3 18285 6868 18285 6868 0 _0008_
rlabel metal2 10902 8942 10902 8942 0 _0009_
rlabel metal3 13087 9588 13087 9588 0 _0010_
rlabel metal3 11868 12580 11868 12580 0 _0011_
rlabel metal1 5382 14042 5382 14042 0 _0012_
rlabel metal1 7084 14790 7084 14790 0 _0013_
rlabel metal1 5336 13158 5336 13158 0 _0014_
rlabel metal1 6578 10744 6578 10744 0 _0015_
rlabel metal1 8004 11866 8004 11866 0 _0016_
rlabel metal3 4761 14620 4761 14620 0 _0017_
rlabel metal1 19143 2346 19143 2346 0 _0018_
rlabel metal1 20838 2455 20838 2455 0 _0019_
rlabel metal1 13662 4488 13662 4488 0 _0020_
rlabel metal2 6118 12852 6118 12852 0 _0021_
rlabel metal1 11776 10438 11776 10438 0 _0022_
rlabel metal2 7682 14144 7682 14144 0 _0023_
rlabel metal2 5934 9112 5934 9112 0 _0024_
rlabel metal2 3588 12036 3588 12036 0 _0025_
rlabel metal3 8027 10268 8027 10268 0 _0026_
rlabel metal3 6233 15572 6233 15572 0 _0027_
rlabel metal1 10442 14246 10442 14246 0 _0028_
rlabel metal1 21022 10071 21022 10071 0 _0029_
rlabel metal2 29854 4352 29854 4352 0 _0030_
rlabel metal1 21213 4590 21213 4590 0 _0031_
rlabel metal1 32982 2822 32982 2822 0 _0032_
rlabel metal1 6447 3502 6447 3502 0 _0033_
rlabel metal1 17119 4590 17119 4590 0 _0034_
rlabel metal1 20983 3502 20983 3502 0 _0035_
rlabel metal1 16146 9486 16146 9486 0 _0036_
rlabel metal2 9246 13804 9246 13804 0 _0037_
rlabel metal1 8333 5610 8333 5610 0 _0038_
rlabel metal1 5796 13362 5796 13362 0 _0039_
rlabel metal2 12650 10234 12650 10234 0 _0040_
rlabel metal2 15686 13838 15686 13838 0 _0041_
rlabel metal1 7452 10438 7452 10438 0 _0042_
rlabel metal1 3174 15946 3174 15946 0 _0043_
rlabel metal1 3312 15334 3312 15334 0 _0044_
rlabel metal2 4002 13328 4002 13328 0 _0045_
rlabel metal1 4048 16422 4048 16422 0 _0046_
rlabel metal1 2668 14790 2668 14790 0 _0047_
rlabel metal1 4009 3434 4009 3434 0 _0048_
rlabel metal1 8740 6834 8740 6834 0 _0049_
rlabel metal2 5014 9758 5014 9758 0 _0050_
rlabel metal3 4991 15300 4991 15300 0 _0051_
rlabel metal1 22218 6086 22218 6086 0 _0052_
rlabel metal1 16921 9622 16921 9622 0 _0053_
rlabel metal2 12466 11764 12466 11764 0 _0054_
rlabel metal2 6854 11271 6854 11271 0 _0055_
rlabel metal1 7406 10234 7406 10234 0 _0056_
rlabel metal1 8411 7446 8411 7446 0 _0057_
rlabel metal1 18630 12920 18630 12920 0 _0058_
rlabel metal2 13662 6086 13662 6086 0 _0059_
rlabel metal1 20700 12614 20700 12614 0 _0060_
rlabel metal1 18775 10710 18775 10710 0 _0061_
rlabel metal1 21206 14824 21206 14824 0 _0062_
rlabel metal1 18860 10166 18860 10166 0 _0063_
rlabel metal1 21298 11016 21298 11016 0 _0064_
rlabel metal2 20240 4182 20240 4182 0 _0065_
rlabel metal1 21489 6698 21489 6698 0 _0066_
rlabel metal1 20339 12886 20339 12886 0 _0067_
rlabel metal1 12788 10778 12788 10778 0 _0068_
rlabel metal1 14352 9146 14352 9146 0 _0069_
rlabel metal1 20010 3128 20010 3128 0 _0070_
rlabel metal1 23046 4631 23046 4631 0 _0071_
rlabel metal2 12466 3740 12466 3740 0 _0072_
rlabel metal4 12788 13940 12788 13940 0 _0073_
rlabel metal2 25898 6919 25898 6919 0 _0074_
rlabel metal1 21512 6358 21512 6358 0 _0075_
rlabel metal1 10672 2822 10672 2822 0 _0076_
rlabel metal1 3641 2346 3641 2346 0 _0077_
rlabel metal3 15272 1700 15272 1700 0 _0078_
rlabel metal1 13386 4699 13386 4699 0 _0079_
rlabel metal1 26450 5814 26450 5814 0 _0080_
rlabel metal1 13800 12138 13800 12138 0 _0081_
rlabel metal2 21114 11169 21114 11169 0 _0082_
rlabel metal1 28474 3366 28474 3366 0 _0083_
rlabel metal1 30544 4114 30544 4114 0 _0084_
rlabel metal1 33488 2890 33488 2890 0 _0085_
rlabel metal1 25944 5882 25944 5882 0 _0086_
rlabel metal3 16905 9996 16905 9996 0 _0087_
rlabel metal1 19826 15674 19826 15674 0 _0088_
rlabel metal1 25438 5746 25438 5746 0 _0089_
rlabel metal1 13255 4182 13255 4182 0 _0090_
rlabel metal1 9338 4216 9338 4216 0 _0091_
rlabel metal1 13623 2346 13623 2346 0 _0092_
rlabel metal1 8234 2523 8234 2523 0 _0093_
rlabel metal1 5849 2346 5849 2346 0 _0094_
rlabel via2 6854 3077 6854 3077 0 _0095_
rlabel metal2 8142 11849 8142 11849 0 _0096_
rlabel metal1 6302 11594 6302 11594 0 _0097_
rlabel metal3 5474 12580 5474 12580 0 _0098_
rlabel metal1 22356 13158 22356 13158 0 _0099_
rlabel metal1 13531 3434 13531 3434 0 _0100_
rlabel metal2 32430 1972 32430 1972 0 _0101_
rlabel metal2 13754 2771 13754 2771 0 _0102_
rlabel metal1 11553 2346 11553 2346 0 _0103_
rlabel metal1 21351 8874 21351 8874 0 _0104_
rlabel metal1 24111 8942 24111 8942 0 _0105_
rlabel metal1 24610 5338 24610 5338 0 _0106_
rlabel metal2 16514 6409 16514 6409 0 _0107_
rlabel metal1 17671 3434 17671 3434 0 _0108_
rlabel metal1 16705 2346 16705 2346 0 _0109_
rlabel metal2 16514 2941 16514 2941 0 _0110_
rlabel metal2 34546 2040 34546 2040 0 _0111_
rlabel metal2 20470 7242 20470 7242 0 _0112_
rlabel metal1 22639 9622 22639 9622 0 _0113_
rlabel metal1 29072 5882 29072 5882 0 _0114_
rlabel metal2 21114 4505 21114 4505 0 _0115_
rlabel metal1 7268 11526 7268 11526 0 _0116_
rlabel metal1 7636 12614 7636 12614 0 _0117_
rlabel metal1 8517 8874 8517 8874 0 _0118_
rlabel metal2 9338 9469 9338 9469 0 _0119_
rlabel metal1 23736 9554 23736 9554 0 _0120_
rlabel metal1 19734 14994 19734 14994 0 _0121_
rlabel metal1 8234 15062 8234 15062 0 _0122_
rlabel metal2 17066 11322 17066 11322 0 _0123_
rlabel metal1 32890 3026 32890 3026 0 _0124_
rlabel metal1 7222 14382 7222 14382 0 _0125_
rlabel metal1 14950 14314 14950 14314 0 _0126_
rlabel metal1 20056 12818 20056 12818 0 _0127_
rlabel metal1 20930 12818 20930 12818 0 _0128_
rlabel metal2 17250 25738 17250 25738 0 _0129_
rlabel metal2 27278 14586 27278 14586 0 _0130_
rlabel metal1 28934 15028 28934 15028 0 _0131_
rlabel metal2 21482 20026 21482 20026 0 _0132_
rlabel metal2 24610 21556 24610 21556 0 _0133_
rlabel metal1 23414 24752 23414 24752 0 _0134_
rlabel metal2 23782 19210 23782 19210 0 _0135_
rlabel metal2 27738 18122 27738 18122 0 _0136_
rlabel metal2 28750 19788 28750 19788 0 _0137_
rlabel metal1 15456 26350 15456 26350 0 _0138_
rlabel metal1 13294 25874 13294 25874 0 _0139_
rlabel metal2 13754 26554 13754 26554 0 _0140_
rlabel metal1 7590 19482 7590 19482 0 _0141_
rlabel metal2 21482 22780 21482 22780 0 _0142_
rlabel metal1 29900 6766 29900 6766 0 _0143_
rlabel metal2 32522 5338 32522 5338 0 _0144_
rlabel metal2 8602 23290 8602 23290 0 _0145_
rlabel metal2 10166 24378 10166 24378 0 _0146_
rlabel metal2 5014 16422 5014 16422 0 _0147_
rlabel metal1 2300 9690 2300 9690 0 _0148_
rlabel metal2 5842 18564 5842 18564 0 _0149_
rlabel metal2 2714 16388 2714 16388 0 _0150_
rlabel metal1 11316 17850 11316 17850 0 _0151_
rlabel metal2 4738 18938 4738 18938 0 _0152_
rlabel metal1 6256 18938 6256 18938 0 _0153_
rlabel metal1 7176 22406 7176 22406 0 _0154_
rlabel metal1 13018 16048 13018 16048 0 _0155_
rlabel metal2 11592 7718 11592 7718 0 _0156_
rlabel metal1 29532 4114 29532 4114 0 _0157_
rlabel metal2 20194 14280 20194 14280 0 _0158_
rlabel metal2 14490 13719 14490 13719 0 _0159_
rlabel metal1 18400 13974 18400 13974 0 _0160_
rlabel metal3 7360 13532 7360 13532 0 _0161_
rlabel metal1 15410 16490 15410 16490 0 _0162_
rlabel metal1 17020 18326 17020 18326 0 _0163_
rlabel metal1 15318 15096 15318 15096 0 _0164_
rlabel metal1 13202 19754 13202 19754 0 _0165_
rlabel metal1 16468 13226 16468 13226 0 _0166_
rlabel metal1 29946 12104 29946 12104 0 _0167_
rlabel metal2 13478 12648 13478 12648 0 _0168_
rlabel metal2 28198 13736 28198 13736 0 _0169_
rlabel metal1 27600 15130 27600 15130 0 _0170_
rlabel metal2 21206 13158 21206 13158 0 _0171_
rlabel metal1 27738 14042 27738 14042 0 _0172_
rlabel metal2 22954 15912 22954 15912 0 _0173_
rlabel metal1 8671 15946 8671 15946 0 _0174_
rlabel metal2 23690 9214 23690 9214 0 _0175_
rlabel metal2 9890 17459 9890 17459 0 _0176_
rlabel metal1 23920 3094 23920 3094 0 _0177_
rlabel metal1 25162 17306 25162 17306 0 _0178_
rlabel metal1 16928 20570 16928 20570 0 _0179_
rlabel metal2 19826 13311 19826 13311 0 _0180_
rlabel metal2 6946 14654 6946 14654 0 _0181_
rlabel metal1 24656 2074 24656 2074 0 _0182_
rlabel metal2 14214 14280 14214 14280 0 _0183_
rlabel metal1 14030 15402 14030 15402 0 _0184_
rlabel metal2 28382 9112 28382 9112 0 _0185_
rlabel metal2 8050 20264 8050 20264 0 _0186_
rlabel metal1 10028 22950 10028 22950 0 _0187_
rlabel metal1 6716 10778 6716 10778 0 _0188_
rlabel metal1 5980 17510 5980 17510 0 _0189_
rlabel metal1 10534 22440 10534 22440 0 _0190_
rlabel metal1 24380 13974 24380 13974 0 _0191_
rlabel metal1 18216 9146 18216 9146 0 _0192_
rlabel metal2 15272 21556 15272 21556 0 _0193_
rlabel metal2 23506 22814 23506 22814 0 _0194_
rlabel metal2 23046 11934 23046 11934 0 _0195_
rlabel metal2 30406 3995 30406 3995 0 _0196_
rlabel metal1 26772 7514 26772 7514 0 _0197_
rlabel metal1 13294 16184 13294 16184 0 _0198_
rlabel metal1 22540 17850 22540 17850 0 _0199_
rlabel metal1 11546 19414 11546 19414 0 _0200_
rlabel metal1 24794 4488 24794 4488 0 _0201_
rlabel metal1 25852 17850 25852 17850 0 _0202_
rlabel metal2 24794 5848 24794 5848 0 _0203_
rlabel metal1 25254 6698 25254 6698 0 _0204_
rlabel metal1 22356 15062 22356 15062 0 _0205_
rlabel metal1 26128 16762 26128 16762 0 _0206_
rlabel metal2 25254 8670 25254 8670 0 _0207_
rlabel metal1 22862 4182 22862 4182 0 _0208_
rlabel metal1 27140 12886 27140 12886 0 _0209_
rlabel metal2 24518 16286 24518 16286 0 _0210_
rlabel metal1 12834 14280 12834 14280 0 _0211_
rlabel metal1 2208 12410 2208 12410 0 _0212_
rlabel metal2 18998 15096 18998 15096 0 _0213_
rlabel metal1 27370 18360 27370 18360 0 _0214_
rlabel metal2 26082 15368 26082 15368 0 _0215_
rlabel metal1 24794 13192 24794 13192 0 _0216_
rlabel metal1 25852 6358 25852 6358 0 _0217_
rlabel metal1 27232 12410 27232 12410 0 _0218_
rlabel metal1 8372 16966 8372 16966 0 _0219_
rlabel metal2 8510 22678 8510 22678 0 _0220_
rlabel metal1 8372 16218 8372 16218 0 _0221_
rlabel metal1 15456 19414 15456 19414 0 _0222_
rlabel metal2 8694 20910 8694 20910 0 _0223_
rlabel metal2 6854 15130 6854 15130 0 _0224_
rlabel metal1 19872 15402 19872 15402 0 _0225_
rlabel metal1 18906 20502 18906 20502 0 _0226_
rlabel metal1 10718 19482 10718 19482 0 _0227_
rlabel metal1 11822 18292 11822 18292 0 _0228_
rlabel metal1 22954 14280 22954 14280 0 _0229_
rlabel metal1 14812 17850 14812 17850 0 _0230_
rlabel metal1 12052 13906 12052 13906 0 _0231_
rlabel metal1 19504 20026 19504 20026 0 _0232_
rlabel metal1 21114 15062 21114 15062 0 _0233_
rlabel metal1 10212 20502 10212 20502 0 _0234_
rlabel metal1 10994 22678 10994 22678 0 _0235_
rlabel metal1 18400 21930 18400 21930 0 _0236_
rlabel metal1 14766 22746 14766 22746 0 _0237_
rlabel metal1 17020 24854 17020 24854 0 _0238_
rlabel metal2 18354 23528 18354 23528 0 _0239_
rlabel metal2 13662 15606 13662 15606 0 _0240_
rlabel metal2 15778 23630 15778 23630 0 _0241_
rlabel metal1 17526 23766 17526 23766 0 _0242_
rlabel metal1 12926 20570 12926 20570 0 _0243_
rlabel metal1 14674 16422 14674 16422 0 _0244_
rlabel metal2 12742 21012 12742 21012 0 _0245_
rlabel metal2 18078 17646 18078 17646 0 _0246_
rlabel metal1 7360 17238 7360 17238 0 _0247_
rlabel metal2 20654 17000 20654 17000 0 _0248_
rlabel metal1 8832 18598 8832 18598 0 _0249_
rlabel metal1 11546 23154 11546 23154 0 _0250_
rlabel metal2 10718 17646 10718 17646 0 _0251_
rlabel metal1 10580 17238 10580 17238 0 _0252_
rlabel metal1 9844 22406 9844 22406 0 _0253_
rlabel metal1 25760 11594 25760 11594 0 _0254_
rlabel metal2 24978 7650 24978 7650 0 _0255_
rlabel metal2 11454 17646 11454 17646 0 _0256_
rlabel viali 15774 18326 15774 18326 0 _0257_
rlabel metal1 19642 14280 19642 14280 0 _0258_
rlabel metal1 19044 16762 19044 16762 0 _0259_
rlabel metal1 6072 11798 6072 11798 0 _0260_
rlabel metal2 5106 15912 5106 15912 0 _0261_
rlabel metal2 9430 16439 9430 16439 0 _0262_
rlabel metal1 16882 16218 16882 16218 0 _0263_
rlabel metal1 9338 15062 9338 15062 0 _0264_
rlabel metal1 17434 16490 17434 16490 0 _0265_
rlabel metal2 17894 15640 17894 15640 0 _0266_
rlabel metal1 25438 4182 25438 4182 0 _0267_
rlabel metal2 33074 3536 33074 3536 0 _0268_
rlabel metal1 4646 14314 4646 14314 0 _0269_
rlabel metal1 9844 13226 9844 13226 0 _0270_
rlabel metal1 23644 7446 23644 7446 0 _0271_
rlabel metal2 27922 7072 27922 7072 0 _0272_
rlabel metal1 27140 11322 27140 11322 0 _0273_
rlabel metal1 16652 19890 16652 19890 0 _0274_
rlabel metal2 8740 19320 8740 19320 0 _0275_
rlabel metal1 18538 13838 18538 13838 0 _0276_
rlabel metal1 15456 18802 15456 18802 0 _0277_
rlabel metal2 12558 19074 12558 19074 0 _0278_
rlabel metal1 13524 20978 13524 20978 0 _0279_
rlabel metal1 11362 20536 11362 20536 0 _0280_
rlabel metal1 14904 20978 14904 20978 0 _0281_
rlabel metal1 7222 21862 7222 21862 0 _0282_
rlabel metal1 7130 17714 7130 17714 0 _0283_
rlabel metal2 6946 20536 6946 20536 0 _0284_
rlabel metal1 8188 18938 8188 18938 0 _0285_
rlabel metal2 4370 18462 4370 18462 0 _0286_
rlabel metal2 16882 17238 16882 17238 0 _0287_
rlabel metal2 9706 17374 9706 17374 0 _0288_
rlabel metal1 13846 17000 13846 17000 0 _0289_
rlabel metal2 2898 15368 2898 15368 0 _0290_
rlabel metal2 6486 17068 6486 17068 0 _0291_
rlabel metal2 3358 15470 3358 15470 0 _0292_
rlabel metal2 6302 16286 6302 16286 0 _0293_
rlabel metal2 2530 10404 2530 10404 0 _0294_
rlabel metal2 5474 16558 5474 16558 0 _0295_
rlabel metal2 1978 10404 1978 10404 0 _0296_
rlabel metal1 21620 11798 21620 11798 0 _0297_
rlabel metal1 11914 21590 11914 21590 0 _0298_
rlabel metal1 10534 21522 10534 21522 0 _0299_
rlabel metal1 9936 23766 9936 23766 0 _0300_
rlabel metal1 12236 22542 12236 22542 0 _0301_
rlabel metal2 27554 4624 27554 4624 0 _0302_
rlabel metal1 28888 6834 28888 6834 0 _0303_
rlabel metal2 28566 5440 28566 5440 0 _0304_
rlabel metal1 28198 8398 28198 8398 0 _0305_
rlabel metal1 22402 22406 22402 22406 0 _0306_
rlabel metal1 6210 20808 6210 20808 0 _0307_
rlabel metal2 19642 21080 19642 21080 0 _0308_
rlabel metal1 9660 18394 9660 18394 0 _0309_
rlabel metal2 14490 24888 14490 24888 0 _0310_
rlabel metal2 14030 25092 14030 25092 0 _0311_
rlabel metal1 15640 24242 15640 24242 0 _0312_
rlabel metal2 14398 25568 14398 25568 0 _0313_
rlabel metal1 13432 23630 13432 23630 0 _0314_
rlabel metal2 16974 24412 16974 24412 0 _0315_
rlabel metal2 27922 17374 27922 17374 0 _0316_
rlabel metal2 28566 18700 28566 18700 0 _0317_
rlabel metal2 23782 18428 23782 18428 0 _0318_
rlabel metal2 26358 18088 26358 18088 0 _0319_
rlabel metal2 29302 17340 29302 17340 0 _0320_
rlabel metal1 27738 19890 27738 19890 0 _0321_
rlabel metal2 23782 21692 23782 21692 0 _0322_
rlabel metal2 22862 24140 22862 24140 0 _0323_
rlabel metal1 20838 19890 20838 19890 0 _0324_
rlabel metal2 24150 20740 24150 20740 0 _0325_
rlabel metal1 20056 22610 20056 22610 0 _0326_
rlabel metal1 20976 20978 20976 20978 0 _0327_
rlabel metal1 28612 13974 28612 13974 0 _0328_
rlabel metal2 30222 14620 30222 14620 0 _0329_
rlabel metal2 17158 23902 17158 23902 0 _0330_
rlabel metal1 22862 15368 22862 15368 0 _0331_
rlabel metal1 28704 12410 28704 12410 0 _0332_
rlabel metal2 18354 25432 18354 25432 0 _0333_
rlabel metal1 23552 12138 23552 12138 0 _0334_
rlabel metal1 23598 9962 23598 9962 0 _0335_
rlabel metal2 22586 18904 22586 18904 0 _0336_
rlabel metal2 24886 18462 24886 18462 0 _0337_
rlabel metal1 12880 16490 12880 16490 0 _0338_
rlabel metal2 22218 16728 22218 16728 0 _0339_
rlabel metal2 20378 17374 20378 17374 0 _0340_
rlabel metal1 23920 15062 23920 15062 0 _0341_
rlabel metal1 23690 12886 23690 12886 0 _0342_
rlabel metal1 16054 17238 16054 17238 0 _0343_
rlabel metal2 13386 16558 13386 16558 0 _0344_
rlabel metal2 20470 17646 20470 17646 0 _0345_
rlabel metal2 31602 6528 31602 6528 0 _0346_
rlabel metal1 27370 5304 27370 5304 0 _0347_
rlabel metal1 13202 18326 13202 18326 0 _0348_
rlabel metal1 19228 18666 19228 18666 0 _0349_
rlabel metal1 27646 10710 27646 10710 0 _0350_
rlabel metal2 17434 16286 17434 16286 0 _0351_
rlabel metal1 24518 17238 24518 17238 0 _0352_
rlabel metal2 17066 15198 17066 15198 0 _0353_
rlabel metal2 24886 9758 24886 9758 0 _0354_
rlabel metal2 29302 3808 29302 3808 0 _0355_
rlabel metal2 29946 9826 29946 9826 0 _0356_
rlabel metal1 18584 12138 18584 12138 0 _0357_
rlabel metal3 1234 19108 1234 19108 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 2806 7701 2806 7701 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal1 5336 37230 5336 37230 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 2990 7769 2990 7769 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal1 36133 3026 36133 3026 0 ccff_head
rlabel metal2 25806 1520 25806 1520 0 ccff_tail
rlabel metal3 1188 22508 1188 22508 0 chanx_left_in[0]
rlabel metal3 1142 6868 1142 6868 0 chanx_left_in[10]
rlabel metal1 18216 37230 18216 37230 0 chanx_left_in[11]
rlabel metal3 1142 38828 1142 38828 0 chanx_left_in[12]
rlabel metal1 15502 3706 15502 3706 0 chanx_left_in[13]
rlabel metal2 29026 1588 29026 1588 0 chanx_left_in[14]
rlabel metal1 25852 37230 25852 37230 0 chanx_left_in[15]
rlabel metal1 6210 37298 6210 37298 0 chanx_left_in[16]
rlabel metal2 32522 3553 32522 3553 0 chanx_left_in[17]
rlabel metal1 9200 36754 9200 36754 0 chanx_left_in[18]
rlabel metal2 20010 1214 20010 1214 0 chanx_left_in[1]
rlabel metal3 1142 17068 1142 17068 0 chanx_left_in[2]
rlabel metal3 1740 2108 1740 2108 0 chanx_left_in[3]
rlabel metal1 27784 37298 27784 37298 0 chanx_left_in[4]
rlabel metal2 11638 1299 11638 1299 0 chanx_left_in[5]
rlabel metal2 38134 32215 38134 32215 0 chanx_left_in[6]
rlabel metal2 38318 27353 38318 27353 0 chanx_left_in[7]
rlabel metal2 9706 1571 9706 1571 0 chanx_left_in[8]
rlabel metal3 1303 748 1303 748 0 chanx_left_in[9]
rlabel metal2 38226 8857 38226 8857 0 chanx_left_out[0]
rlabel metal1 14996 37094 14996 37094 0 chanx_left_out[10]
rlabel metal2 38226 30617 38226 30617 0 chanx_left_out[11]
rlabel metal2 38226 28815 38226 28815 0 chanx_left_out[12]
rlabel metal1 32384 37094 32384 37094 0 chanx_left_out[13]
rlabel metal2 18078 1761 18078 1761 0 chanx_left_out[14]
rlabel metal1 36248 37094 36248 37094 0 chanx_left_out[15]
rlabel metal2 38226 12461 38226 12461 0 chanx_left_out[16]
rlabel metal2 33534 1520 33534 1520 0 chanx_left_out[17]
rlabel metal3 1234 30668 1234 30668 0 chanx_left_out[18]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_out[1]
rlabel metal2 38226 2737 38226 2737 0 chanx_left_out[2]
rlabel metal1 20148 37094 20148 37094 0 chanx_left_out[3]
rlabel via2 38226 35445 38226 35445 0 chanx_left_out[4]
rlabel metal1 36662 2550 36662 2550 0 chanx_left_out[5]
rlabel metal1 19504 36890 19504 36890 0 chanx_left_out[6]
rlabel metal2 34178 1520 34178 1520 0 chanx_left_out[7]
rlabel metal1 31096 37094 31096 37094 0 chanx_left_out[8]
rlabel metal1 34822 37094 34822 37094 0 chanx_left_out[9]
rlabel metal2 38134 37145 38134 37145 0 chanx_right_in[0]
rlabel via1 16606 37179 16606 37179 0 chanx_right_in[10]
rlabel metal2 38318 11033 38318 11033 0 chanx_right_in[11]
rlabel metal1 37352 13838 37352 13838 0 chanx_right_in[12]
rlabel metal2 38134 19227 38134 19227 0 chanx_right_in[13]
rlabel metal2 27738 1588 27738 1588 0 chanx_right_in[14]
rlabel metal3 38786 38828 38786 38828 0 chanx_right_in[15]
rlabel metal2 38134 32759 38134 32759 0 chanx_right_in[16]
rlabel metal1 24610 37230 24610 37230 0 chanx_right_in[17]
rlabel metal1 12512 37230 12512 37230 0 chanx_right_in[18]
rlabel metal2 37490 24021 37490 24021 0 chanx_right_in[1]
rlabel metal1 8786 37298 8786 37298 0 chanx_right_in[2]
rlabel metal1 11776 37230 11776 37230 0 chanx_right_in[3]
rlabel metal1 22632 37298 22632 37298 0 chanx_right_in[4]
rlabel metal1 2622 5610 2622 5610 0 chanx_right_in[5]
rlabel metal1 2898 37230 2898 37230 0 chanx_right_in[6]
rlabel metal1 37352 15470 37352 15470 0 chanx_right_in[7]
rlabel metal1 3956 37298 3956 37298 0 chanx_right_in[8]
rlabel metal2 37490 1921 37490 1921 0 chanx_right_in[9]
rlabel metal3 1234 14348 1234 14348 0 chanx_right_out[0]
rlabel metal2 38226 7633 38226 7633 0 chanx_right_out[10]
rlabel metal3 1234 28628 1234 28628 0 chanx_right_out[11]
rlabel metal1 17250 5814 17250 5814 0 chanx_right_out[12]
rlabel metal3 1234 21148 1234 21148 0 chanx_right_out[13]
rlabel metal2 16146 1163 16146 1163 0 chanx_right_out[14]
rlabel metal3 1234 24548 1234 24548 0 chanx_right_out[15]
rlabel metal1 33212 37094 33212 37094 0 chanx_right_out[16]
rlabel metal3 1234 32708 1234 32708 0 chanx_right_out[17]
rlabel metal2 30314 1520 30314 1520 0 chanx_right_out[18]
rlabel metal2 38226 25177 38226 25177 0 chanx_right_out[1]
rlabel via2 38226 5525 38226 5525 0 chanx_right_out[2]
rlabel metal1 26496 37094 26496 37094 0 chanx_right_out[3]
rlabel metal1 38410 36346 38410 36346 0 chanx_right_out[4]
rlabel metal1 37536 37094 37536 37094 0 chanx_right_out[5]
rlabel metal2 690 2880 690 2880 0 chanx_right_out[6]
rlabel metal1 4462 6086 4462 6086 0 chanx_right_out[7]
rlabel metal2 38686 1792 38686 1792 0 chanx_right_out[8]
rlabel metal3 1234 13668 1234 13668 0 chanx_right_out[9]
rlabel metal2 38318 21913 38318 21913 0 chany_bottom_in[0]
rlabel metal2 38318 15895 38318 15895 0 chany_bottom_in[10]
rlabel metal1 16928 36754 16928 36754 0 chany_bottom_in[11]
rlabel metal1 2438 6732 2438 6732 0 chany_bottom_in[12]
rlabel metal2 38318 3791 38318 3791 0 chany_bottom_in[13]
rlabel metal2 38318 17119 38318 17119 0 chany_bottom_in[14]
rlabel metal3 1234 27268 1234 27268 0 chany_bottom_in[15]
rlabel metal1 2254 36754 2254 36754 0 chany_bottom_in[16]
rlabel metal3 1234 25908 1234 25908 0 chany_bottom_in[17]
rlabel metal3 1234 20468 1234 20468 0 chany_bottom_in[18]
rlabel metal3 1924 39508 1924 39508 0 chany_bottom_in[1]
rlabel metal1 37812 35734 37812 35734 0 chany_bottom_in[2]
rlabel metal1 8510 4590 8510 4590 0 chany_bottom_in[3]
rlabel metal3 1234 17748 1234 17748 0 chany_bottom_in[4]
rlabel metal1 29210 3060 29210 3060 0 chany_bottom_in[5]
rlabel metal2 37398 2132 37398 2132 0 chany_bottom_in[6]
rlabel metal1 13938 37230 13938 37230 0 chany_bottom_in[7]
rlabel metal1 32890 4114 32890 4114 0 chany_bottom_in[8]
rlabel metal1 4416 3910 4416 3910 0 chany_bottom_in[9]
rlabel metal1 14674 4454 14674 4454 0 chany_bottom_out[0]
rlabel metal2 38226 4301 38226 4301 0 chany_bottom_out[10]
rlabel metal2 38226 29393 38226 29393 0 chany_bottom_out[11]
rlabel metal2 38226 20621 38226 20621 0 chany_bottom_out[12]
rlabel metal2 32246 1520 32246 1520 0 chany_bottom_out[13]
rlabel metal3 1234 23868 1234 23868 0 chany_bottom_out[14]
rlabel metal2 38226 10353 38226 10353 0 chany_bottom_out[15]
rlabel metal3 1234 32028 1234 32028 0 chany_bottom_out[16]
rlabel via2 38226 22491 38226 22491 0 chany_bottom_out[17]
rlabel metal2 38226 34221 38226 34221 0 chany_bottom_out[18]
rlabel metal2 36754 1520 36754 1520 0 chany_bottom_out[1]
rlabel metal2 38226 36057 38226 36057 0 chany_bottom_out[2]
rlabel metal3 1234 12308 1234 12308 0 chany_bottom_out[3]
rlabel metal3 1234 34068 1234 34068 0 chany_bottom_out[4]
rlabel metal2 2898 4777 2898 4777 0 chany_bottom_out[5]
rlabel metal2 46 3152 46 3152 0 chany_bottom_out[6]
rlabel metal2 2806 5151 2806 5151 0 chany_bottom_out[7]
rlabel metal2 1794 37179 1794 37179 0 chany_bottom_out[8]
rlabel metal1 10488 37094 10488 37094 0 chany_bottom_out[9]
rlabel metal2 15686 14178 15686 14178 0 clknet_0_prog_clk
rlabel metal1 6716 2482 6716 2482 0 clknet_4_0_0_prog_clk
rlabel metal1 19320 2482 19320 2482 0 clknet_4_10_0_prog_clk
rlabel metal2 16882 6800 16882 6800 0 clknet_4_11_0_prog_clk
rlabel metal2 13294 10370 13294 10370 0 clknet_4_12_0_prog_clk
rlabel metal2 15686 12614 15686 12614 0 clknet_4_13_0_prog_clk
rlabel metal1 16192 7922 16192 7922 0 clknet_4_14_0_prog_clk
rlabel metal1 19734 11220 19734 11220 0 clknet_4_15_0_prog_clk
rlabel metal1 6854 6324 6854 6324 0 clknet_4_1_0_prog_clk
rlabel metal1 9614 2482 9614 2482 0 clknet_4_2_0_prog_clk
rlabel metal2 12282 6528 12282 6528 0 clknet_4_3_0_prog_clk
rlabel metal2 4646 8092 4646 8092 0 clknet_4_4_0_prog_clk
rlabel metal1 6578 9554 6578 9554 0 clknet_4_5_0_prog_clk
rlabel metal1 7222 8534 7222 8534 0 clknet_4_6_0_prog_clk
rlabel metal1 11178 12614 11178 12614 0 clknet_4_7_0_prog_clk
rlabel metal2 14582 3808 14582 3808 0 clknet_4_8_0_prog_clk
rlabel metal2 15134 5406 15134 5406 0 clknet_4_9_0_prog_clk
rlabel metal2 23506 36924 23506 36924 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal3 1234 29308 1234 29308 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 6118 8942 6118 8942 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 1978 4070 1978 4070 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel via2 2898 8925 2898 8925 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 21758 37230 21758 37230 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 19366 1707 19366 1707 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 35604 36754 35604 36754 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 38786 6868 38786 6868 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 36108 1234 36108 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 12374 20434 12374 20434 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal1 13938 12614 13938 12614 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal3 9177 15300 9177 15300 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal3 15709 18020 15709 18020 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal2 18446 2142 18446 2142 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal1 20378 2618 20378 2618 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 19872 3434 19872 3434 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal1 9890 12750 9890 12750 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal1 10718 7718 10718 7718 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal1 7222 18258 7222 18258 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal1 5842 16592 5842 16592 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal1 2898 16048 2898 16048 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal1 2024 3570 2024 3570 0 mem_bottom_track_15.DFFR_0_.Q
rlabel metal1 2070 9588 2070 9588 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal1 10948 5746 10948 5746 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal3 8349 18836 8349 18836 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal1 14030 17646 14030 17646 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal3 12811 17204 12811 17204 0 mem_bottom_track_19.DFFR_1_.Q
rlabel via1 18630 8330 18630 8330 0 mem_bottom_track_21.DFFR_0_.Q
rlabel metal1 30590 6324 30590 6324 0 mem_bottom_track_21.DFFR_1_.Q
rlabel metal1 16192 19346 16192 19346 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal2 16422 12852 16422 12852 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal2 22770 23970 22770 23970 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 21298 11968 21298 11968 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 19688 11662 19688 11662 0 mem_bottom_track_27.DFFR_0_.Q
rlabel metal1 11178 10166 11178 10166 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal1 15824 4658 15824 4658 0 mem_bottom_track_3.DFFR_0_.Q
rlabel via3 17963 15300 17963 15300 0 mem_bottom_track_3.DFFR_1_.Q
rlabel metal3 7015 15300 7015 15300 0 mem_bottom_track_3.DFFR_2_.Q
rlabel metal2 18998 4284 18998 4284 0 mem_bottom_track_3.DFFR_3_.Q
rlabel metal2 21206 4964 21206 4964 0 mem_bottom_track_3.DFFR_4_.Q
rlabel metal1 32522 3944 32522 3944 0 mem_bottom_track_3.DFFR_5_.Q
rlabel metal2 7958 18802 7958 18802 0 mem_bottom_track_37.DFFR_0_.Q
rlabel metal2 19734 21420 19734 21420 0 mem_bottom_track_37.DFFR_1_.Q
rlabel metal2 13616 17238 13616 17238 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal1 15548 16218 15548 16218 0 mem_bottom_track_5.DFFR_1_.Q
rlabel metal2 7866 8806 7866 8806 0 mem_bottom_track_5.DFFR_2_.Q
rlabel metal1 10120 5542 10120 5542 0 mem_bottom_track_5.DFFR_3_.Q
rlabel metal1 12696 12274 12696 12274 0 mem_bottom_track_5.DFFR_4_.Q
rlabel metal1 17940 10166 17940 10166 0 mem_bottom_track_5.DFFR_5_.Q
rlabel metal1 21344 10166 21344 10166 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal3 10557 14620 10557 14620 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal1 16192 16082 16192 16082 0 mem_bottom_track_7.DFFR_2_.Q
rlabel via3 6555 16660 6555 16660 0 mem_bottom_track_7.DFFR_3_.Q
rlabel metal2 6026 10132 6026 10132 0 mem_bottom_track_7.DFFR_4_.Q
rlabel metal1 5796 16694 5796 16694 0 mem_bottom_track_7.DFFR_5_.Q
rlabel metal1 6670 18700 6670 18700 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal1 20470 18292 20470 18292 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 21068 18734 21068 18734 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 20056 12750 20056 12750 0 mem_left_track_1.DFFR_2_.Q
rlabel metal2 21482 5797 21482 5797 0 mem_left_track_1.DFFR_3_.Q
rlabel metal1 20930 4080 20930 4080 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 18768 5066 18768 5066 0 mem_left_track_1.DFFR_5_.Q
rlabel metal1 15456 8874 15456 8874 0 mem_left_track_17.DFFR_0_.D
rlabel metal2 22218 14773 22218 14773 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 19550 17833 19550 17833 0 mem_left_track_17.DFFR_1_.Q
rlabel metal1 8510 21454 8510 21454 0 mem_left_track_17.DFFR_2_.Q
rlabel metal2 5842 16966 5842 16966 0 mem_left_track_17.DFFR_3_.Q
rlabel metal2 7636 13804 7636 13804 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 10396 14790 10396 14790 0 mem_left_track_17.DFFR_5_.Q
rlabel metal3 11247 16660 11247 16660 0 mem_left_track_17.DFFR_6_.Q
rlabel via3 8211 15300 8211 15300 0 mem_left_track_17.DFFR_7_.Q
rlabel metal1 14076 9078 14076 9078 0 mem_left_track_25.DFFR_0_.Q
rlabel metal2 14858 19244 14858 19244 0 mem_left_track_25.DFFR_1_.Q
rlabel metal1 13984 7990 13984 7990 0 mem_left_track_25.DFFR_2_.Q
rlabel metal2 18308 11594 18308 11594 0 mem_left_track_25.DFFR_3_.Q
rlabel metal1 13938 15470 13938 15470 0 mem_left_track_25.DFFR_4_.Q
rlabel metal1 15078 12410 15078 12410 0 mem_left_track_25.DFFR_5_.Q
rlabel metal1 20654 19754 20654 19754 0 mem_left_track_25.DFFR_6_.Q
rlabel metal1 20930 15062 20930 15062 0 mem_left_track_25.DFFR_7_.Q
rlabel metal1 32384 4114 32384 4114 0 mem_left_track_33.DFFR_0_.Q
rlabel metal2 17710 7344 17710 7344 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 14398 5610 14398 5610 0 mem_left_track_33.DFFR_2_.Q
rlabel metal1 21482 4522 21482 4522 0 mem_left_track_33.DFFR_3_.Q
rlabel metal2 19090 3502 19090 3502 0 mem_left_track_33.DFFR_4_.Q
rlabel metal2 18630 3961 18630 3961 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 18078 6800 18078 6800 0 mem_left_track_9.DFFR_1_.Q
rlabel metal1 21160 18258 21160 18258 0 mem_left_track_9.DFFR_2_.Q
rlabel metal2 2162 9724 2162 9724 0 mem_left_track_9.DFFR_3_.Q
rlabel metal1 14674 3094 14674 3094 0 mem_left_track_9.DFFR_4_.Q
rlabel metal1 15456 2482 15456 2482 0 mem_left_track_9.DFFR_5_.Q
rlabel metal2 16330 1972 16330 1972 0 mem_left_track_9.DFFR_6_.Q
rlabel metal1 21252 2890 21252 2890 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 19734 18632 19734 18632 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 17388 18734 17388 18734 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 21206 8398 21206 8398 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 2346 3128 2346 3128 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 2898 2482 2898 2482 0 mem_right_track_0.DFFR_5_.Q
rlabel metal1 4554 2618 4554 2618 0 mem_right_track_0.DFFR_6_.Q
rlabel metal1 4416 14926 4416 14926 0 mem_right_track_0.DFFR_7_.Q
rlabel metal1 20240 15334 20240 15334 0 mem_right_track_16.DFFR_0_.D
rlabel metal1 21252 10574 21252 10574 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 5934 17714 5934 17714 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 8970 11322 8970 11322 0 mem_right_track_16.DFFR_2_.Q
rlabel metal1 6762 10642 6762 10642 0 mem_right_track_16.DFFR_3_.Q
rlabel metal1 5198 2278 5198 2278 0 mem_right_track_16.DFFR_4_.Q
rlabel metal1 7130 2312 7130 2312 0 mem_right_track_16.DFFR_5_.Q
rlabel metal1 12282 2312 12282 2312 0 mem_right_track_16.DFFR_6_.Q
rlabel metal1 14628 2618 14628 2618 0 mem_right_track_16.DFFR_7_.Q
rlabel metal3 18952 16524 18952 16524 0 mem_right_track_24.DFFR_0_.Q
rlabel via2 13294 16779 13294 16779 0 mem_right_track_24.DFFR_1_.Q
rlabel via2 21850 9027 21850 9027 0 mem_right_track_24.DFFR_2_.Q
rlabel metal2 9982 2074 9982 2074 0 mem_right_track_24.DFFR_3_.Q
rlabel metal1 11546 2550 11546 2550 0 mem_right_track_24.DFFR_4_.Q
rlabel metal1 14904 4182 14904 4182 0 mem_right_track_24.DFFR_5_.Q
rlabel metal1 17250 3910 17250 3910 0 mem_right_track_24.DFFR_6_.Q
rlabel metal2 13294 6137 13294 6137 0 mem_right_track_24.DFFR_7_.Q
rlabel metal1 10442 19380 10442 19380 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 12972 20434 12972 20434 0 mem_right_track_32.DFFR_1_.Q
rlabel metal1 8602 18734 8602 18734 0 mem_right_track_32.DFFR_2_.Q
rlabel metal1 8556 17646 8556 17646 0 mem_right_track_32.DFFR_3_.Q
rlabel via3 14467 16660 14467 16660 0 mem_right_track_32.DFFR_4_.Q
rlabel metal3 7107 14212 7107 14212 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 20233 7174 20233 7174 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 24564 14756 24564 14756 0 mem_right_track_8.DFFR_2_.Q
rlabel metal1 17066 20434 17066 20434 0 mem_right_track_8.DFFR_3_.Q
rlabel metal1 20976 13838 20976 13838 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 19550 6800 19550 6800 0 mem_right_track_8.DFFR_5_.Q
rlabel metal1 21022 5134 21022 5134 0 mem_right_track_8.DFFR_6_.Q
rlabel metal2 19826 16932 19826 16932 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal2 13754 17986 13754 17986 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 16836 18190 16836 18190 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 26266 13192 26266 13192 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal1 19964 17034 19964 17034 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 25944 7786 25944 7786 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 33810 4794 33810 4794 0 mux_bottom_track_1.out
rlabel metal1 19228 16014 19228 16014 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal2 16422 16524 16422 16524 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal2 16790 15810 16790 15810 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 4922 17357 4922 17357 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 2990 8432 2990 8432 0 mux_bottom_track_11.out
rlabel metal1 13064 28390 13064 28390 0 mux_bottom_track_13.INVTX1_0_.out
rlabel metal1 6716 15470 6716 15470 0 mux_bottom_track_13.INVTX1_1_.out
rlabel metal1 6992 15334 6992 15334 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 3542 14076 3542 14076 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 3082 7786 3082 7786 0 mux_bottom_track_13.out
rlabel metal1 20286 15538 20286 15538 0 mux_bottom_track_15.INVTX1_0_.out
rlabel metal1 6210 13770 6210 13770 0 mux_bottom_track_15.INVTX1_1_.out
rlabel metal4 2668 12308 2668 12308 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 2070 9690 2070 9690 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 2070 8330 2070 8330 0 mux_bottom_track_15.out
rlabel metal1 15042 23562 15042 23562 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 12006 19278 12006 19278 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 11132 21658 11132 21658 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12558 21420 12558 21420 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5704 33490 5704 33490 0 mux_bottom_track_17.out
rlabel metal1 16790 24276 16790 24276 0 mux_bottom_track_19.INVTX1_0_.out
rlabel metal2 12742 23358 12742 23358 0 mux_bottom_track_19.INVTX1_2_.out
rlabel metal2 15870 24514 15870 24514 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13800 23562 13800 23562 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14444 32402 14444 32402 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 13938 34102 13938 34102 0 mux_bottom_track_19.out
rlabel metal2 26266 14858 26266 14858 0 mux_bottom_track_21.INVTX1_0_.out
rlabel metal2 34362 4998 34362 4998 0 mux_bottom_track_21.INVTX1_1_.out
rlabel metal2 28474 7548 28474 7548 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 29026 4658 29026 4658 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35558 5644 35558 5644 0 mux_bottom_track_21.out
rlabel metal1 26726 19788 26726 19788 0 mux_bottom_track_23.INVTX1_0_.out
rlabel metal1 19458 18156 19458 18156 0 mux_bottom_track_23.INVTX1_1_.out
rlabel metal1 29670 17102 29670 17102 0 mux_bottom_track_23.INVTX1_2_.out
rlabel metal2 26266 18836 26266 18836 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29164 17034 29164 17034 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 28796 17238 28796 17238 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32154 26350 32154 26350 0 mux_bottom_track_23.out
rlabel metal2 20746 21182 20746 21182 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 20194 19924 20194 19924 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal2 20378 24548 20378 24548 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal1 21114 20774 21114 20774 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 23046 23120 23046 23120 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25208 20842 25208 20842 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 30452 20910 30452 20910 0 mux_bottom_track_25.out
rlabel metal1 18170 25194 18170 25194 0 mux_bottom_track_27.INVTX1_0_.out
rlabel metal2 15548 27132 15548 27132 0 mux_bottom_track_27.INVTX1_1_.out
rlabel metal2 28842 12585 28842 12585 0 mux_bottom_track_27.INVTX1_2_.out
rlabel metal2 20424 20468 20424 20468 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 29394 14178 29394 14178 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 29670 14892 29670 14892 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 29946 7514 29946 7514 0 mux_bottom_track_27.out
rlabel metal1 27600 14314 27600 14314 0 mux_bottom_track_3.INVTX1_0_.out
rlabel metal1 4554 14450 4554 14450 0 mux_bottom_track_3.INVTX1_1_.out
rlabel metal1 23322 7310 23322 7310 0 mux_bottom_track_3.INVTX1_3_.out
rlabel metal1 17986 15538 17986 15538 0 mux_bottom_track_3.INVTX1_4_.out
rlabel metal2 22402 15742 22402 15742 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel via2 12466 12971 12466 12971 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 27738 2890 27738 2890 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 31832 4794 31832 4794 0 mux_bottom_track_3.out
rlabel via3 5267 16524 5267 16524 0 mux_bottom_track_37.INVTX1_1_.out
rlabel metal1 17526 21046 17526 21046 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 25668 22066 25668 22066 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 30314 25466 30314 25466 0 mux_bottom_track_37.out
rlabel metal1 14812 19890 14812 19890 0 mux_bottom_track_5.INVTX1_0_.out
rlabel metal2 12650 21522 12650 21522 0 mux_bottom_track_5.INVTX1_3_.out
rlabel metal1 20056 31994 20056 31994 0 mux_bottom_track_5.INVTX1_4_.out
rlabel metal1 16192 21930 16192 21930 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 15410 18598 15410 18598 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 27554 25874 27554 25874 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 30268 26010 30268 26010 0 mux_bottom_track_5.out
rlabel metal1 19044 21658 19044 21658 0 mux_bottom_track_7.INVTX1_0_.out
rlabel metal1 22954 27846 22954 27846 0 mux_bottom_track_7.INVTX1_2_.out
rlabel metal3 7567 18020 7567 18020 0 mux_bottom_track_7.INVTX1_3_.out
rlabel metal2 11822 15776 11822 15776 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 7406 13906 7406 13906 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 4416 16150 4416 16150 0 mux_bottom_track_7.out
rlabel metal1 12512 17510 12512 17510 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 7084 17102 7084 17102 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 7176 17850 7176 17850 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 7498 19312 7498 19312 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 6440 27098 6440 27098 0 mux_bottom_track_9.out
rlabel metal1 12834 14960 12834 14960 0 mux_left_track_1.INVTX1_3_.out
rlabel metal1 5014 7174 5014 7174 0 mux_left_track_1.INVTX1_4_.out
rlabel metal2 18998 16898 18998 16898 0 mux_left_track_1.INVTX1_5_.out
rlabel via3 15709 16660 15709 16660 0 mux_left_track_1.INVTX1_6_.out
rlabel metal2 29854 28832 29854 28832 0 mux_left_track_1.INVTX1_7_.out
rlabel metal1 21114 16014 21114 16014 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 13478 16728 13478 16728 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 19182 17442 19182 17442 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 34546 9316 34546 9316 0 mux_left_track_1.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 36294 8636 36294 8636 0 mux_left_track_1.out
rlabel metal1 8188 31858 8188 31858 0 mux_left_track_17.INVTX1_3_.out
rlabel metal2 29854 8143 29854 8143 0 mux_left_track_17.INVTX1_4_.out
rlabel metal2 15226 20434 15226 20434 0 mux_left_track_17.INVTX1_5_.out
rlabel metal1 8602 20332 8602 20332 0 mux_left_track_17.INVTX1_6_.out
rlabel metal1 6302 13226 6302 13226 0 mux_left_track_17.INVTX1_7_.out
rlabel metal1 11638 24242 11638 24242 0 mux_left_track_17.INVTX1_8_.out
rlabel metal2 20700 17612 20700 17612 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 16238 19448 16238 19448 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 28474 31892 28474 31892 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 29072 36754 29072 36754 0 mux_left_track_17.out
rlabel metal2 24978 22882 24978 22882 0 mux_left_track_25.INVTX1_3_.out
rlabel metal1 15778 22542 15778 22542 0 mux_left_track_25.INVTX1_4_.out
rlabel metal1 10534 14450 10534 14450 0 mux_left_track_25.INVTX1_5_.out
rlabel metal1 12006 15538 12006 15538 0 mux_left_track_25.INVTX1_6_.out
rlabel metal1 18952 31858 18952 31858 0 mux_left_track_25.INVTX1_7_.out
rlabel metal1 20930 31858 20930 31858 0 mux_left_track_25.INVTX1_8_.out
rlabel metal1 18078 23596 18078 23596 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 11178 22474 11178 22474 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 35282 26928 35282 26928 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 35374 27574 35374 27574 0 mux_left_track_25.out
rlabel metal1 16054 13226 16054 13226 0 mux_left_track_33.INVTX1_2_.out
rlabel metal1 29532 9962 29532 9962 0 mux_left_track_33.INVTX1_3_.out
rlabel metal1 28244 10574 28244 10574 0 mux_left_track_33.INVTX1_4_.out
rlabel metal1 10534 19958 10534 19958 0 mux_left_track_33.INVTX1_5_.out
rlabel metal1 26082 3400 26082 3400 0 mux_left_track_33.INVTX1_6_.out
rlabel metal2 13570 18666 13570 18666 0 mux_left_track_33.INVTX1_7_.out
rlabel metal1 20562 14926 20562 14926 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 17618 12682 17618 12682 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 19826 18836 19826 18836 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 29256 7922 29256 7922 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 33258 11526 33258 11526 0 mux_left_track_33.out
rlabel metal1 26082 18190 26082 18190 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 24794 5746 24794 5746 0 mux_left_track_9.INVTX1_4_.out
rlabel metal2 24426 15844 24426 15844 0 mux_left_track_9.INVTX1_5_.out
rlabel metal2 12098 15300 12098 15300 0 mux_left_track_9.INVTX1_6_.out
rlabel metal1 2254 9486 2254 9486 0 mux_left_track_9.INVTX1_7_.out
rlabel metal2 30682 6341 30682 6341 0 mux_left_track_9.INVTX1_8_.out
rlabel metal1 27232 16150 27232 16150 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 26036 13804 26036 13804 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 36754 22644 36754 22644 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36846 32708 36846 32708 0 mux_left_track_9.out
rlabel metal2 27554 21726 27554 21726 0 mux_right_track_0.INVTX1_0_.out
rlabel metal1 13064 19890 13064 19890 0 mux_right_track_0.INVTX1_1_.out
rlabel metal2 13754 20383 13754 20383 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 16376 14926 16376 14926 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 15410 13192 15410 13192 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 3864 11322 3864 11322 0 mux_right_track_0.out
rlabel metal1 23736 22542 23736 22542 0 mux_right_track_16.INVTX1_0_.out
rlabel metal1 3772 12274 3772 12274 0 mux_right_track_16.INVTX1_1_.out
rlabel metal2 4968 12716 4968 12716 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 8096 20366 8096 20366 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 33672 4046 33672 4046 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 35742 3706 35742 3706 0 mux_right_track_16.out
rlabel metal1 26634 30022 26634 30022 0 mux_right_track_24.INVTX1_0_.out
rlabel metal2 35650 4267 35650 4267 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 26864 17102 26864 17102 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 14214 15946 14214 15946 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 26542 9044 26542 9044 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 33166 4624 33166 4624 0 mux_right_track_24.out
rlabel metal1 7912 17578 7912 17578 0 mux_right_track_32.INVTX1_0_.out
rlabel via2 20562 16643 20562 16643 0 mux_right_track_32.INVTX1_1_.out
rlabel metal1 13524 21590 13524 21590 0 mux_right_track_32.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 14444 17714 14444 17714 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel via1 15134 17306 15134 17306 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 14306 21352 14306 21352 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 25254 23834 25254 23834 0 mux_right_track_32.out
rlabel metal1 22402 2516 22402 2516 0 mux_right_track_8.INVTX1_0_.out
rlabel via2 22402 2941 22402 2941 0 mux_right_track_8.INVTX1_1_.out
rlabel metal1 25254 22508 25254 22508 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 20424 13838 20424 13838 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 36386 26146 36386 26146 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36846 36346 36846 36346 0 mux_right_track_8.out
rlabel metal1 1610 19448 1610 19448 0 net1
rlabel metal2 33074 2635 33074 2635 0 net10
rlabel metal1 18492 23290 18492 23290 0 net100
rlabel metal1 34868 2414 34868 2414 0 net101
rlabel metal1 30130 36890 30130 36890 0 net102
rlabel metal2 34914 36924 34914 36924 0 net103
rlabel metal2 2530 13090 2530 13090 0 net104
rlabel metal2 2714 8415 2714 8415 0 net105
rlabel metal1 1978 29138 1978 29138 0 net106
rlabel metal2 17526 5729 17526 5729 0 net107
rlabel metal2 1610 21692 1610 21692 0 net108
rlabel metal1 18262 5644 18262 5644 0 net109
rlabel metal1 30406 23698 30406 23698 0 net11
rlabel metal2 1610 24582 1610 24582 0 net110
rlabel metal1 32752 37230 32752 37230 0 net111
rlabel metal1 2806 32878 2806 32878 0 net112
rlabel metal1 31050 2380 31050 2380 0 net113
rlabel metal2 38042 24378 38042 24378 0 net114
rlabel metal2 38042 6069 38042 6069 0 net115
rlabel metal2 26358 33422 26358 33422 0 net116
rlabel metal1 37306 36176 37306 36176 0 net117
rlabel metal2 37490 37060 37490 37060 0 net118
rlabel metal2 1610 5916 1610 5916 0 net119
rlabel metal1 24380 37094 24380 37094 0 net12
rlabel via3 17549 19380 17549 19380 0 net120
rlabel metal2 36662 3196 36662 3196 0 net121
rlabel metal1 1610 13940 1610 13940 0 net122
rlabel via2 33626 4709 33626 4709 0 net123
rlabel metal2 38042 5066 38042 5066 0 net124
rlabel metal1 35190 26554 35190 26554 0 net125
rlabel metal1 36961 20910 36961 20910 0 net126
rlabel metal2 32338 4114 32338 4114 0 net127
rlabel metal2 2714 24786 2714 24786 0 net128
rlabel metal2 37858 10438 37858 10438 0 net129
rlabel metal1 4876 32878 4876 32878 0 net13
rlabel metal2 2622 29614 2622 29614 0 net130
rlabel metal1 36961 22610 36961 22610 0 net131
rlabel metal2 33810 32198 33810 32198 0 net132
rlabel metal1 36662 2448 36662 2448 0 net133
rlabel metal1 38042 36108 38042 36108 0 net134
rlabel metal2 1610 12206 1610 12206 0 net135
rlabel metal2 1610 32334 1610 32334 0 net136
rlabel metal2 2346 7310 2346 7310 0 net137
rlabel metal2 2530 6154 2530 6154 0 net138
rlabel metal1 1656 6290 1656 6290 0 net139
rlabel metal1 27830 2006 27830 2006 0 net14
rlabel metal1 3128 36686 3128 36686 0 net140
rlabel metal1 12558 37128 12558 37128 0 net141
rlabel metal1 11408 9554 11408 9554 0 net142
rlabel metal2 22862 16286 22862 16286 0 net143
rlabel metal2 27462 9758 27462 9758 0 net144
rlabel metal1 26864 7922 26864 7922 0 net145
rlabel metal1 27508 12750 27508 12750 0 net146
rlabel metal2 14766 22508 14766 22508 0 net147
rlabel metal1 21574 21658 21574 21658 0 net148
rlabel metal1 13018 22066 13018 22066 0 net149
rlabel metal1 8602 36550 8602 36550 0 net15
rlabel metal2 24242 7616 24242 7616 0 net150
rlabel metal1 3818 15402 3818 15402 0 net151
rlabel metal2 33626 3281 33626 3281 0 net152
rlabel metal1 19642 21454 19642 21454 0 net153
rlabel metal2 9246 19040 9246 19040 0 net154
rlabel metal1 4508 17714 4508 17714 0 net155
rlabel metal2 2806 15436 2806 15436 0 net156
rlabel metal2 2806 10812 2806 10812 0 net157
rlabel metal2 12374 21216 12374 21216 0 net158
rlabel metal1 23368 3570 23368 3570 0 net159
rlabel metal2 26358 3349 26358 3349 0 net16
rlabel metal2 22678 21794 22678 21794 0 net160
rlabel metal2 13846 24208 13846 24208 0 net161
rlabel metal2 28382 18428 28382 18428 0 net162
rlabel metal2 22678 23868 22678 23868 0 net163
rlabel metal2 30038 14688 30038 14688 0 net164
rlabel metal2 24886 17952 24886 17952 0 net165
rlabel metal2 19550 19040 19550 19040 0 net166
rlabel metal2 1886 17374 1886 17374 0 net17
rlabel metal1 4370 6630 4370 6630 0 net18
rlabel metal2 28106 37026 28106 37026 0 net19
rlabel metal1 2484 8058 2484 8058 0 net2
rlabel metal2 2254 6494 2254 6494 0 net20
rlabel metal2 23138 30464 23138 30464 0 net21
rlabel metal1 37766 27302 37766 27302 0 net22
rlabel metal1 7268 18734 7268 18734 0 net23
rlabel metal1 3542 7718 3542 7718 0 net24
rlabel metal1 37766 36550 37766 36550 0 net25
rlabel metal1 20378 37366 20378 37366 0 net26
rlabel metal2 38042 10506 38042 10506 0 net27
rlabel metal1 37536 13906 37536 13906 0 net28
rlabel metal2 38226 16728 38226 16728 0 net29
rlabel metal1 7958 29682 7958 29682 0 net3
rlabel metal1 28382 2482 28382 2482 0 net30
rlabel metal2 20654 33354 20654 33354 0 net31
rlabel metal1 38042 32742 38042 32742 0 net32
rlabel metal2 24886 33762 24886 33762 0 net33
rlabel metal1 13846 32470 13846 32470 0 net34
rlabel metal1 37858 24174 37858 24174 0 net35
rlabel metal1 17894 36788 17894 36788 0 net36
rlabel metal2 11730 34510 11730 34510 0 net37
rlabel metal1 22034 37162 22034 37162 0 net38
rlabel via2 12374 17629 12374 17629 0 net39
rlabel metal2 3174 10438 3174 10438 0 net4
rlabel metal2 16606 37502 16606 37502 0 net40
rlabel metal2 37766 21284 37766 21284 0 net41
rlabel metal2 4278 37060 4278 37060 0 net42
rlabel metal1 37766 2550 37766 2550 0 net43
rlabel metal2 34730 20842 34730 20842 0 net44
rlabel metal2 29026 15674 29026 15674 0 net45
rlabel metal1 16192 36550 16192 36550 0 net46
rlabel metal1 2254 6867 2254 6867 0 net47
rlabel metal1 36984 3978 36984 3978 0 net48
rlabel metal2 38134 16796 38134 16796 0 net49
rlabel metal2 36202 2244 36202 2244 0 net5
rlabel metal2 4094 24990 4094 24990 0 net50
rlabel metal1 4554 36618 4554 36618 0 net51
rlabel metal2 5566 25092 5566 25092 0 net52
rlabel metal2 8326 20468 8326 20468 0 net53
rlabel metal1 4416 36550 4416 36550 0 net54
rlabel metal2 34546 33082 34546 33082 0 net55
rlabel metal1 8372 4794 8372 4794 0 net56
rlabel metal2 6578 17850 6578 17850 0 net57
rlabel metal1 29026 2924 29026 2924 0 net58
rlabel metal2 36754 4930 36754 4930 0 net59
rlabel metal2 1794 22304 1794 22304 0 net6
rlabel metal1 14352 29138 14352 29138 0 net60
rlabel metal1 31556 4250 31556 4250 0 net61
rlabel metal2 3818 8636 3818 8636 0 net62
rlabel metal1 22494 36550 22494 36550 0 net63
rlabel metal2 5658 27132 5658 27132 0 net64
rlabel metal1 4002 3604 4002 3604 0 net65
rlabel metal2 2898 7922 2898 7922 0 net66
rlabel metal1 3680 9146 3680 9146 0 net67
rlabel metal1 21206 37094 21206 37094 0 net68
rlabel metal2 32614 4386 32614 4386 0 net69
rlabel metal2 2530 22559 2530 22559 0 net7
rlabel metal1 34362 36550 34362 36550 0 net70
rlabel metal1 33902 6766 33902 6766 0 net71
rlabel metal1 2162 36006 2162 36006 0 net72
rlabel metal2 2714 12087 2714 12087 0 net73
rlabel metal2 35558 2635 35558 2635 0 net74
rlabel metal2 23874 2822 23874 2822 0 net75
rlabel metal2 38134 24106 38134 24106 0 net76
rlabel metal1 25300 2414 25300 2414 0 net77
rlabel metal1 30130 37094 30130 37094 0 net78
rlabel metal1 28474 37094 28474 37094 0 net79
rlabel metal1 18124 37094 18124 37094 0 net8
rlabel metal1 3680 35462 3680 35462 0 net80
rlabel metal1 9476 37162 9476 37162 0 net81
rlabel metal2 33718 3230 33718 3230 0 net82
rlabel metal1 2208 11866 2208 11866 0 net83
rlabel metal2 29578 3740 29578 3740 0 net84
rlabel metal2 36110 8772 36110 8772 0 net85
rlabel via2 14950 37213 14950 37213 0 net86
rlabel metal2 38042 30396 38042 30396 0 net87
rlabel metal2 36294 28662 36294 28662 0 net88
rlabel metal1 32246 37230 32246 37230 0 net89
rlabel metal2 1886 36555 1886 36555 0 net9
rlabel metal1 21919 3502 21919 3502 0 net90
rlabel metal1 35880 37230 35880 37230 0 net91
rlabel metal2 36938 12342 36938 12342 0 net92
rlabel metal1 33580 2414 33580 2414 0 net93
rlabel metal1 1610 30736 1610 30736 0 net94
rlabel via2 1610 16099 1610 16099 0 net95
rlabel metal1 37996 3502 37996 3502 0 net96
rlabel metal1 18078 36890 18078 36890 0 net97
rlabel metal1 37720 33082 37720 33082 0 net98
rlabel metal2 35926 4657 35926 4657 0 net99
rlabel metal3 1142 10948 1142 10948 0 pReset
rlabel metal1 8280 3706 8280 3706 0 prog_clk
rlabel metal2 13570 1163 13570 1163 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 21298 1146 21298 1146 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal3 38786 25908 38786 25908 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 23276 3910 23276 3910 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 30406 37230 30406 37230 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 29486 37230 29486 37230 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 1242 35666 1242 35666 0 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 7590 37230 7590 37230 0 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 34730 3145 34730 3145 0 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 10268 1234 10268 0 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
