magic
tech sky130A
magscale 1 2
timestamp 1674174325
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 662 39200 718 39800
rect 2594 39200 2650 39800
rect 3882 39200 3938 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9678 39200 9734 39800
rect 10966 39200 11022 39800
rect 12898 39200 12954 39800
rect 14830 39200 14886 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21914 39200 21970 39800
rect 23846 39200 23902 39800
rect 25134 39200 25190 39800
rect 27066 39200 27122 39800
rect 28998 39200 29054 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 34150 39200 34206 39800
rect 36082 39200 36138 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 1306 200 1362 800
rect 3238 200 3294 800
rect 5170 200 5226 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 10322 200 10378 800
rect 12254 200 12310 800
rect 14186 200 14242 800
rect 15474 200 15530 800
rect 17406 200 17462 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 24490 200 24546 800
rect 26422 200 26478 800
rect 28354 200 28410 800
rect 29642 200 29698 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 38658 200 38714 800
<< obsm2 >>
rect 20 39144 606 39250
rect 774 39144 2538 39250
rect 2706 39144 3826 39250
rect 3994 39144 5758 39250
rect 5926 39144 7690 39250
rect 7858 39144 9622 39250
rect 9790 39144 10910 39250
rect 11078 39144 12842 39250
rect 13010 39144 14774 39250
rect 14942 39144 16706 39250
rect 16874 39144 17994 39250
rect 18162 39144 19926 39250
rect 20094 39144 21858 39250
rect 22026 39144 23790 39250
rect 23958 39144 25078 39250
rect 25246 39144 27010 39250
rect 27178 39144 28942 39250
rect 29110 39144 30874 39250
rect 31042 39144 32162 39250
rect 32330 39144 34094 39250
rect 34262 39144 36026 39250
rect 36194 39144 37958 39250
rect 38126 39144 39246 39250
rect 20 856 39356 39144
rect 130 800 1250 856
rect 1418 800 3182 856
rect 3350 800 5114 856
rect 5282 800 7046 856
rect 7214 800 8334 856
rect 8502 800 10266 856
rect 10434 800 12198 856
rect 12366 800 14130 856
rect 14298 800 15418 856
rect 15586 800 17350 856
rect 17518 800 19282 856
rect 19450 800 21214 856
rect 21382 800 22502 856
rect 22670 800 24434 856
rect 24602 800 26366 856
rect 26534 800 28298 856
rect 28466 800 29586 856
rect 29754 800 31518 856
rect 31686 800 33450 856
rect 33618 800 35382 856
rect 35550 800 36670 856
rect 36838 800 38602 856
rect 38770 800 39356 856
<< metal3 >>
rect 200 38768 800 38888
rect 39200 38088 39800 38208
rect 200 36728 800 36848
rect 39200 36048 39800 36168
rect 200 35368 800 35488
rect 39200 34008 39800 34128
rect 200 33328 800 33448
rect 39200 32648 39800 32768
rect 200 31288 800 31408
rect 39200 30608 39800 30728
rect 200 29248 800 29368
rect 39200 28568 39800 28688
rect 200 27888 800 28008
rect 39200 26528 39800 26648
rect 200 25848 800 25968
rect 39200 25168 39800 25288
rect 200 23808 800 23928
rect 39200 23128 39800 23248
rect 200 21768 800 21888
rect 39200 21088 39800 21208
rect 200 20408 800 20528
rect 39200 19048 39800 19168
rect 200 18368 800 18488
rect 39200 17688 39800 17808
rect 200 16328 800 16448
rect 39200 15648 39800 15768
rect 200 14288 800 14408
rect 39200 13608 39800 13728
rect 200 12928 800 13048
rect 39200 11568 39800 11688
rect 200 10888 800 11008
rect 39200 10208 39800 10328
rect 200 8848 800 8968
rect 39200 8168 39800 8288
rect 200 6808 800 6928
rect 39200 6128 39800 6248
rect 200 5448 800 5568
rect 39200 4088 39800 4208
rect 200 3408 800 3528
rect 39200 2728 39800 2848
rect 200 1368 800 1488
rect 39200 688 39800 808
<< obsm3 >>
rect 880 38688 39314 38861
rect 800 38288 39314 38688
rect 800 38008 39120 38288
rect 800 36928 39314 38008
rect 880 36648 39314 36928
rect 800 36248 39314 36648
rect 800 35968 39120 36248
rect 800 35568 39314 35968
rect 880 35288 39314 35568
rect 800 34208 39314 35288
rect 800 33928 39120 34208
rect 800 33528 39314 33928
rect 880 33248 39314 33528
rect 800 32848 39314 33248
rect 800 32568 39120 32848
rect 800 31488 39314 32568
rect 880 31208 39314 31488
rect 800 30808 39314 31208
rect 800 30528 39120 30808
rect 800 29448 39314 30528
rect 880 29168 39314 29448
rect 800 28768 39314 29168
rect 800 28488 39120 28768
rect 800 28088 39314 28488
rect 880 27808 39314 28088
rect 800 26728 39314 27808
rect 800 26448 39120 26728
rect 800 26048 39314 26448
rect 880 25768 39314 26048
rect 800 25368 39314 25768
rect 800 25088 39120 25368
rect 800 24008 39314 25088
rect 880 23728 39314 24008
rect 800 23328 39314 23728
rect 800 23048 39120 23328
rect 800 21968 39314 23048
rect 880 21688 39314 21968
rect 800 21288 39314 21688
rect 800 21008 39120 21288
rect 800 20608 39314 21008
rect 880 20328 39314 20608
rect 800 19248 39314 20328
rect 800 18968 39120 19248
rect 800 18568 39314 18968
rect 880 18288 39314 18568
rect 800 17888 39314 18288
rect 800 17608 39120 17888
rect 800 16528 39314 17608
rect 880 16248 39314 16528
rect 800 15848 39314 16248
rect 800 15568 39120 15848
rect 800 14488 39314 15568
rect 880 14208 39314 14488
rect 800 13808 39314 14208
rect 800 13528 39120 13808
rect 800 13128 39314 13528
rect 880 12848 39314 13128
rect 800 11768 39314 12848
rect 800 11488 39120 11768
rect 800 11088 39314 11488
rect 880 10808 39314 11088
rect 800 10408 39314 10808
rect 800 10128 39120 10408
rect 800 9048 39314 10128
rect 880 8768 39314 9048
rect 800 8368 39314 8768
rect 800 8088 39120 8368
rect 800 7008 39314 8088
rect 880 6728 39314 7008
rect 800 6328 39314 6728
rect 800 6048 39120 6328
rect 800 5648 39314 6048
rect 880 5368 39314 5648
rect 800 4288 39314 5368
rect 800 4008 39120 4288
rect 800 3608 39314 4008
rect 880 3328 39314 3608
rect 800 2928 39314 3328
rect 800 2648 39120 2928
rect 800 1568 39314 2648
rect 880 1288 39314 1568
rect 800 888 39314 1288
rect 800 718 39120 888
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal2 s 8390 200 8446 800 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 200 25848 800 25968 6 ccff_tail
port 2 nsew signal output
rlabel metal3 s 200 31288 800 31408 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 18050 39200 18106 39800 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal2 s 5814 39200 5870 39800 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal3 s 39200 6128 39800 6248 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal3 s 39200 32648 39800 32768 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal3 s 39200 8168 39800 8288 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 28354 200 28410 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal3 s 39200 36048 39800 36168 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal3 s 200 36728 800 36848 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal2 s 14186 200 14242 800 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal3 s 39200 28568 39800 28688 6 chany_bottom_in[1]
port 13 nsew signal input
rlabel metal3 s 39200 688 39800 808 6 chany_bottom_in[2]
port 14 nsew signal input
rlabel metal3 s 39200 25168 39800 25288 6 chany_bottom_in[3]
port 15 nsew signal input
rlabel metal3 s 200 14288 800 14408 6 chany_bottom_in[4]
port 16 nsew signal input
rlabel metal2 s 38014 39200 38070 39800 6 chany_bottom_in[5]
port 17 nsew signal input
rlabel metal3 s 39200 13608 39800 13728 6 chany_bottom_in[6]
port 18 nsew signal input
rlabel metal2 s 16762 39200 16818 39800 6 chany_bottom_in[7]
port 19 nsew signal input
rlabel metal2 s 36726 200 36782 800 6 chany_bottom_in[8]
port 20 nsew signal input
rlabel metal2 s 33506 200 33562 800 6 chany_bottom_in[9]
port 21 nsew signal input
rlabel metal2 s 35438 200 35494 800 6 chany_bottom_out[0]
port 22 nsew signal output
rlabel metal2 s 25134 39200 25190 39800 6 chany_bottom_out[10]
port 23 nsew signal output
rlabel metal3 s 39200 26528 39800 26648 6 chany_bottom_out[11]
port 24 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 chany_bottom_out[12]
port 25 nsew signal output
rlabel metal3 s 200 23808 800 23928 6 chany_bottom_out[13]
port 26 nsew signal output
rlabel metal3 s 39200 15648 39800 15768 6 chany_bottom_out[14]
port 27 nsew signal output
rlabel metal2 s 21914 39200 21970 39800 6 chany_bottom_out[15]
port 28 nsew signal output
rlabel metal3 s 200 29248 800 29368 6 chany_bottom_out[16]
port 29 nsew signal output
rlabel metal2 s 28998 39200 29054 39800 6 chany_bottom_out[17]
port 30 nsew signal output
rlabel metal3 s 200 3408 800 3528 6 chany_bottom_out[18]
port 31 nsew signal output
rlabel metal3 s 39200 30608 39800 30728 6 chany_bottom_out[1]
port 32 nsew signal output
rlabel metal3 s 200 1368 800 1488 6 chany_bottom_out[2]
port 33 nsew signal output
rlabel metal2 s 19982 39200 20038 39800 6 chany_bottom_out[3]
port 34 nsew signal output
rlabel metal3 s 200 8848 800 8968 6 chany_bottom_out[4]
port 35 nsew signal output
rlabel metal3 s 200 21768 800 21888 6 chany_bottom_out[5]
port 36 nsew signal output
rlabel metal2 s 27066 39200 27122 39800 6 chany_bottom_out[6]
port 37 nsew signal output
rlabel metal2 s 34150 39200 34206 39800 6 chany_bottom_out[7]
port 38 nsew signal output
rlabel metal2 s 662 39200 718 39800 6 chany_bottom_out[8]
port 39 nsew signal output
rlabel metal2 s 2594 39200 2650 39800 6 chany_bottom_out[9]
port 40 nsew signal output
rlabel metal2 s 15474 200 15530 800 6 chany_top_in[0]
port 41 nsew signal input
rlabel metal3 s 200 6808 800 6928 6 chany_top_in[10]
port 42 nsew signal input
rlabel metal3 s 39200 34008 39800 34128 6 chany_top_in[11]
port 43 nsew signal input
rlabel metal3 s 200 20408 800 20528 6 chany_top_in[12]
port 44 nsew signal input
rlabel metal2 s 3238 200 3294 800 6 chany_top_in[13]
port 45 nsew signal input
rlabel metal2 s 10322 200 10378 800 6 chany_top_in[14]
port 46 nsew signal input
rlabel metal2 s 31574 200 31630 800 6 chany_top_in[15]
port 47 nsew signal input
rlabel metal3 s 39200 11568 39800 11688 6 chany_top_in[16]
port 48 nsew signal input
rlabel metal3 s 39200 4088 39800 4208 6 chany_top_in[17]
port 49 nsew signal input
rlabel metal2 s 24490 200 24546 800 6 chany_top_in[18]
port 50 nsew signal input
rlabel metal3 s 200 38768 800 38888 6 chany_top_in[1]
port 51 nsew signal input
rlabel metal2 s 38658 200 38714 800 6 chany_top_in[2]
port 52 nsew signal input
rlabel metal2 s 10966 39200 11022 39800 6 chany_top_in[3]
port 53 nsew signal input
rlabel metal3 s 39200 10208 39800 10328 6 chany_top_in[4]
port 54 nsew signal input
rlabel metal3 s 39200 19048 39800 19168 6 chany_top_in[5]
port 55 nsew signal input
rlabel metal2 s 29642 200 29698 800 6 chany_top_in[6]
port 56 nsew signal input
rlabel metal3 s 200 18368 800 18488 6 chany_top_in[7]
port 57 nsew signal input
rlabel metal2 s 7746 39200 7802 39800 6 chany_top_in[8]
port 58 nsew signal input
rlabel metal2 s 14830 39200 14886 39800 6 chany_top_in[9]
port 59 nsew signal input
rlabel metal3 s 200 33328 800 33448 6 chany_top_out[0]
port 60 nsew signal output
rlabel metal2 s 18 200 74 800 6 chany_top_out[10]
port 61 nsew signal output
rlabel metal2 s 22558 200 22614 800 6 chany_top_out[11]
port 62 nsew signal output
rlabel metal2 s 12898 39200 12954 39800 6 chany_top_out[12]
port 63 nsew signal output
rlabel metal2 s 23846 39200 23902 39800 6 chany_top_out[13]
port 64 nsew signal output
rlabel metal2 s 36082 39200 36138 39800 6 chany_top_out[14]
port 65 nsew signal output
rlabel metal3 s 200 27888 800 28008 6 chany_top_out[15]
port 66 nsew signal output
rlabel metal2 s 5170 200 5226 800 6 chany_top_out[16]
port 67 nsew signal output
rlabel metal2 s 1306 200 1362 800 6 chany_top_out[17]
port 68 nsew signal output
rlabel metal2 s 39302 39200 39358 39800 6 chany_top_out[18]
port 69 nsew signal output
rlabel metal3 s 200 5448 800 5568 6 chany_top_out[1]
port 70 nsew signal output
rlabel metal2 s 17406 200 17462 800 6 chany_top_out[2]
port 71 nsew signal output
rlabel metal3 s 39200 38088 39800 38208 6 chany_top_out[3]
port 72 nsew signal output
rlabel metal3 s 39200 2728 39800 2848 6 chany_top_out[4]
port 73 nsew signal output
rlabel metal3 s 200 10888 800 11008 6 chany_top_out[5]
port 74 nsew signal output
rlabel metal3 s 39200 21088 39800 21208 6 chany_top_out[6]
port 75 nsew signal output
rlabel metal2 s 7102 200 7158 800 6 chany_top_out[7]
port 76 nsew signal output
rlabel metal2 s 12254 200 12310 800 6 chany_top_out[8]
port 77 nsew signal output
rlabel metal3 s 200 16328 800 16448 6 chany_top_out[9]
port 78 nsew signal output
rlabel metal3 s 39200 23128 39800 23248 6 left_grid_right_width_0_height_0_subtile_0__pin_I_1_
port 79 nsew signal output
rlabel metal2 s 21270 200 21326 800 6 left_grid_right_width_0_height_0_subtile_0__pin_I_5_
port 80 nsew signal output
rlabel metal2 s 32218 39200 32274 39800 6 left_grid_right_width_0_height_0_subtile_0__pin_I_9_
port 81 nsew signal output
rlabel metal2 s 30930 39200 30986 39800 6 pReset
port 82 nsew signal input
rlabel metal2 s 3882 39200 3938 39800 6 prog_clk
port 83 nsew signal input
rlabel metal2 s 9678 39200 9734 39800 6 right_grid_left_width_0_height_0_subtile_0__pin_I_11_
port 84 nsew signal output
rlabel metal2 s 26422 200 26478 800 6 right_grid_left_width_0_height_0_subtile_0__pin_I_3_
port 85 nsew signal output
rlabel metal3 s 200 12928 800 13048 6 right_grid_left_width_0_height_0_subtile_0__pin_I_7_
port 86 nsew signal output
rlabel metal3 s 200 35368 800 35488 6 vccd1
port 87 nsew signal bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 87 nsew signal bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 87 nsew signal bidirectional
rlabel metal3 s 39200 17688 39800 17808 6 vssd1
port 88 nsew signal bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 88 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1295302
string GDS_FILE /home/baungarten/Proyectos_caravel/FPGA_3/openlane/cby_1__1_/runs/23_01_19_18_25/results/signoff/cby_1__1_.magic.gds
string GDS_START 134360
<< end >>

