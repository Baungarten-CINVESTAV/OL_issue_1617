magic
tech sky130A
magscale 1 2
timestamp 1674175616
<< viali >>
rect 1593 37213 1627 37247
rect 2513 37213 2547 37247
rect 3157 37213 3191 37247
rect 4169 37213 4203 37247
rect 4813 37213 4847 37247
rect 6561 37213 6595 37247
rect 7849 37213 7883 37247
rect 9321 37213 9355 37247
rect 10425 37213 10459 37247
rect 12357 37213 12391 37247
rect 14473 37213 14507 37247
rect 15577 37213 15611 37247
rect 16865 37213 16899 37247
rect 18337 37213 18371 37247
rect 20085 37213 20119 37247
rect 22017 37213 22051 37247
rect 22937 37213 22971 37247
rect 24777 37213 24811 37247
rect 26065 37213 26099 37247
rect 27813 37213 27847 37247
rect 29745 37213 29779 37247
rect 30665 37213 30699 37247
rect 32505 37213 32539 37247
rect 33793 37213 33827 37247
rect 34897 37213 34931 37247
rect 36921 37213 36955 37247
rect 37473 37213 37507 37247
rect 1777 37077 1811 37111
rect 2329 37077 2363 37111
rect 2973 37077 3007 37111
rect 3985 37077 4019 37111
rect 4629 37077 4663 37111
rect 6745 37077 6779 37111
rect 8033 37077 8067 37111
rect 9137 37077 9171 37111
rect 10609 37077 10643 37111
rect 12541 37077 12575 37111
rect 14289 37077 14323 37111
rect 15761 37077 15795 37111
rect 17049 37077 17083 37111
rect 18153 37077 18187 37111
rect 20269 37077 20303 37111
rect 22201 37077 22235 37111
rect 22753 37077 22787 37111
rect 24593 37077 24627 37111
rect 25881 37077 25915 37111
rect 27997 37077 28031 37111
rect 29929 37077 29963 37111
rect 30481 37077 30515 37111
rect 32321 37077 32355 37111
rect 33609 37077 33643 37111
rect 35081 37077 35115 37111
rect 36737 37077 36771 37111
rect 37657 37077 37691 37111
rect 1777 36873 1811 36907
rect 3525 36873 3559 36907
rect 25329 36873 25363 36907
rect 31493 36873 31527 36907
rect 36001 36873 36035 36907
rect 38209 36873 38243 36907
rect 1593 36737 1627 36771
rect 3709 36737 3743 36771
rect 4905 36737 4939 36771
rect 25513 36737 25547 36771
rect 31677 36737 31711 36771
rect 33149 36737 33183 36771
rect 36185 36737 36219 36771
rect 36921 36737 36955 36771
rect 38025 36737 38059 36771
rect 4721 36601 4755 36635
rect 32965 36601 32999 36635
rect 36737 36533 36771 36567
rect 3985 36329 4019 36363
rect 11621 36329 11655 36363
rect 29837 36329 29871 36363
rect 34989 36329 35023 36363
rect 4077 36125 4111 36159
rect 11805 36125 11839 36159
rect 29745 36125 29779 36159
rect 34897 36125 34931 36159
rect 38301 36125 38335 36159
rect 38117 35989 38151 36023
rect 24501 35785 24535 35819
rect 24409 35649 24443 35683
rect 8309 35241 8343 35275
rect 15485 35241 15519 35275
rect 8217 35037 8251 35071
rect 15669 35037 15703 35071
rect 38025 35037 38059 35071
rect 38209 34901 38243 34935
rect 5549 34697 5583 34731
rect 6837 34697 6871 34731
rect 14657 34697 14691 34731
rect 15301 34697 15335 34731
rect 17693 34697 17727 34731
rect 18797 34697 18831 34731
rect 27445 34697 27479 34731
rect 5733 34561 5767 34595
rect 7021 34561 7055 34595
rect 14841 34561 14875 34595
rect 15485 34561 15519 34595
rect 17877 34561 17911 34595
rect 18981 34561 19015 34595
rect 27629 34561 27663 34595
rect 15853 34085 15887 34119
rect 9137 33949 9171 33983
rect 14289 33949 14323 33983
rect 15761 33949 15795 33983
rect 23029 33949 23063 33983
rect 25053 33949 25087 33983
rect 27997 33949 28031 33983
rect 9229 33813 9263 33847
rect 14381 33813 14415 33847
rect 23121 33813 23155 33847
rect 25145 33813 25179 33847
rect 28089 33813 28123 33847
rect 1777 33473 1811 33507
rect 38301 33473 38335 33507
rect 1593 33269 1627 33303
rect 38117 33269 38151 33303
rect 27629 33065 27663 33099
rect 5641 32861 5675 32895
rect 27537 32861 27571 32895
rect 5733 32725 5767 32759
rect 1777 32385 1811 32419
rect 38025 32385 38059 32419
rect 1593 32181 1627 32215
rect 38209 32181 38243 32215
rect 6561 31977 6595 32011
rect 12173 31977 12207 32011
rect 21005 31841 21039 31875
rect 6469 31773 6503 31807
rect 12081 31773 12115 31807
rect 20913 31773 20947 31807
rect 33609 31773 33643 31807
rect 33701 31773 33735 31807
rect 10241 31297 10275 31331
rect 13829 31297 13863 31331
rect 27169 31297 27203 31331
rect 10333 31093 10367 31127
rect 13921 31093 13955 31127
rect 27261 31093 27295 31127
rect 34897 30889 34931 30923
rect 1777 30685 1811 30719
rect 24869 30685 24903 30719
rect 29745 30685 29779 30719
rect 35081 30685 35115 30719
rect 1593 30549 1627 30583
rect 24961 30549 24995 30583
rect 29837 30549 29871 30583
rect 8861 30209 8895 30243
rect 29929 30209 29963 30243
rect 38025 30209 38059 30243
rect 8953 30005 8987 30039
rect 30021 30005 30055 30039
rect 38209 30005 38243 30039
rect 14841 29801 14875 29835
rect 16957 29801 16991 29835
rect 34989 29801 35023 29835
rect 6193 29597 6227 29631
rect 14749 29597 14783 29631
rect 16865 29597 16899 29631
rect 35173 29597 35207 29631
rect 6285 29461 6319 29495
rect 14197 29257 14231 29291
rect 17509 29257 17543 29291
rect 27261 29257 27295 29291
rect 1777 29121 1811 29155
rect 14105 29121 14139 29155
rect 17417 29121 17451 29155
rect 27169 29121 27203 29155
rect 38301 29121 38335 29155
rect 1593 28985 1627 29019
rect 38117 28985 38151 29019
rect 5641 28713 5675 28747
rect 17141 28713 17175 28747
rect 32873 28713 32907 28747
rect 5549 28509 5583 28543
rect 17049 28509 17083 28543
rect 32781 28509 32815 28543
rect 4261 28033 4295 28067
rect 30389 28033 30423 28067
rect 4353 27829 4387 27863
rect 30481 27829 30515 27863
rect 1777 27421 1811 27455
rect 21005 27421 21039 27455
rect 38025 27421 38059 27455
rect 1593 27285 1627 27319
rect 20821 27285 20855 27319
rect 38209 27285 38243 27319
rect 29193 27081 29227 27115
rect 6561 26945 6595 26979
rect 20913 26945 20947 26979
rect 29101 26945 29135 26979
rect 6653 26741 6687 26775
rect 20729 26741 20763 26775
rect 12725 26469 12759 26503
rect 13369 26469 13403 26503
rect 15945 26469 15979 26503
rect 12265 26333 12299 26367
rect 12909 26333 12943 26367
rect 13553 26333 13587 26367
rect 16129 26333 16163 26367
rect 17233 26333 17267 26367
rect 21005 26333 21039 26367
rect 21097 26265 21131 26299
rect 12081 26197 12115 26231
rect 17049 26197 17083 26231
rect 33609 25993 33643 26027
rect 36737 25993 36771 26027
rect 10609 25857 10643 25891
rect 11989 25857 12023 25891
rect 12633 25857 12667 25891
rect 14197 25857 14231 25891
rect 15301 25857 15335 25891
rect 16865 25857 16899 25891
rect 17693 25857 17727 25891
rect 23581 25857 23615 25891
rect 33793 25857 33827 25891
rect 36921 25857 36955 25891
rect 13553 25789 13587 25823
rect 15945 25789 15979 25823
rect 10701 25653 10735 25687
rect 11805 25653 11839 25687
rect 12449 25653 12483 25687
rect 14289 25653 14323 25687
rect 15393 25653 15427 25687
rect 16957 25653 16991 25687
rect 17509 25653 17543 25687
rect 23397 25653 23431 25687
rect 9781 25449 9815 25483
rect 14749 25449 14783 25483
rect 1593 25381 1627 25415
rect 11069 25381 11103 25415
rect 10425 25313 10459 25347
rect 10609 25313 10643 25347
rect 12725 25313 12759 25347
rect 14289 25313 14323 25347
rect 14473 25313 14507 25347
rect 15945 25313 15979 25347
rect 16129 25313 16163 25347
rect 1777 25245 1811 25279
rect 5181 25245 5215 25279
rect 9965 25245 9999 25279
rect 12541 25245 12575 25279
rect 17233 25245 17267 25279
rect 23581 25245 23615 25279
rect 38301 25245 38335 25279
rect 4997 25109 5031 25143
rect 13185 25109 13219 25143
rect 16589 25109 16623 25143
rect 17049 25109 17083 25143
rect 20361 25109 20395 25143
rect 23397 25109 23431 25143
rect 38117 25109 38151 25143
rect 14381 24905 14415 24939
rect 15209 24837 15243 24871
rect 17049 24837 17083 24871
rect 5181 24769 5215 24803
rect 7297 24769 7331 24803
rect 8861 24769 8895 24803
rect 9965 24769 9999 24803
rect 11989 24769 12023 24803
rect 12633 24769 12667 24803
rect 13277 24769 13311 24803
rect 13921 24769 13955 24803
rect 20361 24769 20395 24803
rect 20545 24769 20579 24803
rect 22201 24769 22235 24803
rect 23305 24769 23339 24803
rect 33333 24769 33367 24803
rect 35541 24769 35575 24803
rect 35633 24769 35667 24803
rect 9045 24701 9079 24735
rect 10057 24701 10091 24735
rect 13737 24701 13771 24735
rect 15117 24701 15151 24735
rect 16957 24701 16991 24735
rect 22661 24701 22695 24735
rect 9505 24633 9539 24667
rect 12449 24633 12483 24667
rect 15669 24633 15703 24667
rect 17509 24633 17543 24667
rect 4997 24565 5031 24599
rect 7113 24565 7147 24599
rect 11805 24565 11839 24599
rect 13093 24565 13127 24599
rect 20821 24565 20855 24599
rect 22017 24565 22051 24599
rect 23397 24565 23431 24599
rect 33425 24565 33459 24599
rect 15209 24361 15243 24395
rect 16589 24361 16623 24395
rect 20821 24361 20855 24395
rect 21925 24293 21959 24327
rect 15025 24225 15059 24259
rect 16221 24225 16255 24259
rect 16405 24225 16439 24259
rect 20177 24225 20211 24259
rect 20361 24225 20395 24259
rect 21373 24225 21407 24259
rect 22753 24225 22787 24259
rect 1593 24157 1627 24191
rect 2329 24157 2363 24191
rect 4169 24157 4203 24191
rect 7573 24157 7607 24191
rect 11621 24157 11655 24191
rect 12449 24157 12483 24191
rect 12909 24157 12943 24191
rect 13737 24157 13771 24191
rect 14841 24157 14875 24191
rect 22569 24157 22603 24191
rect 24777 24157 24811 24191
rect 38301 24157 38335 24191
rect 21465 24089 21499 24123
rect 1777 24021 1811 24055
rect 2421 24021 2455 24055
rect 3985 24021 4019 24055
rect 6745 24021 6779 24055
rect 7389 24021 7423 24055
rect 11713 24021 11747 24055
rect 12265 24021 12299 24055
rect 13001 24021 13035 24055
rect 13553 24021 13587 24055
rect 23213 24021 23247 24055
rect 24593 24021 24627 24055
rect 38117 24021 38151 24055
rect 1777 23817 1811 23851
rect 10333 23817 10367 23851
rect 12541 23817 12575 23851
rect 13185 23817 13219 23851
rect 14473 23817 14507 23851
rect 20361 23817 20395 23851
rect 22017 23817 22051 23851
rect 23305 23817 23339 23851
rect 15301 23749 15335 23783
rect 15853 23749 15887 23783
rect 1961 23681 1995 23715
rect 2513 23681 2547 23715
rect 3157 23681 3191 23715
rect 3893 23681 3927 23715
rect 4537 23681 4571 23715
rect 5365 23681 5399 23715
rect 7021 23681 7055 23715
rect 7665 23681 7699 23715
rect 9413 23681 9447 23715
rect 10517 23681 10551 23715
rect 11161 23681 11195 23715
rect 12725 23681 12759 23715
rect 13369 23681 13403 23715
rect 13829 23681 13863 23715
rect 14657 23681 14691 23715
rect 17601 23681 17635 23715
rect 18429 23681 18463 23715
rect 19257 23681 19291 23715
rect 20545 23681 20579 23715
rect 21189 23681 21223 23715
rect 22201 23681 22235 23715
rect 22661 23681 22695 23715
rect 22845 23681 22879 23715
rect 23949 23681 23983 23715
rect 25237 23681 25271 23715
rect 11897 23613 11931 23647
rect 15209 23613 15243 23647
rect 16865 23613 16899 23647
rect 24409 23613 24443 23647
rect 3985 23545 4019 23579
rect 7113 23545 7147 23579
rect 2605 23477 2639 23511
rect 3249 23477 3283 23511
rect 4629 23477 4663 23511
rect 5181 23477 5215 23511
rect 7757 23477 7791 23511
rect 9229 23477 9263 23511
rect 10977 23477 11011 23511
rect 13921 23477 13955 23511
rect 17693 23477 17727 23511
rect 18521 23477 18555 23511
rect 19073 23477 19107 23511
rect 21005 23477 21039 23511
rect 23765 23477 23799 23511
rect 25053 23477 25087 23511
rect 8401 23273 8435 23307
rect 20085 23273 20119 23307
rect 1593 23205 1627 23239
rect 4077 23205 4111 23239
rect 12541 23205 12575 23239
rect 14657 23205 14691 23239
rect 17785 23205 17819 23239
rect 4905 23137 4939 23171
rect 5089 23137 5123 23171
rect 6745 23137 6779 23171
rect 7389 23137 7423 23171
rect 9689 23137 9723 23171
rect 11897 23137 11931 23171
rect 12081 23137 12115 23171
rect 13093 23137 13127 23171
rect 13737 23137 13771 23171
rect 14473 23137 14507 23171
rect 17141 23137 17175 23171
rect 17325 23137 17359 23171
rect 18429 23137 18463 23171
rect 21005 23137 21039 23171
rect 22385 23137 22419 23171
rect 24593 23137 24627 23171
rect 24777 23137 24811 23171
rect 1777 23069 1811 23103
rect 2605 23069 2639 23103
rect 3157 23069 3191 23103
rect 3985 23069 4019 23103
rect 6009 23069 6043 23103
rect 8585 23069 8619 23103
rect 9505 23069 9539 23103
rect 11253 23069 11287 23103
rect 14289 23069 14323 23103
rect 15393 23069 15427 23103
rect 16221 23069 16255 23103
rect 18245 23069 18279 23103
rect 19625 23069 19659 23103
rect 20269 23069 20303 23103
rect 20821 23069 20855 23103
rect 24041 23069 24075 23103
rect 33977 23069 34011 23103
rect 5549 23001 5583 23035
rect 6837 23001 6871 23035
rect 13185 23001 13219 23035
rect 21465 23001 21499 23035
rect 22477 23001 22511 23035
rect 23397 23001 23431 23035
rect 2421 22933 2455 22967
rect 3249 22933 3283 22967
rect 6101 22933 6135 22967
rect 10149 22933 10183 22967
rect 10609 22933 10643 22967
rect 11345 22933 11379 22967
rect 15485 22933 15519 22967
rect 16037 22933 16071 22967
rect 18889 22933 18923 22967
rect 19441 22933 19475 22967
rect 23857 22933 23891 22967
rect 25237 22933 25271 22967
rect 34069 22933 34103 22967
rect 1593 22729 1627 22763
rect 9413 22729 9447 22763
rect 18613 22729 18647 22763
rect 20177 22729 20211 22763
rect 25053 22729 25087 22763
rect 25513 22729 25547 22763
rect 12173 22661 12207 22695
rect 12265 22661 12299 22695
rect 12817 22661 12851 22695
rect 15117 22661 15151 22695
rect 15669 22661 15703 22695
rect 21373 22661 21407 22695
rect 22201 22661 22235 22695
rect 23305 22661 23339 22695
rect 23397 22661 23431 22695
rect 1777 22593 1811 22627
rect 4905 22593 4939 22627
rect 5549 22593 5583 22627
rect 6561 22593 6595 22627
rect 7297 22593 7331 22627
rect 8493 22593 8527 22627
rect 10057 22593 10091 22627
rect 13829 22593 13863 22627
rect 16129 22593 16163 22627
rect 17049 22593 17083 22627
rect 17969 22593 18003 22627
rect 18153 22593 18187 22627
rect 19257 22593 19291 22627
rect 20361 22593 20395 22627
rect 21281 22593 21315 22627
rect 25697 22593 25731 22627
rect 32321 22593 32355 22627
rect 2605 22525 2639 22559
rect 2881 22525 2915 22559
rect 10241 22525 10275 22559
rect 14013 22525 14047 22559
rect 15025 22525 15059 22559
rect 19073 22525 19107 22559
rect 22109 22525 22143 22559
rect 24409 22525 24443 22559
rect 24593 22525 24627 22559
rect 7389 22457 7423 22491
rect 22661 22457 22695 22491
rect 23857 22457 23891 22491
rect 4353 22389 4387 22423
rect 4997 22389 5031 22423
rect 5641 22389 5675 22423
rect 6653 22389 6687 22423
rect 8309 22389 8343 22423
rect 10701 22389 10735 22423
rect 14197 22389 14231 22423
rect 16221 22389 16255 22423
rect 16865 22389 16899 22423
rect 19441 22389 19475 22423
rect 32413 22389 32447 22423
rect 1948 22185 1982 22219
rect 4077 22185 4111 22219
rect 8217 22185 8251 22219
rect 9689 22185 9723 22219
rect 10596 22185 10630 22219
rect 12081 22117 12115 22151
rect 24961 22117 24995 22151
rect 4169 22049 4203 22083
rect 5917 22049 5951 22083
rect 8033 22049 8067 22083
rect 12726 22049 12760 22083
rect 18705 22049 18739 22083
rect 19441 22049 19475 22083
rect 19625 22049 19659 22083
rect 24777 22049 24811 22083
rect 26433 22049 26467 22083
rect 1685 21981 1719 22015
rect 6377 21981 6411 22015
rect 7205 21981 7239 22015
rect 7849 21981 7883 22015
rect 9873 21981 9907 22015
rect 10333 21981 10367 22015
rect 12541 21981 12575 22015
rect 15393 21981 15427 22015
rect 16037 21981 16071 22015
rect 16497 21981 16531 22015
rect 20729 21981 20763 22015
rect 21189 21981 21223 22015
rect 22109 21981 22143 22015
rect 22845 21981 22879 22015
rect 23029 21981 23063 22015
rect 24593 21981 24627 22015
rect 26341 21981 26375 22015
rect 31677 21981 31711 22015
rect 38301 21981 38335 22015
rect 4445 21913 4479 21947
rect 14749 21913 14783 21947
rect 14841 21913 14875 21947
rect 17601 21913 17635 21947
rect 17693 21913 17727 21947
rect 18245 21913 18279 21947
rect 25697 21913 25731 21947
rect 31861 21913 31895 21947
rect 3433 21845 3467 21879
rect 6193 21845 6227 21879
rect 7297 21845 7331 21879
rect 13185 21845 13219 21879
rect 15853 21845 15887 21879
rect 16589 21845 16623 21879
rect 20085 21845 20119 21879
rect 20545 21845 20579 21879
rect 21281 21845 21315 21879
rect 21925 21845 21959 21879
rect 23489 21845 23523 21879
rect 38117 21845 38151 21879
rect 6561 21641 6595 21675
rect 12081 21641 12115 21675
rect 18521 21641 18555 21675
rect 22017 21641 22051 21675
rect 22661 21641 22695 21675
rect 25329 21641 25363 21675
rect 33793 21641 33827 21675
rect 2697 21573 2731 21607
rect 8769 21573 8803 21607
rect 13553 21573 13587 21607
rect 14105 21573 14139 21607
rect 17233 21573 17267 21607
rect 20913 21573 20947 21607
rect 21465 21573 21499 21607
rect 23673 21573 23707 21607
rect 24225 21573 24259 21607
rect 24777 21573 24811 21607
rect 1777 21505 1811 21539
rect 5089 21505 5123 21539
rect 5825 21505 5859 21539
rect 6745 21505 6779 21539
rect 7389 21505 7423 21539
rect 7849 21505 7883 21539
rect 10977 21505 11011 21539
rect 12909 21505 12943 21539
rect 14565 21505 14599 21539
rect 15853 21505 15887 21539
rect 18705 21505 18739 21539
rect 19257 21505 19291 21539
rect 20085 21505 20119 21539
rect 22201 21505 22235 21539
rect 22845 21505 22879 21539
rect 24685 21505 24719 21539
rect 25513 21505 25547 21539
rect 26157 21505 26191 21539
rect 33701 21505 33735 21539
rect 2421 21437 2455 21471
rect 4445 21437 4479 21471
rect 8493 21437 8527 21471
rect 13461 21437 13495 21471
rect 14749 21437 14783 21471
rect 15669 21437 15703 21471
rect 17141 21437 17175 21471
rect 20821 21437 20855 21471
rect 23581 21437 23615 21471
rect 11069 21369 11103 21403
rect 17693 21369 17727 21403
rect 19349 21369 19383 21403
rect 1593 21301 1627 21335
rect 4905 21301 4939 21335
rect 5917 21301 5951 21335
rect 7205 21301 7239 21335
rect 7941 21301 7975 21335
rect 10241 21301 10275 21335
rect 12725 21301 12759 21335
rect 14933 21301 14967 21335
rect 16037 21301 16071 21335
rect 20177 21301 20211 21335
rect 25973 21301 26007 21335
rect 4248 21097 4282 21131
rect 11989 21097 12023 21131
rect 16681 21097 16715 21131
rect 22753 21097 22787 21131
rect 27905 21097 27939 21131
rect 38117 21097 38151 21131
rect 8585 21029 8619 21063
rect 9597 21029 9631 21063
rect 14841 21029 14875 21063
rect 3985 20961 4019 20995
rect 6009 20961 6043 20995
rect 7113 20961 7147 20995
rect 10241 20961 10275 20995
rect 10517 20961 10551 20995
rect 12817 20961 12851 20995
rect 13461 20961 13495 20995
rect 14473 20961 14507 20995
rect 16497 20961 16531 20995
rect 20453 20961 20487 20995
rect 23581 20961 23615 20995
rect 24777 20961 24811 20995
rect 27169 20961 27203 20995
rect 1593 20893 1627 20927
rect 6837 20893 6871 20927
rect 9781 20893 9815 20927
rect 14657 20893 14691 20927
rect 15853 20893 15887 20927
rect 16313 20893 16347 20927
rect 19625 20893 19659 20927
rect 20269 20893 20303 20927
rect 21557 20893 21591 20927
rect 22293 20893 22327 20927
rect 22937 20893 22971 20927
rect 23397 20893 23431 20927
rect 24961 20893 24995 20927
rect 25881 20893 25915 20927
rect 26709 20893 26743 20927
rect 27813 20893 27847 20927
rect 38301 20893 38335 20927
rect 1869 20825 1903 20859
rect 12909 20825 12943 20859
rect 17693 20825 17727 20859
rect 17785 20825 17819 20859
rect 18337 20825 18371 20859
rect 3341 20757 3375 20791
rect 15669 20757 15703 20791
rect 19441 20757 19475 20791
rect 20913 20757 20947 20791
rect 21373 20757 21407 20791
rect 22109 20757 22143 20791
rect 24041 20757 24075 20791
rect 25421 20757 25455 20791
rect 25973 20757 26007 20791
rect 26525 20757 26559 20791
rect 11161 20553 11195 20587
rect 13921 20553 13955 20587
rect 16957 20553 16991 20587
rect 18797 20553 18831 20587
rect 22109 20553 22143 20587
rect 23673 20553 23707 20587
rect 25421 20553 25455 20587
rect 25881 20553 25915 20587
rect 1869 20485 1903 20519
rect 4537 20485 4571 20519
rect 13369 20485 13403 20519
rect 15393 20485 15427 20519
rect 17785 20485 17819 20519
rect 18337 20485 18371 20519
rect 3617 20417 3651 20451
rect 4261 20417 4295 20451
rect 9413 20417 9447 20451
rect 12173 20417 12207 20451
rect 12817 20417 12851 20451
rect 13277 20417 13311 20451
rect 14105 20417 14139 20451
rect 14749 20417 14783 20451
rect 18981 20417 19015 20451
rect 20177 20417 20211 20451
rect 20821 20417 20855 20451
rect 22293 20417 22327 20451
rect 22753 20417 22787 20451
rect 23857 20417 23891 20451
rect 24777 20417 24811 20451
rect 24961 20417 24995 20451
rect 26065 20417 26099 20451
rect 1593 20349 1627 20383
rect 6745 20349 6779 20383
rect 7021 20349 7055 20383
rect 8493 20349 8527 20383
rect 9689 20349 9723 20383
rect 15301 20349 15335 20383
rect 15577 20349 15611 20383
rect 17693 20349 17727 20383
rect 20637 20349 20671 20383
rect 6009 20213 6043 20247
rect 11989 20213 12023 20247
rect 12633 20213 12667 20247
rect 14565 20213 14599 20247
rect 19993 20213 20027 20247
rect 21281 20213 21315 20247
rect 22845 20213 22879 20247
rect 6837 20009 6871 20043
rect 9137 20009 9171 20043
rect 14565 20009 14599 20043
rect 17509 20009 17543 20043
rect 18153 20009 18187 20043
rect 21097 20009 21131 20043
rect 8309 19941 8343 19975
rect 9873 19941 9907 19975
rect 15577 19941 15611 19975
rect 16681 19941 16715 19975
rect 23673 19941 23707 19975
rect 25605 19941 25639 19975
rect 1869 19873 1903 19907
rect 5089 19873 5123 19907
rect 10425 19873 10459 19907
rect 13277 19873 13311 19907
rect 15393 19873 15427 19907
rect 16497 19873 16531 19907
rect 22845 19873 22879 19907
rect 25053 19873 25087 19907
rect 1593 19805 1627 19839
rect 4629 19805 4663 19839
rect 9321 19805 9355 19839
rect 9781 19805 9815 19839
rect 13093 19805 13127 19839
rect 14749 19805 14783 19839
rect 15209 19805 15243 19839
rect 16313 19805 16347 19839
rect 17417 19805 17451 19839
rect 18061 19805 18095 19839
rect 18889 19805 18923 19839
rect 19441 19805 19475 19839
rect 20545 19805 20579 19839
rect 21281 19805 21315 19839
rect 23305 19805 23339 19839
rect 23489 19805 23523 19839
rect 26341 19805 26375 19839
rect 5365 19737 5399 19771
rect 7757 19737 7791 19771
rect 7849 19737 7883 19771
rect 10701 19737 10735 19771
rect 22201 19737 22235 19771
rect 22293 19737 22327 19771
rect 25145 19737 25179 19771
rect 3341 19669 3375 19703
rect 4445 19669 4479 19703
rect 12173 19669 12207 19703
rect 13737 19669 13771 19703
rect 18705 19669 18739 19703
rect 19533 19669 19567 19703
rect 20361 19669 20395 19703
rect 26157 19669 26191 19703
rect 4721 19465 4755 19499
rect 8769 19465 8803 19499
rect 12449 19465 12483 19499
rect 20361 19465 20395 19499
rect 22937 19465 22971 19499
rect 24685 19465 24719 19499
rect 25881 19465 25915 19499
rect 3801 19397 3835 19431
rect 6745 19397 6779 19431
rect 8125 19397 8159 19431
rect 14381 19397 14415 19431
rect 21465 19397 21499 19431
rect 23581 19397 23615 19431
rect 4905 19329 4939 19363
rect 6009 19329 6043 19363
rect 8953 19329 8987 19363
rect 9413 19329 9447 19363
rect 11805 19329 11839 19363
rect 13093 19329 13127 19363
rect 13185 19329 13219 19363
rect 16865 19329 16899 19363
rect 18521 19329 18555 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 20821 19329 20855 19363
rect 24593 19329 24627 19363
rect 25421 19329 25455 19363
rect 26065 19329 26099 19363
rect 1777 19261 1811 19295
rect 2053 19261 2087 19295
rect 5365 19261 5399 19295
rect 5549 19261 5583 19295
rect 6653 19261 6687 19295
rect 11161 19261 11195 19295
rect 11989 19261 12023 19295
rect 13737 19261 13771 19295
rect 13921 19261 13955 19295
rect 15117 19261 15151 19295
rect 15301 19261 15335 19295
rect 17049 19261 17083 19295
rect 17509 19261 17543 19295
rect 18705 19261 18739 19295
rect 21005 19261 21039 19295
rect 22293 19261 22327 19295
rect 22477 19261 22511 19295
rect 23489 19261 23523 19295
rect 7205 19193 7239 19227
rect 15485 19193 15519 19227
rect 24041 19193 24075 19227
rect 9670 19125 9704 19159
rect 19165 19125 19199 19159
rect 25237 19125 25271 19159
rect 3341 18921 3375 18955
rect 9689 18921 9723 18955
rect 13737 18921 13771 18955
rect 14473 18921 14507 18955
rect 15485 18921 15519 18955
rect 5733 18853 5767 18887
rect 8217 18853 8251 18887
rect 12081 18853 12115 18887
rect 23949 18853 23983 18887
rect 3985 18785 4019 18819
rect 4261 18785 4295 18819
rect 7665 18785 7699 18819
rect 10333 18785 10367 18819
rect 13093 18785 13127 18819
rect 15301 18785 15335 18819
rect 17693 18785 17727 18819
rect 18429 18785 18463 18819
rect 19441 18785 19475 18819
rect 22385 18785 22419 18819
rect 23397 18785 23431 18819
rect 1593 18717 1627 18751
rect 7113 18717 7147 18751
rect 9873 18717 9907 18751
rect 13277 18717 13311 18751
rect 14657 18717 14691 18751
rect 15117 18717 15151 18751
rect 16497 18717 16531 18751
rect 17141 18717 17175 18751
rect 17601 18717 17635 18751
rect 18245 18717 18279 18751
rect 19625 18717 19659 18751
rect 20545 18717 20579 18751
rect 24593 18717 24627 18751
rect 25237 18717 25271 18751
rect 1869 18649 1903 18683
rect 6285 18649 6319 18683
rect 7750 18649 7784 18683
rect 10609 18649 10643 18683
rect 23489 18649 23523 18683
rect 6929 18581 6963 18615
rect 16313 18581 16347 18615
rect 16957 18581 16991 18615
rect 18889 18581 18923 18615
rect 20085 18581 20119 18615
rect 20637 18581 20671 18615
rect 24685 18581 24719 18615
rect 25329 18581 25363 18615
rect 1777 18377 1811 18411
rect 6837 18377 6871 18411
rect 9781 18377 9815 18411
rect 16129 18377 16163 18411
rect 21281 18377 21315 18411
rect 23949 18377 23983 18411
rect 24501 18377 24535 18411
rect 3341 18309 3375 18343
rect 7665 18309 7699 18343
rect 11897 18309 11931 18343
rect 14289 18309 14323 18343
rect 19165 18309 19199 18343
rect 19257 18309 19291 18343
rect 1593 18241 1627 18275
rect 3249 18241 3283 18275
rect 3893 18241 3927 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 6009 18241 6043 18275
rect 7021 18241 7055 18275
rect 9229 18241 9263 18275
rect 9689 18241 9723 18275
rect 10333 18241 10367 18275
rect 11161 18241 11195 18275
rect 13277 18241 13311 18275
rect 15117 18241 15151 18275
rect 15577 18241 15611 18275
rect 16313 18241 16347 18275
rect 17969 18241 18003 18275
rect 18153 18241 18187 18275
rect 21189 18241 21223 18275
rect 22109 18241 22143 18275
rect 22937 18241 22971 18275
rect 23857 18241 23891 18275
rect 24685 18241 24719 18275
rect 2605 18173 2639 18207
rect 7573 18173 7607 18207
rect 10425 18173 10459 18207
rect 11805 18173 11839 18207
rect 13093 18173 13127 18207
rect 14933 18173 14967 18207
rect 16865 18173 16899 18207
rect 17049 18173 17083 18207
rect 20177 18173 20211 18207
rect 22753 18173 22787 18207
rect 23397 18173 23431 18207
rect 3985 18105 4019 18139
rect 5181 18105 5215 18139
rect 5825 18105 5859 18139
rect 8125 18105 8159 18139
rect 9045 18105 9079 18139
rect 12357 18105 12391 18139
rect 4537 18037 4571 18071
rect 10977 18037 11011 18071
rect 13461 18037 13495 18071
rect 17509 18037 17543 18071
rect 18613 18037 18647 18071
rect 22201 18037 22235 18071
rect 9689 17833 9723 17867
rect 11897 17833 11931 17867
rect 19441 17833 19475 17867
rect 2053 17765 2087 17799
rect 4537 17765 4571 17799
rect 5825 17765 5859 17799
rect 8217 17765 8251 17799
rect 11161 17765 11195 17799
rect 17141 17765 17175 17799
rect 20085 17765 20119 17799
rect 23949 17765 23983 17799
rect 6469 17697 6503 17731
rect 6653 17697 6687 17731
rect 7665 17697 7699 17731
rect 9137 17697 9171 17731
rect 9321 17697 9355 17731
rect 12633 17697 12667 17731
rect 13093 17697 13127 17731
rect 13553 17697 13587 17731
rect 14473 17697 14507 17731
rect 15577 17697 15611 17731
rect 16589 17697 16623 17731
rect 17693 17697 17727 17731
rect 17877 17697 17911 17731
rect 1961 17629 1995 17663
rect 2789 17629 2823 17663
rect 3433 17629 3467 17663
rect 4721 17629 4755 17663
rect 10517 17629 10551 17663
rect 11345 17629 11379 17663
rect 11805 17629 11839 17663
rect 12449 17629 12483 17663
rect 14289 17629 14323 17663
rect 15393 17629 15427 17663
rect 19625 17629 19659 17663
rect 20269 17629 20303 17663
rect 21373 17629 21407 17663
rect 24593 17629 24627 17663
rect 5273 17561 5307 17595
rect 5365 17561 5399 17595
rect 7757 17561 7791 17595
rect 10609 17561 10643 17595
rect 16681 17561 16715 17595
rect 23397 17561 23431 17595
rect 23489 17561 23523 17595
rect 2605 17493 2639 17527
rect 3249 17493 3283 17527
rect 7113 17493 7147 17527
rect 14933 17493 14967 17527
rect 16037 17493 16071 17527
rect 18337 17493 18371 17527
rect 21189 17493 21223 17527
rect 24685 17493 24719 17527
rect 16221 17289 16255 17323
rect 18153 17289 18187 17323
rect 18797 17289 18831 17323
rect 22845 17289 22879 17323
rect 38117 17289 38151 17323
rect 3157 17221 3191 17255
rect 8861 17221 8895 17255
rect 9689 17221 9723 17255
rect 14749 17221 14783 17255
rect 1593 17153 1627 17187
rect 6009 17153 6043 17187
rect 8769 17153 8803 17187
rect 9413 17153 9447 17187
rect 14105 17153 14139 17187
rect 16129 17153 16163 17187
rect 17049 17153 17083 17187
rect 18981 17153 19015 17187
rect 19625 17153 19659 17187
rect 20085 17153 20119 17187
rect 21465 17153 21499 17187
rect 22385 17153 22419 17187
rect 23489 17153 23523 17187
rect 24409 17153 24443 17187
rect 25881 17153 25915 17187
rect 33701 17153 33735 17187
rect 38301 17153 38335 17187
rect 2881 17085 2915 17119
rect 4905 17085 4939 17119
rect 6561 17085 6595 17119
rect 6837 17085 6871 17119
rect 12265 17085 12299 17119
rect 12449 17085 12483 17119
rect 14657 17085 14691 17119
rect 15301 17085 15335 17119
rect 17509 17085 17543 17119
rect 17693 17085 17727 17119
rect 22201 17085 22235 17119
rect 23305 17085 23339 17119
rect 25053 17085 25087 17119
rect 33793 17017 33827 17051
rect 1777 16949 1811 16983
rect 5825 16949 5859 16983
rect 8309 16949 8343 16983
rect 11161 16949 11195 16983
rect 12633 16949 12667 16983
rect 13921 16949 13955 16983
rect 16865 16949 16899 16983
rect 19441 16949 19475 16983
rect 20177 16949 20211 16983
rect 21281 16949 21315 16983
rect 23673 16949 23707 16983
rect 24501 16949 24535 16983
rect 25697 16949 25731 16983
rect 16681 16745 16715 16779
rect 18337 16745 18371 16779
rect 20085 16745 20119 16779
rect 21557 16745 21591 16779
rect 23213 16745 23247 16779
rect 1961 16609 1995 16643
rect 4261 16609 4295 16643
rect 6929 16609 6963 16643
rect 7573 16609 7607 16643
rect 10885 16609 10919 16643
rect 12081 16609 12115 16643
rect 16497 16609 16531 16643
rect 17969 16609 18003 16643
rect 18153 16609 18187 16643
rect 21189 16609 21223 16643
rect 21373 16609 21407 16643
rect 22569 16609 22603 16643
rect 24593 16609 24627 16643
rect 1685 16541 1719 16575
rect 3985 16541 4019 16575
rect 9137 16541 9171 16575
rect 11621 16541 11655 16575
rect 12265 16541 12299 16575
rect 14473 16541 14507 16575
rect 16313 16541 16347 16575
rect 19625 16541 19659 16575
rect 20269 16541 20303 16575
rect 22753 16541 22787 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 6285 16473 6319 16507
rect 6377 16473 6411 16507
rect 7665 16473 7699 16507
rect 8217 16473 8251 16507
rect 9413 16473 9447 16507
rect 15209 16473 15243 16507
rect 15301 16473 15335 16507
rect 15853 16473 15887 16507
rect 3433 16405 3467 16439
rect 5733 16405 5767 16439
rect 11437 16405 11471 16439
rect 12725 16405 12759 16439
rect 13553 16405 13587 16439
rect 14565 16405 14599 16439
rect 19441 16405 19475 16439
rect 23673 16405 23707 16439
rect 25237 16405 25271 16439
rect 11161 16201 11195 16235
rect 13277 16201 13311 16235
rect 22017 16201 22051 16235
rect 22753 16201 22787 16235
rect 24041 16201 24075 16235
rect 24501 16201 24535 16235
rect 3617 16133 3651 16167
rect 7481 16133 7515 16167
rect 14105 16133 14139 16167
rect 18337 16133 18371 16167
rect 18889 16133 18923 16167
rect 19533 16133 19567 16167
rect 20085 16133 20119 16167
rect 6561 16065 6595 16099
rect 9413 16065 9447 16099
rect 13461 16065 13495 16099
rect 16865 16065 16899 16099
rect 20729 16065 20763 16099
rect 22201 16065 22235 16099
rect 22937 16065 22971 16099
rect 24685 16065 24719 16099
rect 29745 16065 29779 16099
rect 38025 16065 38059 16099
rect 1593 15997 1627 16031
rect 1869 15997 1903 16031
rect 4077 15997 4111 16031
rect 4353 15997 4387 16031
rect 5825 15997 5859 16031
rect 7194 15997 7228 16031
rect 9689 15997 9723 16031
rect 11713 15997 11747 16031
rect 11897 15997 11931 16031
rect 14013 15997 14047 16031
rect 15117 15997 15151 16031
rect 15301 15997 15335 16031
rect 17049 15997 17083 16031
rect 18245 15997 18279 16031
rect 19441 15997 19475 16031
rect 20545 15997 20579 16031
rect 23397 15997 23431 16031
rect 23581 15997 23615 16031
rect 14565 15929 14599 15963
rect 6653 15861 6687 15895
rect 8953 15861 8987 15895
rect 12081 15861 12115 15895
rect 15485 15861 15519 15895
rect 17233 15861 17267 15895
rect 20913 15861 20947 15895
rect 29837 15861 29871 15895
rect 38209 15861 38243 15895
rect 3433 15657 3467 15691
rect 11345 15657 11379 15691
rect 13645 15657 13679 15691
rect 14565 15657 14599 15691
rect 20269 15657 20303 15691
rect 6653 15589 6687 15623
rect 9965 15589 9999 15623
rect 16865 15589 16899 15623
rect 2145 15521 2179 15555
rect 2789 15521 2823 15555
rect 2973 15521 3007 15555
rect 5181 15521 5215 15555
rect 7665 15521 7699 15555
rect 9781 15521 9815 15555
rect 10977 15521 11011 15555
rect 12081 15521 12115 15555
rect 17693 15521 17727 15555
rect 17969 15521 18003 15555
rect 19809 15521 19843 15555
rect 20913 15521 20947 15555
rect 22293 15521 22327 15555
rect 1869 15453 1903 15487
rect 3985 15453 4019 15487
rect 4905 15453 4939 15487
rect 9597 15453 9631 15487
rect 11161 15453 11195 15487
rect 12265 15453 12299 15487
rect 13553 15453 13587 15487
rect 14749 15453 14783 15487
rect 16497 15453 16531 15487
rect 16681 15453 16715 15487
rect 19625 15453 19659 15487
rect 20729 15453 20763 15487
rect 22477 15453 22511 15487
rect 24593 15453 24627 15487
rect 4261 15385 4295 15419
rect 7757 15385 7791 15419
rect 8309 15385 8343 15419
rect 15301 15385 15335 15419
rect 15393 15385 15427 15419
rect 15945 15385 15979 15419
rect 17785 15385 17819 15419
rect 12725 15317 12759 15351
rect 21373 15317 21407 15351
rect 22937 15317 22971 15351
rect 23397 15317 23431 15351
rect 24685 15317 24719 15351
rect 10609 15113 10643 15147
rect 14473 15113 14507 15147
rect 15761 15113 15795 15147
rect 18613 15113 18647 15147
rect 22937 15113 22971 15147
rect 34713 15113 34747 15147
rect 3801 15045 3835 15079
rect 6837 15045 6871 15079
rect 17417 15045 17451 15079
rect 19257 15045 19291 15079
rect 19349 15045 19383 15079
rect 4261 14977 4295 15011
rect 8861 14977 8895 15011
rect 13001 14977 13035 15011
rect 14657 14977 14691 15011
rect 18521 14977 18555 15011
rect 19901 14977 19935 15011
rect 22293 14977 22327 15011
rect 23581 14977 23615 15011
rect 24041 14977 24075 15011
rect 24869 14977 24903 15011
rect 33517 14977 33551 15011
rect 34897 14977 34931 15011
rect 35541 14977 35575 15011
rect 1777 14909 1811 14943
rect 2053 14909 2087 14943
rect 4537 14909 4571 14943
rect 6561 14909 6595 14943
rect 9137 14909 9171 14943
rect 11713 14909 11747 14943
rect 11897 14909 11931 14943
rect 12817 14909 12851 14943
rect 15117 14909 15151 14943
rect 15301 14909 15335 14943
rect 17325 14909 17359 14943
rect 20545 14909 20579 14943
rect 20729 14909 20763 14943
rect 22477 14909 22511 14943
rect 25329 14909 25363 14943
rect 25513 14909 25547 14943
rect 17877 14841 17911 14875
rect 23397 14841 23431 14875
rect 24133 14841 24167 14875
rect 24685 14841 24719 14875
rect 33609 14841 33643 14875
rect 6009 14773 6043 14807
rect 8309 14773 8343 14807
rect 12081 14773 12115 14807
rect 13185 14773 13219 14807
rect 20913 14773 20947 14807
rect 25697 14773 25731 14807
rect 35357 14773 35391 14807
rect 3433 14569 3467 14603
rect 6377 14569 6411 14603
rect 15577 14569 15611 14603
rect 18429 14569 18463 14603
rect 30021 14569 30055 14603
rect 3801 14501 3835 14535
rect 14657 14501 14691 14535
rect 25237 14501 25271 14535
rect 26065 14501 26099 14535
rect 1961 14433 1995 14467
rect 9137 14433 9171 14467
rect 9413 14433 9447 14467
rect 10885 14433 10919 14467
rect 11437 14433 11471 14467
rect 13645 14433 13679 14467
rect 14473 14433 14507 14467
rect 16129 14433 16163 14467
rect 17325 14433 17359 14467
rect 17785 14433 17819 14467
rect 19533 14433 19567 14467
rect 20637 14433 20671 14467
rect 21741 14433 21775 14467
rect 23029 14433 23063 14467
rect 23213 14433 23247 14467
rect 33793 14433 33827 14467
rect 1685 14365 1719 14399
rect 3985 14365 4019 14399
rect 4629 14365 4663 14399
rect 6837 14365 6871 14399
rect 13001 14365 13035 14399
rect 13185 14365 13219 14399
rect 14289 14365 14323 14399
rect 15485 14365 15519 14399
rect 16313 14365 16347 14399
rect 18613 14365 18647 14399
rect 21925 14365 21959 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 25697 14365 25731 14399
rect 25881 14365 25915 14399
rect 26985 14365 27019 14399
rect 29929 14365 29963 14399
rect 33701 14365 33735 14399
rect 38301 14365 38335 14399
rect 4353 14297 4387 14331
rect 4905 14297 4939 14331
rect 7113 14297 7147 14331
rect 11529 14297 11563 14331
rect 12081 14297 12115 14331
rect 17417 14297 17451 14331
rect 20729 14297 20763 14331
rect 21281 14297 21315 14331
rect 8585 14229 8619 14263
rect 16773 14229 16807 14263
rect 22385 14229 22419 14263
rect 23673 14229 23707 14263
rect 26801 14229 26835 14263
rect 38117 14229 38151 14263
rect 1685 14025 1719 14059
rect 5825 14025 5859 14059
rect 7573 14025 7607 14059
rect 11161 14025 11195 14059
rect 13185 14025 13219 14059
rect 15761 14025 15795 14059
rect 18153 14025 18187 14059
rect 19441 14025 19475 14059
rect 20085 14025 20119 14059
rect 22109 14025 22143 14059
rect 23857 14025 23891 14059
rect 25329 14025 25363 14059
rect 26525 14025 26559 14059
rect 12357 13957 12391 13991
rect 13921 13957 13955 13991
rect 14013 13957 14047 13991
rect 14565 13957 14599 13991
rect 17049 13957 17083 13991
rect 17601 13957 17635 13991
rect 20913 13957 20947 13991
rect 2329 13889 2363 13923
rect 6009 13889 6043 13923
rect 8217 13889 8251 13923
rect 10517 13889 10551 13923
rect 13369 13889 13403 13923
rect 18337 13889 18371 13923
rect 18797 13889 18831 13923
rect 19625 13889 19659 13923
rect 22293 13889 22327 13923
rect 23213 13889 23247 13923
rect 25789 13889 25823 13923
rect 26433 13889 26467 13923
rect 2513 13821 2547 13855
rect 3249 13821 3283 13855
rect 3525 13821 3559 13855
rect 5273 13821 5307 13855
rect 6929 13821 6963 13855
rect 7113 13821 7147 13855
rect 8493 13821 8527 13855
rect 9965 13821 9999 13855
rect 10701 13821 10735 13855
rect 11713 13821 11747 13855
rect 11897 13821 11931 13855
rect 15117 13821 15151 13855
rect 15301 13821 15335 13855
rect 16957 13821 16991 13855
rect 18889 13821 18923 13855
rect 20821 13821 20855 13855
rect 21465 13821 21499 13855
rect 23397 13821 23431 13855
rect 24685 13821 24719 13855
rect 24869 13821 24903 13855
rect 25881 13821 25915 13855
rect 3433 13481 3467 13515
rect 4248 13481 4282 13515
rect 13645 13481 13679 13515
rect 14749 13481 14783 13515
rect 15669 13481 15703 13515
rect 21925 13481 21959 13515
rect 22569 13481 22603 13515
rect 25881 13481 25915 13515
rect 26525 13481 26559 13515
rect 17417 13413 17451 13447
rect 18889 13413 18923 13447
rect 19809 13413 19843 13447
rect 21373 13413 21407 13447
rect 1961 13345 1995 13379
rect 6745 13345 6779 13379
rect 7021 13345 7055 13379
rect 9137 13345 9171 13379
rect 11345 13345 11379 13379
rect 14289 13345 14323 13379
rect 20821 13345 20855 13379
rect 23305 13345 23339 13379
rect 24593 13345 24627 13379
rect 1685 13277 1719 13311
rect 3985 13277 4019 13311
rect 11529 13277 11563 13311
rect 11989 13277 12023 13311
rect 12449 13277 12483 13311
rect 12633 13277 12667 13311
rect 13553 13277 13587 13311
rect 14473 13277 14507 13311
rect 15577 13277 15611 13311
rect 17601 13277 17635 13311
rect 18245 13277 18279 13311
rect 18429 13277 18463 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 21005 13277 21039 13311
rect 22109 13277 22143 13311
rect 22753 13277 22787 13311
rect 25421 13277 25455 13311
rect 26065 13277 26099 13311
rect 26709 13277 26743 13311
rect 6009 13209 6043 13243
rect 9413 13209 9447 13243
rect 16313 13209 16347 13243
rect 16405 13209 16439 13243
rect 16957 13209 16991 13243
rect 23397 13209 23431 13243
rect 23949 13209 23983 13243
rect 8493 13141 8527 13175
rect 10885 13141 10919 13175
rect 13093 13141 13127 13175
rect 25237 13141 25271 13175
rect 10793 12937 10827 12971
rect 16957 12937 16991 12971
rect 18153 12937 18187 12971
rect 19073 12937 19107 12971
rect 19809 12937 19843 12971
rect 21281 12937 21315 12971
rect 22385 12937 22419 12971
rect 24225 12937 24259 12971
rect 25605 12937 25639 12971
rect 1869 12869 1903 12903
rect 4353 12869 4387 12903
rect 6837 12869 6871 12903
rect 12541 12869 12575 12903
rect 13737 12869 13771 12903
rect 14933 12869 14967 12903
rect 23121 12869 23155 12903
rect 23213 12869 23247 12903
rect 24961 12869 24995 12903
rect 4077 12801 4111 12835
rect 6561 12801 6595 12835
rect 9229 12801 9263 12835
rect 10149 12801 10183 12835
rect 11713 12801 11747 12835
rect 18337 12801 18371 12835
rect 19257 12801 19291 12835
rect 19717 12801 19751 12835
rect 20637 12801 20671 12835
rect 22569 12801 22603 12835
rect 24409 12801 24443 12835
rect 24869 12801 24903 12835
rect 25789 12801 25823 12835
rect 38025 12801 38059 12835
rect 1593 12733 1627 12767
rect 3617 12733 3651 12767
rect 8309 12733 8343 12767
rect 9045 12733 9079 12767
rect 10333 12733 10367 12767
rect 12449 12733 12483 12767
rect 13645 12733 13679 12767
rect 15577 12733 15611 12767
rect 15761 12733 15795 12767
rect 20821 12733 20855 12767
rect 23765 12733 23799 12767
rect 5825 12665 5859 12699
rect 13001 12665 13035 12699
rect 14197 12665 14231 12699
rect 9413 12597 9447 12631
rect 11805 12597 11839 12631
rect 15945 12597 15979 12631
rect 38209 12597 38243 12631
rect 3433 12393 3467 12427
rect 4077 12393 4111 12427
rect 16773 12393 16807 12427
rect 17417 12393 17451 12427
rect 20177 12393 20211 12427
rect 23029 12393 23063 12427
rect 24593 12393 24627 12427
rect 30665 12393 30699 12427
rect 8585 12325 8619 12359
rect 10425 12325 10459 12359
rect 11529 12325 11563 12359
rect 16037 12325 16071 12359
rect 18061 12325 18095 12359
rect 1961 12257 1995 12291
rect 4721 12257 4755 12291
rect 6745 12257 6779 12291
rect 7297 12257 7331 12291
rect 7941 12257 7975 12291
rect 10057 12257 10091 12291
rect 11161 12257 11195 12291
rect 18705 12257 18739 12291
rect 20913 12257 20947 12291
rect 22385 12257 22419 12291
rect 22569 12257 22603 12291
rect 23581 12257 23615 12291
rect 1685 12189 1719 12223
rect 3985 12189 4019 12223
rect 8125 12189 8159 12223
rect 9597 12189 9631 12223
rect 10241 12189 10275 12223
rect 11345 12189 11379 12223
rect 12541 12189 12575 12223
rect 13737 12189 13771 12223
rect 16221 12189 16255 12223
rect 16681 12189 16715 12223
rect 17601 12189 17635 12223
rect 18245 12189 18279 12223
rect 19717 12189 19751 12223
rect 20361 12189 20395 12223
rect 23489 12189 23523 12223
rect 24777 12189 24811 12223
rect 25421 12189 25455 12223
rect 30573 12189 30607 12223
rect 4997 12121 5031 12155
rect 13093 12121 13127 12155
rect 13194 12121 13228 12155
rect 14381 12121 14415 12155
rect 14473 12121 14507 12155
rect 15025 12121 15059 12155
rect 21005 12121 21039 12155
rect 21557 12121 21591 12155
rect 9413 12053 9447 12087
rect 12357 12053 12391 12087
rect 19533 12053 19567 12087
rect 25237 12053 25271 12087
rect 7205 11849 7239 11883
rect 10609 11849 10643 11883
rect 12357 11849 12391 11883
rect 13369 11849 13403 11883
rect 15301 11849 15335 11883
rect 16129 11849 16163 11883
rect 16865 11849 16899 11883
rect 19073 11849 19107 11883
rect 19625 11849 19659 11883
rect 20453 11849 20487 11883
rect 22017 11849 22051 11883
rect 2881 11781 2915 11815
rect 4629 11781 4663 11815
rect 14657 11781 14691 11815
rect 21189 11781 21223 11815
rect 1685 11713 1719 11747
rect 6009 11697 6043 11731
rect 7113 11713 7147 11747
rect 9965 11713 9999 11747
rect 13277 11713 13311 11747
rect 14105 11713 14139 11747
rect 14565 11713 14599 11747
rect 15209 11713 15243 11747
rect 16313 11713 16347 11747
rect 17693 11713 17727 11747
rect 18981 11713 19015 11747
rect 19809 11713 19843 11747
rect 20637 11713 20671 11747
rect 21097 11713 21131 11747
rect 22201 11713 22235 11747
rect 22845 11713 22879 11747
rect 1869 11645 1903 11679
rect 2605 11645 2639 11679
rect 5181 11645 5215 11679
rect 7757 11645 7791 11679
rect 8033 11645 8067 11679
rect 10149 11645 10183 11679
rect 11713 11645 11747 11679
rect 11897 11645 11931 11679
rect 18245 11645 18279 11679
rect 9505 11577 9539 11611
rect 17509 11577 17543 11611
rect 22661 11577 22695 11611
rect 5825 11509 5859 11543
rect 13921 11509 13955 11543
rect 3433 11305 3467 11339
rect 7297 11305 7331 11339
rect 11621 11305 11655 11339
rect 12357 11305 12391 11339
rect 13185 11305 13219 11339
rect 15761 11305 15795 11339
rect 18521 11305 18555 11339
rect 20729 11305 20763 11339
rect 38117 11305 38151 11339
rect 15117 11237 15151 11271
rect 4905 11169 4939 11203
rect 7849 11169 7883 11203
rect 8033 11169 8067 11203
rect 9965 11169 9999 11203
rect 16405 11169 16439 11203
rect 18153 11169 18187 11203
rect 20177 11169 20211 11203
rect 21649 11169 21683 11203
rect 22477 11169 22511 11203
rect 1685 11101 1719 11135
rect 4261 11101 4295 11135
rect 7205 11101 7239 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 10425 11101 10459 11135
rect 10609 11101 10643 11135
rect 11529 11101 11563 11135
rect 12541 11101 12575 11135
rect 13093 11101 13127 11135
rect 14473 11101 14507 11135
rect 15301 11101 15335 11135
rect 15945 11101 15979 11135
rect 16589 11101 16623 11135
rect 17693 11101 17727 11135
rect 18337 11101 18371 11135
rect 20637 11101 20671 11135
rect 38301 11101 38335 11135
rect 1961 11033 1995 11067
rect 4353 11033 4387 11067
rect 5181 11033 5215 11067
rect 8493 11033 8527 11067
rect 11069 11033 11103 11067
rect 17049 11033 17083 11067
rect 19533 11033 19567 11067
rect 19625 11033 19659 11067
rect 21373 11033 21407 11067
rect 21465 11033 21499 11067
rect 6653 10965 6687 10999
rect 14289 10965 14323 10999
rect 17509 10965 17543 10999
rect 1777 10761 1811 10795
rect 2421 10761 2455 10795
rect 3065 10761 3099 10795
rect 4077 10761 4111 10795
rect 7573 10761 7607 10795
rect 13553 10761 13587 10795
rect 14749 10761 14783 10795
rect 15301 10761 15335 10795
rect 15945 10761 15979 10795
rect 16865 10761 16899 10795
rect 19625 10761 19659 10795
rect 21097 10761 21131 10795
rect 6929 10693 6963 10727
rect 9689 10693 9723 10727
rect 12265 10693 12299 10727
rect 12357 10693 12391 10727
rect 1685 10625 1719 10659
rect 2329 10625 2363 10659
rect 2973 10625 3007 10659
rect 3985 10625 4019 10659
rect 5181 10625 5215 10659
rect 6009 10625 6043 10659
rect 6837 10625 6871 10659
rect 7481 10625 7515 10659
rect 8125 10625 8159 10659
rect 8953 10625 8987 10659
rect 9413 10625 9447 10659
rect 13461 10625 13495 10659
rect 14657 10625 14691 10659
rect 16129 10625 16163 10659
rect 17049 10625 17083 10659
rect 17969 10625 18003 10659
rect 19533 10625 19567 10659
rect 21281 10625 21315 10659
rect 22753 10625 22787 10659
rect 27169 10625 27203 10659
rect 27261 10625 27295 10659
rect 28549 10625 28583 10659
rect 33793 10625 33827 10659
rect 5273 10557 5307 10591
rect 8217 10557 8251 10591
rect 18429 10557 18463 10591
rect 18613 10557 18647 10591
rect 12817 10489 12851 10523
rect 18797 10489 18831 10523
rect 28641 10489 28675 10523
rect 5825 10421 5859 10455
rect 8769 10421 8803 10455
rect 11161 10421 11195 10455
rect 17785 10421 17819 10455
rect 22845 10421 22879 10455
rect 33885 10421 33919 10455
rect 2053 10217 2087 10251
rect 3341 10217 3375 10251
rect 4077 10217 4111 10251
rect 4892 10217 4926 10251
rect 7205 10217 7239 10251
rect 8401 10217 8435 10251
rect 12173 10217 12207 10251
rect 12817 10217 12851 10251
rect 14289 10217 14323 10251
rect 15577 10217 15611 10251
rect 18521 10217 18555 10251
rect 19533 10217 19567 10251
rect 20545 10217 20579 10251
rect 33977 10217 34011 10251
rect 2697 10149 2731 10183
rect 11529 10149 11563 10183
rect 14933 10149 14967 10183
rect 4629 10081 4663 10115
rect 9229 10081 9263 10115
rect 9505 10081 9539 10115
rect 13553 10081 13587 10115
rect 1961 10013 1995 10047
rect 2605 10013 2639 10047
rect 3249 10013 3283 10047
rect 3985 10013 4019 10047
rect 7113 10013 7147 10047
rect 7757 10013 7791 10047
rect 8585 10013 8619 10047
rect 11713 10013 11747 10047
rect 12357 10013 12391 10047
rect 13001 10013 13035 10047
rect 13461 10013 13495 10047
rect 14473 10013 14507 10047
rect 15117 10013 15151 10047
rect 15761 10013 15795 10047
rect 16773 10013 16807 10047
rect 18705 10013 18739 10047
rect 19441 10013 19475 10047
rect 20729 10013 20763 10047
rect 28273 10013 28307 10047
rect 29745 10013 29779 10047
rect 33885 10013 33919 10047
rect 6377 9877 6411 9911
rect 10977 9877 11011 9911
rect 16865 9877 16899 9911
rect 28365 9877 28399 9911
rect 29837 9877 29871 9911
rect 1869 9605 1903 9639
rect 2513 9605 2547 9639
rect 11069 9605 11103 9639
rect 12541 9605 12575 9639
rect 13093 9605 13127 9639
rect 14565 9605 14599 9639
rect 1777 9537 1811 9571
rect 2421 9537 2455 9571
rect 5549 9537 5583 9571
rect 5641 9537 5675 9571
rect 6561 9537 6595 9571
rect 9229 9537 9263 9571
rect 9873 9537 9907 9571
rect 10517 9537 10551 9571
rect 10977 9537 11011 9571
rect 12081 9537 12115 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 14473 9537 14507 9571
rect 15301 9537 15335 9571
rect 34529 9537 34563 9571
rect 3065 9469 3099 9503
rect 3341 9469 3375 9503
rect 5089 9469 5123 9503
rect 6837 9469 6871 9503
rect 11897 9469 11931 9503
rect 8309 9401 8343 9435
rect 9689 9401 9723 9435
rect 10333 9401 10367 9435
rect 9045 9333 9079 9367
rect 13829 9333 13863 9367
rect 15117 9333 15151 9367
rect 34345 9333 34379 9367
rect 7100 9129 7134 9163
rect 9689 9129 9723 9163
rect 12081 9129 12115 9163
rect 12633 9129 12667 9163
rect 14933 9129 14967 9163
rect 25237 9129 25271 9163
rect 3341 9061 3375 9095
rect 8585 9061 8619 9095
rect 14381 9061 14415 9095
rect 1869 8993 1903 9027
rect 4353 8993 4387 9027
rect 6837 8993 6871 9027
rect 10609 8993 10643 9027
rect 1593 8925 1627 8959
rect 9873 8925 9907 8959
rect 10333 8925 10367 8959
rect 12541 8925 12575 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 15117 8925 15151 8959
rect 25145 8925 25179 8959
rect 38025 8925 38059 8959
rect 4629 8857 4663 8891
rect 6377 8857 6411 8891
rect 13185 8789 13219 8823
rect 38209 8789 38243 8823
rect 1685 8585 1719 8619
rect 4629 8585 4663 8619
rect 5273 8585 5307 8619
rect 5917 8585 5951 8619
rect 9413 8585 9447 8619
rect 10333 8585 10367 8619
rect 11069 8585 11103 8619
rect 11805 8585 11839 8619
rect 12357 8585 12391 8619
rect 13001 8585 13035 8619
rect 14013 8585 14047 8619
rect 14749 8585 14783 8619
rect 2513 8517 2547 8551
rect 1593 8449 1627 8483
rect 4537 8449 4571 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 7021 8449 7055 8483
rect 10517 8449 10551 8483
rect 10977 8449 11011 8483
rect 11713 8449 11747 8483
rect 12541 8449 12575 8483
rect 13185 8449 13219 8483
rect 14197 8449 14231 8483
rect 14657 8449 14691 8483
rect 20177 8449 20211 8483
rect 21189 8449 21223 8483
rect 33977 8449 34011 8483
rect 2237 8381 2271 8415
rect 3985 8381 4019 8415
rect 7665 8381 7699 8415
rect 7941 8381 7975 8415
rect 21281 8381 21315 8415
rect 7113 8313 7147 8347
rect 20269 8313 20303 8347
rect 34069 8313 34103 8347
rect 4721 8041 4755 8075
rect 7941 8041 7975 8075
rect 9781 8041 9815 8075
rect 12725 8041 12759 8075
rect 13277 8041 13311 8075
rect 27997 8041 28031 8075
rect 38117 8041 38151 8075
rect 3341 7973 3375 8007
rect 4077 7973 4111 8007
rect 6193 7905 6227 7939
rect 1593 7837 1627 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 5273 7837 5307 7871
rect 9689 7837 9723 7871
rect 10333 7837 10367 7871
rect 12633 7837 12667 7871
rect 13461 7837 13495 7871
rect 27905 7837 27939 7871
rect 38301 7837 38335 7871
rect 1869 7769 1903 7803
rect 5365 7769 5399 7803
rect 6469 7769 6503 7803
rect 10609 7769 10643 7803
rect 12081 7701 12115 7735
rect 3433 7497 3467 7531
rect 5365 7497 5399 7531
rect 6653 7497 6687 7531
rect 13461 7497 13495 7531
rect 1961 7429 1995 7463
rect 4077 7429 4111 7463
rect 7481 7429 7515 7463
rect 9689 7429 9723 7463
rect 1685 7361 1719 7395
rect 3985 7361 4019 7395
rect 4629 7361 4663 7395
rect 5273 7361 5307 7395
rect 6561 7361 6595 7395
rect 7205 7361 7239 7395
rect 9413 7361 9447 7395
rect 11713 7361 11747 7395
rect 16865 7361 16899 7395
rect 36369 7361 36403 7395
rect 11989 7293 12023 7327
rect 4721 7225 4755 7259
rect 8953 7157 8987 7191
rect 11161 7157 11195 7191
rect 16957 7157 16991 7191
rect 36185 7157 36219 7191
rect 10406 6953 10440 6987
rect 6009 6817 6043 6851
rect 6653 6817 6687 6851
rect 10149 6817 10183 6851
rect 12541 6817 12575 6851
rect 25421 6817 25455 6851
rect 1777 6749 1811 6783
rect 2329 6749 2363 6783
rect 2973 6749 3007 6783
rect 3985 6749 4019 6783
rect 4077 6749 4111 6783
rect 4629 6749 4663 6783
rect 5273 6749 5307 6783
rect 5917 6749 5951 6783
rect 6561 6749 6595 6783
rect 7573 6749 7607 6783
rect 8217 6749 8251 6783
rect 8309 6749 8343 6783
rect 9321 6749 9355 6783
rect 12449 6749 12483 6783
rect 25329 6749 25363 6783
rect 34161 6749 34195 6783
rect 1593 6613 1627 6647
rect 2421 6613 2455 6647
rect 3065 6613 3099 6647
rect 4721 6613 4755 6647
rect 5365 6613 5399 6647
rect 7665 6613 7699 6647
rect 9137 6613 9171 6647
rect 11897 6613 11931 6647
rect 33977 6613 34011 6647
rect 1593 6409 1627 6443
rect 2513 6409 2547 6443
rect 3157 6409 3191 6443
rect 3801 6409 3835 6443
rect 6653 6409 6687 6443
rect 7757 6409 7791 6443
rect 8401 6409 8435 6443
rect 10701 6409 10735 6443
rect 13921 6409 13955 6443
rect 18429 6409 18463 6443
rect 22109 6409 22143 6443
rect 38117 6409 38151 6443
rect 1777 6273 1811 6307
rect 2421 6273 2455 6307
rect 3065 6273 3099 6307
rect 3709 6273 3743 6307
rect 4629 6273 4663 6307
rect 5273 6273 5307 6307
rect 6561 6273 6595 6307
rect 7665 6273 7699 6307
rect 8309 6273 8343 6307
rect 8953 6273 8987 6307
rect 13829 6273 13863 6307
rect 18337 6273 18371 6307
rect 22017 6273 22051 6307
rect 31033 6273 31067 6307
rect 32965 6273 32999 6307
rect 38301 6273 38335 6307
rect 5365 6205 5399 6239
rect 9229 6205 9263 6239
rect 33057 6205 33091 6239
rect 31125 6137 31159 6171
rect 4721 6069 4755 6103
rect 2421 5865 2455 5899
rect 4077 5865 4111 5899
rect 4721 5865 4755 5899
rect 5365 5865 5399 5899
rect 6009 5865 6043 5899
rect 11253 5865 11287 5899
rect 1777 5797 1811 5831
rect 6653 5797 6687 5831
rect 8125 5797 8159 5831
rect 7297 5729 7331 5763
rect 1685 5661 1719 5695
rect 2329 5661 2363 5695
rect 3157 5661 3191 5695
rect 3985 5661 4019 5695
rect 4629 5661 4663 5695
rect 5273 5661 5307 5695
rect 5917 5661 5951 5695
rect 6561 5661 6595 5695
rect 7205 5661 7239 5695
rect 8033 5661 8067 5695
rect 11161 5661 11195 5695
rect 11989 5661 12023 5695
rect 17877 5661 17911 5695
rect 18521 5661 18555 5695
rect 21189 5661 21223 5695
rect 23581 5661 23615 5695
rect 3249 5593 3283 5627
rect 12081 5593 12115 5627
rect 17693 5525 17727 5559
rect 18337 5525 18371 5559
rect 21005 5525 21039 5559
rect 23397 5525 23431 5559
rect 2421 5321 2455 5355
rect 3709 5321 3743 5355
rect 4353 5321 4387 5355
rect 4997 5321 5031 5355
rect 3065 5253 3099 5287
rect 8861 5253 8895 5287
rect 1593 5185 1627 5219
rect 2329 5185 2363 5219
rect 2973 5185 3007 5219
rect 3617 5185 3651 5219
rect 4269 5185 4303 5219
rect 4905 5185 4939 5219
rect 5549 5185 5583 5219
rect 6745 5185 6779 5219
rect 7205 5185 7239 5219
rect 7849 5185 7883 5219
rect 8769 5185 8803 5219
rect 9597 5185 9631 5219
rect 33793 5185 33827 5219
rect 6561 5049 6595 5083
rect 7941 5049 7975 5083
rect 1777 4981 1811 5015
rect 5641 4981 5675 5015
rect 7297 4981 7331 5015
rect 9413 4981 9447 5015
rect 33609 4981 33643 5015
rect 2697 4777 2731 4811
rect 3341 4777 3375 4811
rect 5641 4777 5675 4811
rect 6929 4777 6963 4811
rect 10057 4777 10091 4811
rect 1961 4709 1995 4743
rect 6285 4709 6319 4743
rect 4261 4641 4295 4675
rect 1869 4573 1903 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 4169 4573 4203 4607
rect 4905 4573 4939 4607
rect 5549 4573 5583 4607
rect 6193 4573 6227 4607
rect 6837 4573 6871 4607
rect 9965 4573 9999 4607
rect 26249 4573 26283 4607
rect 38025 4573 38059 4607
rect 4997 4437 5031 4471
rect 26341 4437 26375 4471
rect 38209 4437 38243 4471
rect 2329 4233 2363 4267
rect 1777 4097 1811 4131
rect 2237 4097 2271 4131
rect 2881 4097 2915 4131
rect 3525 4097 3559 4131
rect 3617 4097 3651 4131
rect 4445 4097 4479 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 5825 4097 5859 4131
rect 2973 4029 3007 4063
rect 4537 4029 4571 4063
rect 5181 4029 5215 4063
rect 1593 3961 1627 3995
rect 1777 3689 1811 3723
rect 3341 3689 3375 3723
rect 5733 3689 5767 3723
rect 6377 3689 6411 3723
rect 38117 3689 38151 3723
rect 4077 3621 4111 3655
rect 1685 3485 1719 3519
rect 2329 3485 2363 3519
rect 3249 3485 3283 3519
rect 3985 3485 4019 3519
rect 5089 3485 5123 3519
rect 5917 3485 5951 3519
rect 6561 3485 6595 3519
rect 38301 3485 38335 3519
rect 2605 3417 2639 3451
rect 5181 3349 5215 3383
rect 5273 3145 5307 3179
rect 6561 3145 6595 3179
rect 36737 3145 36771 3179
rect 2973 3077 3007 3111
rect 1593 3009 1627 3043
rect 2697 3009 2731 3043
rect 3801 3009 3835 3043
rect 4261 3009 4295 3043
rect 5181 3009 5215 3043
rect 6745 3009 6779 3043
rect 10057 3009 10091 3043
rect 28181 3009 28215 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 3617 2873 3651 2907
rect 1777 2805 1811 2839
rect 4353 2805 4387 2839
rect 9873 2805 9907 2839
rect 27997 2805 28031 2839
rect 38209 2805 38243 2839
rect 3985 2601 4019 2635
rect 4629 2601 4663 2635
rect 7297 2601 7331 2635
rect 11713 2601 11747 2635
rect 14289 2601 14323 2635
rect 14933 2601 14967 2635
rect 16865 2601 16899 2635
rect 22017 2601 22051 2635
rect 22661 2601 22695 2635
rect 29745 2601 29779 2635
rect 33609 2601 33643 2635
rect 36185 2601 36219 2635
rect 5273 2533 5307 2567
rect 30389 2533 30423 2567
rect 27445 2465 27479 2499
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 2789 2397 2823 2431
rect 4169 2397 4203 2431
rect 4813 2397 4847 2431
rect 5457 2397 5491 2431
rect 6561 2397 6595 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 11897 2397 11931 2431
rect 14473 2397 14507 2431
rect 15117 2397 15151 2431
rect 17049 2397 17083 2431
rect 18153 2397 18187 2431
rect 19441 2397 19475 2431
rect 22201 2397 22235 2431
rect 22845 2397 22879 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 29929 2397 29963 2431
rect 30573 2397 30607 2431
rect 32321 2397 32355 2431
rect 33793 2397 33827 2431
rect 35081 2397 35115 2431
rect 36369 2397 36403 2431
rect 38025 2397 38059 2431
rect 27261 2329 27295 2363
rect 1777 2261 1811 2295
rect 6745 2261 6779 2295
rect 9321 2261 9355 2295
rect 10609 2261 10643 2295
rect 18337 2261 18371 2295
rect 19625 2261 19659 2295
rect 24777 2261 24811 2295
rect 26065 2261 26099 2295
rect 32505 2261 32539 2295
rect 34897 2261 34931 2295
rect 38209 2261 38243 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 2501 37247 2559 37253
rect 2501 37213 2513 37247
rect 2547 37244 2559 37247
rect 2774 37244 2780 37256
rect 2547 37216 2780 37244
rect 2547 37213 2559 37216
rect 2501 37207 2559 37213
rect 2774 37204 2780 37216
rect 2832 37204 2838 37256
rect 3142 37244 3148 37256
rect 3103 37216 3148 37244
rect 3142 37204 3148 37216
rect 3200 37204 3206 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 4157 37247 4215 37253
rect 4157 37244 4169 37247
rect 3292 37216 4169 37244
rect 3292 37204 3298 37216
rect 4157 37213 4169 37216
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 4801 37247 4859 37253
rect 4801 37244 4813 37247
rect 4672 37216 4813 37244
rect 4672 37204 4678 37216
rect 4801 37213 4813 37216
rect 4847 37213 4859 37247
rect 6546 37244 6552 37256
rect 6507 37216 6552 37244
rect 4801 37207 4859 37213
rect 6546 37204 6552 37216
rect 6604 37204 6610 37256
rect 7834 37244 7840 37256
rect 7795 37216 7840 37244
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 9030 37204 9036 37256
rect 9088 37244 9094 37256
rect 9309 37247 9367 37253
rect 9309 37244 9321 37247
rect 9088 37216 9321 37244
rect 9088 37204 9094 37216
rect 9309 37213 9321 37216
rect 9355 37213 9367 37247
rect 9309 37207 9367 37213
rect 10413 37247 10471 37253
rect 10413 37213 10425 37247
rect 10459 37244 10471 37247
rect 11606 37244 11612 37256
rect 10459 37216 11612 37244
rect 10459 37213 10471 37216
rect 10413 37207 10471 37213
rect 11606 37204 11612 37216
rect 11664 37204 11670 37256
rect 12345 37247 12403 37253
rect 12345 37213 12357 37247
rect 12391 37213 12403 37247
rect 12345 37207 12403 37213
rect 5626 37176 5632 37188
rect 2976 37148 5632 37176
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 1765 37111 1823 37117
rect 1765 37108 1777 37111
rect 1360 37080 1777 37108
rect 1360 37068 1366 37080
rect 1765 37077 1777 37080
rect 1811 37077 1823 37111
rect 2314 37108 2320 37120
rect 2275 37080 2320 37108
rect 1765 37071 1823 37077
rect 2314 37068 2320 37080
rect 2372 37068 2378 37120
rect 2976 37117 3004 37148
rect 5626 37136 5632 37148
rect 5684 37136 5690 37188
rect 12360 37176 12388 37207
rect 13538 37204 13544 37256
rect 13596 37244 13602 37256
rect 14461 37247 14519 37253
rect 14461 37244 14473 37247
rect 13596 37216 14473 37244
rect 13596 37204 13602 37216
rect 14461 37213 14473 37216
rect 14507 37213 14519 37247
rect 15562 37244 15568 37256
rect 15523 37216 15568 37244
rect 14461 37207 14519 37213
rect 15562 37204 15568 37216
rect 15620 37204 15626 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18506 37204 18512 37256
rect 18564 37244 18570 37256
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 18564 37216 20085 37244
rect 18564 37204 18570 37216
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 20073 37207 20131 37213
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 20680 37216 22017 37244
rect 20680 37204 20686 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22925 37247 22983 37253
rect 22925 37244 22937 37247
rect 22612 37216 22937 37244
rect 22612 37204 22618 37216
rect 22925 37213 22937 37216
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 24544 37216 24777 37244
rect 24544 37204 24550 37216
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 25774 37204 25780 37256
rect 25832 37244 25838 37256
rect 26053 37247 26111 37253
rect 26053 37244 26065 37247
rect 25832 37216 26065 37244
rect 25832 37204 25838 37216
rect 26053 37213 26065 37216
rect 26099 37213 26111 37247
rect 27798 37244 27804 37256
rect 27759 37216 27804 37244
rect 26053 37207 26111 37213
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 27890 37204 27896 37256
rect 27948 37244 27954 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 27948 37216 29745 37244
rect 27948 37204 27954 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 30653 37247 30711 37253
rect 30653 37244 30665 37247
rect 30432 37216 30665 37244
rect 30432 37204 30438 37216
rect 30653 37213 30665 37216
rect 30699 37213 30711 37247
rect 30653 37207 30711 37213
rect 32214 37204 32220 37256
rect 32272 37244 32278 37256
rect 32493 37247 32551 37253
rect 32493 37244 32505 37247
rect 32272 37216 32505 37244
rect 32272 37204 32278 37216
rect 32493 37213 32505 37216
rect 32539 37213 32551 37247
rect 32493 37207 32551 37213
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 34882 37244 34888 37256
rect 34843 37216 34888 37244
rect 33781 37207 33839 37213
rect 34882 37204 34888 37216
rect 34940 37204 34946 37256
rect 36906 37244 36912 37256
rect 36867 37216 36912 37244
rect 36906 37204 36912 37216
rect 36964 37204 36970 37256
rect 37458 37244 37464 37256
rect 37419 37216 37464 37244
rect 37458 37204 37464 37216
rect 37516 37204 37522 37256
rect 14642 37176 14648 37188
rect 12360 37148 14648 37176
rect 14642 37136 14648 37148
rect 14700 37136 14706 37188
rect 15838 37136 15844 37188
rect 15896 37176 15902 37188
rect 15896 37148 18184 37176
rect 15896 37136 15902 37148
rect 2961 37111 3019 37117
rect 2961 37077 2973 37111
rect 3007 37077 3019 37111
rect 3970 37108 3976 37120
rect 3931 37080 3976 37108
rect 2961 37071 3019 37077
rect 3970 37068 3976 37080
rect 4028 37068 4034 37120
rect 4614 37108 4620 37120
rect 4575 37080 4620 37108
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 5810 37068 5816 37120
rect 5868 37108 5874 37120
rect 6733 37111 6791 37117
rect 6733 37108 6745 37111
rect 5868 37080 6745 37108
rect 5868 37068 5874 37080
rect 6733 37077 6745 37080
rect 6779 37077 6791 37111
rect 6733 37071 6791 37077
rect 7742 37068 7748 37120
rect 7800 37108 7806 37120
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7800 37080 8033 37108
rect 7800 37068 7806 37080
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 9122 37108 9128 37120
rect 9083 37080 9128 37108
rect 8021 37071 8079 37077
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10376 37080 10609 37108
rect 10376 37068 10382 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 10597 37071 10655 37077
rect 12434 37068 12440 37120
rect 12492 37108 12498 37120
rect 12529 37111 12587 37117
rect 12529 37108 12541 37111
rect 12492 37080 12541 37108
rect 12492 37068 12498 37080
rect 12529 37077 12541 37080
rect 12575 37077 12587 37111
rect 14274 37108 14280 37120
rect 14235 37080 14280 37108
rect 12529 37071 12587 37077
rect 14274 37068 14280 37080
rect 14332 37068 14338 37120
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 15749 37111 15807 37117
rect 15749 37108 15761 37111
rect 15528 37080 15761 37108
rect 15528 37068 15534 37080
rect 15749 37077 15761 37080
rect 15795 37077 15807 37111
rect 15749 37071 15807 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 18156 37117 18184 37148
rect 20898 37136 20904 37188
rect 20956 37176 20962 37188
rect 20956 37148 22784 37176
rect 20956 37136 20962 37148
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 18141 37111 18199 37117
rect 18141 37077 18153 37111
rect 18187 37077 18199 37111
rect 18141 37071 18199 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 22756 37117 22784 37148
rect 28074 37136 28080 37188
rect 28132 37176 28138 37188
rect 28132 37148 33640 37176
rect 28132 37136 28138 37148
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 22741 37111 22799 37117
rect 22741 37077 22753 37111
rect 22787 37077 22799 37111
rect 22741 37071 22799 37077
rect 23014 37068 23020 37120
rect 23072 37108 23078 37120
rect 24581 37111 24639 37117
rect 24581 37108 24593 37111
rect 23072 37080 24593 37108
rect 23072 37068 23078 37080
rect 24581 37077 24593 37080
rect 24627 37077 24639 37111
rect 24581 37071 24639 37077
rect 25038 37068 25044 37120
rect 25096 37108 25102 37120
rect 25869 37111 25927 37117
rect 25869 37108 25881 37111
rect 25096 37080 25881 37108
rect 25096 37068 25102 37080
rect 25869 37077 25881 37080
rect 25915 37077 25927 37111
rect 25869 37071 25927 37077
rect 27706 37068 27712 37120
rect 27764 37108 27770 37120
rect 27985 37111 28043 37117
rect 27985 37108 27997 37111
rect 27764 37080 27997 37108
rect 27764 37068 27770 37080
rect 27985 37077 27997 37080
rect 28031 37077 28043 37111
rect 27985 37071 28043 37077
rect 28994 37068 29000 37120
rect 29052 37108 29058 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29052 37080 29929 37108
rect 29052 37068 29058 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 30006 37068 30012 37120
rect 30064 37108 30070 37120
rect 30469 37111 30527 37117
rect 30469 37108 30481 37111
rect 30064 37080 30481 37108
rect 30064 37068 30070 37080
rect 30469 37077 30481 37080
rect 30515 37077 30527 37111
rect 30469 37071 30527 37077
rect 30650 37068 30656 37120
rect 30708 37108 30714 37120
rect 33612 37117 33640 37148
rect 34422 37136 34428 37188
rect 34480 37176 34486 37188
rect 34480 37148 35894 37176
rect 34480 37136 34486 37148
rect 32309 37111 32367 37117
rect 32309 37108 32321 37111
rect 30708 37080 32321 37108
rect 30708 37068 30714 37080
rect 32309 37077 32321 37080
rect 32355 37077 32367 37111
rect 32309 37071 32367 37077
rect 33597 37111 33655 37117
rect 33597 37077 33609 37111
rect 33643 37077 33655 37111
rect 33597 37071 33655 37077
rect 34790 37068 34796 37120
rect 34848 37108 34854 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34848 37080 35081 37108
rect 34848 37068 34854 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35866 37108 35894 37148
rect 36725 37111 36783 37117
rect 36725 37108 36737 37111
rect 35866 37080 36737 37108
rect 35069 37071 35127 37077
rect 36725 37077 36737 37080
rect 36771 37077 36783 37111
rect 36725 37071 36783 37077
rect 36814 37068 36820 37120
rect 36872 37108 36878 37120
rect 37645 37111 37703 37117
rect 37645 37108 37657 37111
rect 36872 37080 37657 37108
rect 36872 37068 36878 37080
rect 37645 37077 37657 37080
rect 37691 37077 37703 37111
rect 37645 37071 37703 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 14 36864 20 36916
rect 72 36904 78 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 72 36876 1777 36904
rect 72 36864 78 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 3513 36907 3571 36913
rect 3513 36873 3525 36907
rect 3559 36873 3571 36907
rect 3513 36867 3571 36873
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 3528 36768 3556 36867
rect 3970 36864 3976 36916
rect 4028 36904 4034 36916
rect 10226 36904 10232 36916
rect 4028 36876 10232 36904
rect 4028 36864 4034 36876
rect 10226 36864 10232 36876
rect 10284 36864 10290 36916
rect 25317 36907 25375 36913
rect 25317 36873 25329 36907
rect 25363 36904 25375 36907
rect 27798 36904 27804 36916
rect 25363 36876 27804 36904
rect 25363 36873 25375 36876
rect 25317 36867 25375 36873
rect 27798 36864 27804 36876
rect 27856 36864 27862 36916
rect 31481 36907 31539 36913
rect 31481 36873 31493 36907
rect 31527 36904 31539 36907
rect 34882 36904 34888 36916
rect 31527 36876 34888 36904
rect 31527 36873 31539 36876
rect 31481 36867 31539 36873
rect 34882 36864 34888 36876
rect 34940 36864 34946 36916
rect 35989 36907 36047 36913
rect 35989 36873 36001 36907
rect 36035 36873 36047 36907
rect 35989 36867 36047 36873
rect 38197 36907 38255 36913
rect 38197 36873 38209 36907
rect 38243 36904 38255 36907
rect 39298 36904 39304 36916
rect 38243 36876 39304 36904
rect 38243 36873 38255 36876
rect 38197 36867 38255 36873
rect 9122 36796 9128 36848
rect 9180 36836 9186 36848
rect 13814 36836 13820 36848
rect 9180 36808 13820 36836
rect 9180 36796 9186 36808
rect 13814 36796 13820 36808
rect 13872 36796 13878 36848
rect 36004 36836 36032 36867
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 36004 36808 38056 36836
rect 1627 36740 3556 36768
rect 3697 36771 3755 36777
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 3697 36737 3709 36771
rect 3743 36768 3755 36771
rect 3970 36768 3976 36780
rect 3743 36740 3976 36768
rect 3743 36737 3755 36740
rect 3697 36731 3755 36737
rect 3970 36728 3976 36740
rect 4028 36728 4034 36780
rect 4893 36771 4951 36777
rect 4893 36737 4905 36771
rect 4939 36768 4951 36771
rect 8294 36768 8300 36780
rect 4939 36740 8300 36768
rect 4939 36737 4951 36740
rect 4893 36731 4951 36737
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 25498 36768 25504 36780
rect 25459 36740 25504 36768
rect 25498 36728 25504 36740
rect 25556 36728 25562 36780
rect 29822 36728 29828 36780
rect 29880 36768 29886 36780
rect 31665 36771 31723 36777
rect 31665 36768 31677 36771
rect 29880 36740 31677 36768
rect 29880 36728 29886 36740
rect 31665 36737 31677 36740
rect 31711 36737 31723 36771
rect 31665 36731 31723 36737
rect 31754 36728 31760 36780
rect 31812 36768 31818 36780
rect 33137 36771 33195 36777
rect 33137 36768 33149 36771
rect 31812 36740 33149 36768
rect 31812 36728 31818 36740
rect 33137 36737 33149 36740
rect 33183 36737 33195 36771
rect 36170 36768 36176 36780
rect 36131 36740 36176 36768
rect 33137 36731 33195 36737
rect 36170 36728 36176 36740
rect 36228 36728 36234 36780
rect 36909 36771 36967 36777
rect 36909 36737 36921 36771
rect 36955 36768 36967 36771
rect 36998 36768 37004 36780
rect 36955 36740 37004 36768
rect 36955 36737 36967 36740
rect 36909 36731 36967 36737
rect 36998 36728 37004 36740
rect 37056 36728 37062 36780
rect 38028 36777 38056 36808
rect 38013 36771 38071 36777
rect 38013 36737 38025 36771
rect 38059 36737 38071 36771
rect 38013 36731 38071 36737
rect 2314 36660 2320 36712
rect 2372 36700 2378 36712
rect 8846 36700 8852 36712
rect 2372 36672 8852 36700
rect 2372 36660 2378 36672
rect 8846 36660 8852 36672
rect 8904 36660 8910 36712
rect 1578 36592 1584 36644
rect 1636 36632 1642 36644
rect 4709 36635 4767 36641
rect 4709 36632 4721 36635
rect 1636 36604 4721 36632
rect 1636 36592 1642 36604
rect 4709 36601 4721 36604
rect 4755 36601 4767 36635
rect 4709 36595 4767 36601
rect 32953 36635 33011 36641
rect 32953 36601 32965 36635
rect 32999 36632 33011 36635
rect 37458 36632 37464 36644
rect 32999 36604 37464 36632
rect 32999 36601 33011 36604
rect 32953 36595 33011 36601
rect 37458 36592 37464 36604
rect 37516 36592 37522 36644
rect 36722 36564 36728 36576
rect 36683 36536 36728 36564
rect 36722 36524 36728 36536
rect 36780 36524 36786 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 3970 36360 3976 36372
rect 3931 36332 3976 36360
rect 3970 36320 3976 36332
rect 4028 36320 4034 36372
rect 11606 36360 11612 36372
rect 11567 36332 11612 36360
rect 11606 36320 11612 36332
rect 11664 36320 11670 36372
rect 29822 36360 29828 36372
rect 29783 36332 29828 36360
rect 29822 36320 29828 36332
rect 29880 36320 29886 36372
rect 34977 36363 35035 36369
rect 34977 36329 34989 36363
rect 35023 36360 35035 36363
rect 36170 36360 36176 36372
rect 35023 36332 36176 36360
rect 35023 36329 35035 36332
rect 34977 36323 35035 36329
rect 36170 36320 36176 36332
rect 36228 36320 36234 36372
rect 4062 36156 4068 36168
rect 4023 36128 4068 36156
rect 4062 36116 4068 36128
rect 4120 36116 4126 36168
rect 11790 36156 11796 36168
rect 11751 36128 11796 36156
rect 11790 36116 11796 36128
rect 11848 36116 11854 36168
rect 29730 36156 29736 36168
rect 29691 36128 29736 36156
rect 29730 36116 29736 36128
rect 29788 36116 29794 36168
rect 34790 36116 34796 36168
rect 34848 36156 34854 36168
rect 34885 36159 34943 36165
rect 34885 36156 34897 36159
rect 34848 36128 34897 36156
rect 34848 36116 34854 36128
rect 34885 36125 34897 36128
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 38010 36116 38016 36168
rect 38068 36156 38074 36168
rect 38289 36159 38347 36165
rect 38289 36156 38301 36159
rect 38068 36128 38301 36156
rect 38068 36116 38074 36128
rect 38289 36125 38301 36128
rect 38335 36125 38347 36159
rect 38289 36119 38347 36125
rect 37274 35980 37280 36032
rect 37332 36020 37338 36032
rect 38105 36023 38163 36029
rect 38105 36020 38117 36023
rect 37332 35992 38117 36020
rect 37332 35980 37338 35992
rect 38105 35989 38117 35992
rect 38151 35989 38163 36023
rect 38105 35983 38163 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 24489 35819 24547 35825
rect 24489 35785 24501 35819
rect 24535 35816 24547 35819
rect 25498 35816 25504 35828
rect 24535 35788 25504 35816
rect 24535 35785 24547 35788
rect 24489 35779 24547 35785
rect 25498 35776 25504 35788
rect 25556 35776 25562 35828
rect 21910 35640 21916 35692
rect 21968 35680 21974 35692
rect 24397 35683 24455 35689
rect 24397 35680 24409 35683
rect 21968 35652 24409 35680
rect 21968 35640 21974 35652
rect 24397 35649 24409 35652
rect 24443 35649 24455 35683
rect 24397 35643 24455 35649
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 8294 35272 8300 35284
rect 8255 35244 8300 35272
rect 8294 35232 8300 35244
rect 8352 35232 8358 35284
rect 15473 35275 15531 35281
rect 15473 35241 15485 35275
rect 15519 35272 15531 35275
rect 16850 35272 16856 35284
rect 15519 35244 16856 35272
rect 15519 35241 15531 35244
rect 15473 35235 15531 35241
rect 16850 35232 16856 35244
rect 16908 35232 16914 35284
rect 8202 35068 8208 35080
rect 8163 35040 8208 35068
rect 8202 35028 8208 35040
rect 8260 35028 8266 35080
rect 14826 35028 14832 35080
rect 14884 35068 14890 35080
rect 15657 35071 15715 35077
rect 15657 35068 15669 35071
rect 14884 35040 15669 35068
rect 14884 35028 14890 35040
rect 15657 35037 15669 35040
rect 15703 35037 15715 35071
rect 15657 35031 15715 35037
rect 35342 35028 35348 35080
rect 35400 35068 35406 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 35400 35040 38025 35068
rect 35400 35028 35406 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 38194 34932 38200 34944
rect 38155 34904 38200 34932
rect 38194 34892 38200 34904
rect 38252 34892 38258 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 5537 34731 5595 34737
rect 5537 34697 5549 34731
rect 5583 34728 5595 34731
rect 6546 34728 6552 34740
rect 5583 34700 6552 34728
rect 5583 34697 5595 34700
rect 5537 34691 5595 34697
rect 6546 34688 6552 34700
rect 6604 34688 6610 34740
rect 6825 34731 6883 34737
rect 6825 34697 6837 34731
rect 6871 34728 6883 34731
rect 7834 34728 7840 34740
rect 6871 34700 7840 34728
rect 6871 34697 6883 34700
rect 6825 34691 6883 34697
rect 7834 34688 7840 34700
rect 7892 34688 7898 34740
rect 14642 34728 14648 34740
rect 14603 34700 14648 34728
rect 14642 34688 14648 34700
rect 14700 34688 14706 34740
rect 15289 34731 15347 34737
rect 15289 34697 15301 34731
rect 15335 34728 15347 34731
rect 15562 34728 15568 34740
rect 15335 34700 15568 34728
rect 15335 34697 15347 34700
rect 15289 34691 15347 34697
rect 15562 34688 15568 34700
rect 15620 34688 15626 34740
rect 17681 34731 17739 34737
rect 17681 34697 17693 34731
rect 17727 34728 17739 34731
rect 18506 34728 18512 34740
rect 17727 34700 18512 34728
rect 17727 34697 17739 34700
rect 17681 34691 17739 34697
rect 18506 34688 18512 34700
rect 18564 34688 18570 34740
rect 18785 34731 18843 34737
rect 18785 34697 18797 34731
rect 18831 34728 18843 34731
rect 20622 34728 20628 34740
rect 18831 34700 20628 34728
rect 18831 34697 18843 34700
rect 18785 34691 18843 34697
rect 20622 34688 20628 34700
rect 20680 34688 20686 34740
rect 27433 34731 27491 34737
rect 27433 34697 27445 34731
rect 27479 34728 27491 34731
rect 27890 34728 27896 34740
rect 27479 34700 27896 34728
rect 27479 34697 27491 34700
rect 27433 34691 27491 34697
rect 27890 34688 27896 34700
rect 27948 34688 27954 34740
rect 5721 34595 5779 34601
rect 5721 34561 5733 34595
rect 5767 34592 5779 34595
rect 5810 34592 5816 34604
rect 5767 34564 5816 34592
rect 5767 34561 5779 34564
rect 5721 34555 5779 34561
rect 5810 34552 5816 34564
rect 5868 34552 5874 34604
rect 6546 34552 6552 34604
rect 6604 34592 6610 34604
rect 7009 34595 7067 34601
rect 7009 34592 7021 34595
rect 6604 34564 7021 34592
rect 6604 34552 6610 34564
rect 7009 34561 7021 34564
rect 7055 34561 7067 34595
rect 7009 34555 7067 34561
rect 14734 34552 14740 34604
rect 14792 34592 14798 34604
rect 14829 34595 14887 34601
rect 14829 34592 14841 34595
rect 14792 34564 14841 34592
rect 14792 34552 14798 34564
rect 14829 34561 14841 34564
rect 14875 34561 14887 34595
rect 14829 34555 14887 34561
rect 15010 34552 15016 34604
rect 15068 34592 15074 34604
rect 15473 34595 15531 34601
rect 15473 34592 15485 34595
rect 15068 34564 15485 34592
rect 15068 34552 15074 34564
rect 15473 34561 15485 34564
rect 15519 34561 15531 34595
rect 17862 34592 17868 34604
rect 17823 34564 17868 34592
rect 15473 34555 15531 34561
rect 17862 34552 17868 34564
rect 17920 34552 17926 34604
rect 18969 34595 19027 34601
rect 18969 34561 18981 34595
rect 19015 34561 19027 34595
rect 18969 34555 19027 34561
rect 17494 34484 17500 34536
rect 17552 34524 17558 34536
rect 18984 34524 19012 34555
rect 27246 34552 27252 34604
rect 27304 34592 27310 34604
rect 27617 34595 27675 34601
rect 27617 34592 27629 34595
rect 27304 34564 27629 34592
rect 27304 34552 27310 34564
rect 27617 34561 27629 34564
rect 27663 34561 27675 34595
rect 27617 34555 27675 34561
rect 17552 34496 19012 34524
rect 17552 34484 17558 34496
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 14550 34076 14556 34128
rect 14608 34116 14614 34128
rect 15841 34119 15899 34125
rect 15841 34116 15853 34119
rect 14608 34088 15853 34116
rect 14608 34076 14614 34088
rect 15841 34085 15853 34088
rect 15887 34085 15899 34119
rect 15841 34079 15899 34085
rect 4614 33940 4620 33992
rect 4672 33980 4678 33992
rect 9125 33983 9183 33989
rect 9125 33980 9137 33983
rect 4672 33952 9137 33980
rect 4672 33940 4678 33952
rect 9125 33949 9137 33952
rect 9171 33949 9183 33983
rect 14274 33980 14280 33992
rect 14235 33952 14280 33980
rect 9125 33943 9183 33949
rect 14274 33940 14280 33952
rect 14332 33940 14338 33992
rect 15749 33983 15807 33989
rect 15749 33949 15761 33983
rect 15795 33980 15807 33983
rect 15838 33980 15844 33992
rect 15795 33952 15844 33980
rect 15795 33949 15807 33952
rect 15749 33943 15807 33949
rect 15838 33940 15844 33952
rect 15896 33940 15902 33992
rect 23014 33980 23020 33992
rect 22975 33952 23020 33980
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 25038 33980 25044 33992
rect 24999 33952 25044 33980
rect 25038 33940 25044 33952
rect 25096 33940 25102 33992
rect 27985 33983 28043 33989
rect 27985 33949 27997 33983
rect 28031 33980 28043 33983
rect 28074 33980 28080 33992
rect 28031 33952 28080 33980
rect 28031 33949 28043 33952
rect 27985 33943 28043 33949
rect 28074 33940 28080 33952
rect 28132 33940 28138 33992
rect 9217 33847 9275 33853
rect 9217 33813 9229 33847
rect 9263 33844 9275 33847
rect 11882 33844 11888 33856
rect 9263 33816 11888 33844
rect 9263 33813 9275 33816
rect 9217 33807 9275 33813
rect 11882 33804 11888 33816
rect 11940 33804 11946 33856
rect 14369 33847 14427 33853
rect 14369 33813 14381 33847
rect 14415 33844 14427 33847
rect 15102 33844 15108 33856
rect 14415 33816 15108 33844
rect 14415 33813 14427 33816
rect 14369 33807 14427 33813
rect 15102 33804 15108 33816
rect 15160 33804 15166 33856
rect 20162 33804 20168 33856
rect 20220 33844 20226 33856
rect 23109 33847 23167 33853
rect 23109 33844 23121 33847
rect 20220 33816 23121 33844
rect 20220 33804 20226 33816
rect 23109 33813 23121 33816
rect 23155 33813 23167 33847
rect 25130 33844 25136 33856
rect 25091 33816 25136 33844
rect 23109 33807 23167 33813
rect 25130 33804 25136 33816
rect 25188 33804 25194 33856
rect 28074 33844 28080 33856
rect 28035 33816 28080 33844
rect 28074 33804 28080 33816
rect 28132 33804 28138 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1762 33504 1768 33516
rect 1723 33476 1768 33504
rect 1762 33464 1768 33476
rect 1820 33464 1826 33516
rect 38286 33504 38292 33516
rect 38247 33476 38292 33504
rect 38286 33464 38292 33476
rect 38344 33464 38350 33516
rect 1581 33303 1639 33309
rect 1581 33269 1593 33303
rect 1627 33300 1639 33303
rect 3878 33300 3884 33312
rect 1627 33272 3884 33300
rect 1627 33269 1639 33272
rect 1581 33263 1639 33269
rect 3878 33260 3884 33272
rect 3936 33260 3942 33312
rect 38102 33300 38108 33312
rect 38063 33272 38108 33300
rect 38102 33260 38108 33272
rect 38160 33260 38166 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 27617 33099 27675 33105
rect 27617 33065 27629 33099
rect 27663 33096 27675 33099
rect 31754 33096 31760 33108
rect 27663 33068 31760 33096
rect 27663 33065 27675 33068
rect 27617 33059 27675 33065
rect 31754 33056 31760 33068
rect 31812 33056 31818 33108
rect 5626 32892 5632 32904
rect 5587 32864 5632 32892
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 27522 32892 27528 32904
rect 27483 32864 27528 32892
rect 27522 32852 27528 32864
rect 27580 32852 27586 32904
rect 5718 32756 5724 32768
rect 5679 32728 5724 32756
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1762 32416 1768 32428
rect 1723 32388 1768 32416
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 35434 32376 35440 32428
rect 35492 32416 35498 32428
rect 38013 32419 38071 32425
rect 38013 32416 38025 32419
rect 35492 32388 38025 32416
rect 35492 32376 35498 32388
rect 38013 32385 38025 32388
rect 38059 32385 38071 32419
rect 38013 32379 38071 32385
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 3970 32212 3976 32224
rect 1627 32184 3976 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 3970 32172 3976 32184
rect 4028 32172 4034 32224
rect 38194 32212 38200 32224
rect 38155 32184 38200 32212
rect 38194 32172 38200 32184
rect 38252 32172 38258 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 6546 32008 6552 32020
rect 6507 31980 6552 32008
rect 6546 31968 6552 31980
rect 6604 31968 6610 32020
rect 11790 31968 11796 32020
rect 11848 32008 11854 32020
rect 12161 32011 12219 32017
rect 12161 32008 12173 32011
rect 11848 31980 12173 32008
rect 11848 31968 11854 31980
rect 12161 31977 12173 31980
rect 12207 31977 12219 32011
rect 12161 31971 12219 31977
rect 16298 31832 16304 31884
rect 16356 31872 16362 31884
rect 20993 31875 21051 31881
rect 20993 31872 21005 31875
rect 16356 31844 21005 31872
rect 16356 31832 16362 31844
rect 20993 31841 21005 31844
rect 21039 31841 21051 31875
rect 34422 31872 34428 31884
rect 20993 31835 21051 31841
rect 33612 31844 34428 31872
rect 6457 31807 6515 31813
rect 6457 31773 6469 31807
rect 6503 31804 6515 31807
rect 7374 31804 7380 31816
rect 6503 31776 7380 31804
rect 6503 31773 6515 31776
rect 6457 31767 6515 31773
rect 7374 31764 7380 31776
rect 7432 31764 7438 31816
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31804 12127 31807
rect 12894 31804 12900 31816
rect 12115 31776 12900 31804
rect 12115 31773 12127 31776
rect 12069 31767 12127 31773
rect 12894 31764 12900 31776
rect 12952 31764 12958 31816
rect 20898 31804 20904 31816
rect 20859 31776 20904 31804
rect 20898 31764 20904 31776
rect 20956 31764 20962 31816
rect 33612 31813 33640 31844
rect 34422 31832 34428 31844
rect 34480 31832 34486 31884
rect 33597 31807 33655 31813
rect 33597 31773 33609 31807
rect 33643 31773 33655 31807
rect 33597 31767 33655 31773
rect 33686 31764 33692 31816
rect 33744 31804 33750 31816
rect 33744 31776 33789 31804
rect 33744 31764 33750 31776
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 10226 31328 10232 31340
rect 10187 31300 10232 31328
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 13814 31328 13820 31340
rect 13775 31300 13820 31328
rect 13814 31288 13820 31300
rect 13872 31288 13878 31340
rect 27157 31331 27215 31337
rect 27157 31297 27169 31331
rect 27203 31328 27215 31331
rect 30650 31328 30656 31340
rect 27203 31300 30656 31328
rect 27203 31297 27215 31300
rect 27157 31291 27215 31297
rect 30650 31288 30656 31300
rect 30708 31288 30714 31340
rect 10321 31127 10379 31133
rect 10321 31093 10333 31127
rect 10367 31124 10379 31127
rect 11514 31124 11520 31136
rect 10367 31096 11520 31124
rect 10367 31093 10379 31096
rect 10321 31087 10379 31093
rect 11514 31084 11520 31096
rect 11572 31084 11578 31136
rect 13909 31127 13967 31133
rect 13909 31093 13921 31127
rect 13955 31124 13967 31127
rect 16206 31124 16212 31136
rect 13955 31096 16212 31124
rect 13955 31093 13967 31096
rect 13909 31087 13967 31093
rect 16206 31084 16212 31096
rect 16264 31084 16270 31136
rect 24578 31084 24584 31136
rect 24636 31124 24642 31136
rect 27249 31127 27307 31133
rect 27249 31124 27261 31127
rect 24636 31096 27261 31124
rect 24636 31084 24642 31096
rect 27249 31093 27261 31096
rect 27295 31093 27307 31127
rect 27249 31087 27307 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 34885 30923 34943 30929
rect 34885 30889 34897 30923
rect 34931 30920 34943 30923
rect 35342 30920 35348 30932
rect 34931 30892 35348 30920
rect 34931 30889 34943 30892
rect 34885 30883 34943 30889
rect 35342 30880 35348 30892
rect 35400 30880 35406 30932
rect 37274 30784 37280 30796
rect 29748 30756 37280 30784
rect 1762 30716 1768 30728
rect 1723 30688 1768 30716
rect 1762 30676 1768 30688
rect 1820 30676 1826 30728
rect 29748 30725 29776 30756
rect 37274 30744 37280 30756
rect 37332 30744 37338 30796
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30716 24915 30719
rect 29733 30719 29791 30725
rect 24903 30688 26234 30716
rect 24903 30685 24915 30688
rect 24857 30679 24915 30685
rect 26206 30648 26234 30688
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 29914 30676 29920 30728
rect 29972 30716 29978 30728
rect 35069 30719 35127 30725
rect 35069 30716 35081 30719
rect 29972 30688 35081 30716
rect 29972 30676 29978 30688
rect 35069 30685 35081 30688
rect 35115 30685 35127 30719
rect 35069 30679 35127 30685
rect 30006 30648 30012 30660
rect 26206 30620 30012 30648
rect 30006 30608 30012 30620
rect 30064 30608 30070 30660
rect 1486 30540 1492 30592
rect 1544 30580 1550 30592
rect 1581 30583 1639 30589
rect 1581 30580 1593 30583
rect 1544 30552 1593 30580
rect 1544 30540 1550 30552
rect 1581 30549 1593 30552
rect 1627 30549 1639 30583
rect 24946 30580 24952 30592
rect 24907 30552 24952 30580
rect 1581 30543 1639 30549
rect 24946 30540 24952 30552
rect 25004 30540 25010 30592
rect 29822 30580 29828 30592
rect 29783 30552 29828 30580
rect 29822 30540 29828 30552
rect 29880 30540 29886 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 36722 30308 36728 30320
rect 29932 30280 36728 30308
rect 8846 30240 8852 30252
rect 8807 30212 8852 30240
rect 8846 30200 8852 30212
rect 8904 30200 8910 30252
rect 29932 30249 29960 30280
rect 36722 30268 36728 30280
rect 36780 30268 36786 30320
rect 29917 30243 29975 30249
rect 29917 30209 29929 30243
rect 29963 30209 29975 30243
rect 29917 30203 29975 30209
rect 33594 30200 33600 30252
rect 33652 30240 33658 30252
rect 38013 30243 38071 30249
rect 38013 30240 38025 30243
rect 33652 30212 38025 30240
rect 33652 30200 33658 30212
rect 38013 30209 38025 30212
rect 38059 30209 38071 30243
rect 38013 30203 38071 30209
rect 8941 30039 8999 30045
rect 8941 30005 8953 30039
rect 8987 30036 8999 30039
rect 12434 30036 12440 30048
rect 8987 30008 12440 30036
rect 8987 30005 8999 30008
rect 8941 29999 8999 30005
rect 12434 29996 12440 30008
rect 12492 29996 12498 30048
rect 30006 30036 30012 30048
rect 29967 30008 30012 30036
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 38194 30036 38200 30048
rect 38155 30008 38200 30036
rect 38194 29996 38200 30008
rect 38252 29996 38258 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 14826 29832 14832 29844
rect 14787 29804 14832 29832
rect 14826 29792 14832 29804
rect 14884 29792 14890 29844
rect 16945 29835 17003 29841
rect 16945 29801 16957 29835
rect 16991 29832 17003 29835
rect 17862 29832 17868 29844
rect 16991 29804 17868 29832
rect 16991 29801 17003 29804
rect 16945 29795 17003 29801
rect 17862 29792 17868 29804
rect 17920 29792 17926 29844
rect 34977 29835 35035 29841
rect 34977 29801 34989 29835
rect 35023 29832 35035 29835
rect 35434 29832 35440 29844
rect 35023 29804 35440 29832
rect 35023 29801 35035 29804
rect 34977 29795 35035 29801
rect 35434 29792 35440 29804
rect 35492 29792 35498 29844
rect 3878 29588 3884 29640
rect 3936 29628 3942 29640
rect 6181 29631 6239 29637
rect 6181 29628 6193 29631
rect 3936 29600 6193 29628
rect 3936 29588 3942 29600
rect 6181 29597 6193 29600
rect 6227 29597 6239 29631
rect 14734 29628 14740 29640
rect 14695 29600 14740 29628
rect 6181 29591 6239 29597
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 15838 29588 15844 29640
rect 15896 29628 15902 29640
rect 16853 29631 16911 29637
rect 16853 29628 16865 29631
rect 15896 29600 16865 29628
rect 15896 29588 15902 29600
rect 16853 29597 16865 29600
rect 16899 29597 16911 29631
rect 16853 29591 16911 29597
rect 33778 29588 33784 29640
rect 33836 29628 33842 29640
rect 35161 29631 35219 29637
rect 35161 29628 35173 29631
rect 33836 29600 35173 29628
rect 33836 29588 33842 29600
rect 35161 29597 35173 29600
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 6273 29495 6331 29501
rect 6273 29461 6285 29495
rect 6319 29492 6331 29495
rect 8110 29492 8116 29504
rect 6319 29464 8116 29492
rect 6319 29461 6331 29464
rect 6273 29455 6331 29461
rect 8110 29452 8116 29464
rect 8168 29452 8174 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 14185 29291 14243 29297
rect 14185 29257 14197 29291
rect 14231 29288 14243 29291
rect 15010 29288 15016 29300
rect 14231 29260 15016 29288
rect 14231 29257 14243 29260
rect 14185 29251 14243 29257
rect 15010 29248 15016 29260
rect 15068 29248 15074 29300
rect 17494 29288 17500 29300
rect 17455 29260 17500 29288
rect 17494 29248 17500 29260
rect 17552 29248 17558 29300
rect 27246 29288 27252 29300
rect 27207 29260 27252 29288
rect 27246 29248 27252 29260
rect 27304 29248 27310 29300
rect 1762 29152 1768 29164
rect 1723 29124 1768 29152
rect 1762 29112 1768 29124
rect 1820 29112 1826 29164
rect 14090 29152 14096 29164
rect 14051 29124 14096 29152
rect 14090 29112 14096 29124
rect 14148 29112 14154 29164
rect 15654 29112 15660 29164
rect 15712 29152 15718 29164
rect 17405 29155 17463 29161
rect 17405 29152 17417 29155
rect 15712 29124 17417 29152
rect 15712 29112 15718 29124
rect 17405 29121 17417 29124
rect 17451 29121 17463 29155
rect 17405 29115 17463 29121
rect 24486 29112 24492 29164
rect 24544 29152 24550 29164
rect 27157 29155 27215 29161
rect 27157 29152 27169 29155
rect 24544 29124 27169 29152
rect 24544 29112 24550 29124
rect 27157 29121 27169 29124
rect 27203 29121 27215 29155
rect 38286 29152 38292 29164
rect 38247 29124 38292 29152
rect 27157 29115 27215 29121
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 1581 29019 1639 29025
rect 1581 28985 1593 29019
rect 1627 29016 1639 29019
rect 6546 29016 6552 29028
rect 1627 28988 6552 29016
rect 1627 28985 1639 28988
rect 1581 28979 1639 28985
rect 6546 28976 6552 28988
rect 6604 28976 6610 29028
rect 33318 28976 33324 29028
rect 33376 29016 33382 29028
rect 38105 29019 38163 29025
rect 38105 29016 38117 29019
rect 33376 28988 38117 29016
rect 33376 28976 33382 28988
rect 38105 28985 38117 28988
rect 38151 28985 38163 29019
rect 38105 28979 38163 28985
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 5629 28747 5687 28753
rect 5629 28713 5641 28747
rect 5675 28744 5687 28747
rect 5810 28744 5816 28756
rect 5675 28716 5816 28744
rect 5675 28713 5687 28716
rect 5629 28707 5687 28713
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 17129 28747 17187 28753
rect 17129 28744 17141 28747
rect 14884 28716 17141 28744
rect 14884 28704 14890 28716
rect 17129 28713 17141 28716
rect 17175 28713 17187 28747
rect 17129 28707 17187 28713
rect 32861 28747 32919 28753
rect 32861 28713 32873 28747
rect 32907 28744 32919 28747
rect 33778 28744 33784 28756
rect 32907 28716 33784 28744
rect 32907 28713 32919 28716
rect 32861 28707 32919 28713
rect 33778 28704 33784 28716
rect 33836 28704 33842 28756
rect 5537 28543 5595 28549
rect 5537 28509 5549 28543
rect 5583 28540 5595 28543
rect 6178 28540 6184 28552
rect 5583 28512 6184 28540
rect 5583 28509 5595 28512
rect 5537 28503 5595 28509
rect 6178 28500 6184 28512
rect 6236 28500 6242 28552
rect 17037 28543 17095 28549
rect 17037 28509 17049 28543
rect 17083 28540 17095 28543
rect 18322 28540 18328 28552
rect 17083 28512 18328 28540
rect 17083 28509 17095 28512
rect 17037 28503 17095 28509
rect 18322 28500 18328 28512
rect 18380 28500 18386 28552
rect 32766 28540 32772 28552
rect 32727 28512 32772 28540
rect 32766 28500 32772 28512
rect 32824 28500 32830 28552
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3970 28024 3976 28076
rect 4028 28064 4034 28076
rect 4249 28067 4307 28073
rect 4249 28064 4261 28067
rect 4028 28036 4261 28064
rect 4028 28024 4034 28036
rect 4249 28033 4261 28036
rect 4295 28033 4307 28067
rect 4249 28027 4307 28033
rect 30377 28067 30435 28073
rect 30377 28033 30389 28067
rect 30423 28064 30435 28067
rect 38102 28064 38108 28076
rect 30423 28036 38108 28064
rect 30423 28033 30435 28036
rect 30377 28027 30435 28033
rect 38102 28024 38108 28036
rect 38160 28024 38166 28076
rect 4341 27863 4399 27869
rect 4341 27829 4353 27863
rect 4387 27860 4399 27863
rect 4798 27860 4804 27872
rect 4387 27832 4804 27860
rect 4387 27829 4399 27832
rect 4341 27823 4399 27829
rect 4798 27820 4804 27832
rect 4856 27820 4862 27872
rect 30466 27860 30472 27872
rect 30427 27832 30472 27860
rect 30466 27820 30472 27832
rect 30524 27820 30530 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1762 27452 1768 27464
rect 1723 27424 1768 27452
rect 1762 27412 1768 27424
rect 1820 27412 1826 27464
rect 20622 27412 20628 27464
rect 20680 27452 20686 27464
rect 20993 27455 21051 27461
rect 20993 27452 21005 27455
rect 20680 27424 21005 27452
rect 20680 27412 20686 27424
rect 20993 27421 21005 27424
rect 21039 27421 21051 27455
rect 20993 27415 21051 27421
rect 36722 27412 36728 27464
rect 36780 27452 36786 27464
rect 38013 27455 38071 27461
rect 38013 27452 38025 27455
rect 36780 27424 38025 27452
rect 36780 27412 36786 27424
rect 38013 27421 38025 27424
rect 38059 27421 38071 27455
rect 38013 27415 38071 27421
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 5718 27316 5724 27328
rect 1627 27288 5724 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 5718 27276 5724 27288
rect 5776 27276 5782 27328
rect 20809 27319 20867 27325
rect 20809 27285 20821 27319
rect 20855 27316 20867 27319
rect 20898 27316 20904 27328
rect 20855 27288 20904 27316
rect 20855 27285 20867 27288
rect 20809 27279 20867 27285
rect 20898 27276 20904 27288
rect 20956 27276 20962 27328
rect 38194 27316 38200 27328
rect 38155 27288 38200 27316
rect 38194 27276 38200 27288
rect 38252 27276 38258 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 29181 27115 29239 27121
rect 29181 27081 29193 27115
rect 29227 27112 29239 27115
rect 29914 27112 29920 27124
rect 29227 27084 29920 27112
rect 29227 27081 29239 27084
rect 29181 27075 29239 27081
rect 29914 27072 29920 27084
rect 29972 27072 29978 27124
rect 6546 26976 6552 26988
rect 6507 26948 6552 26976
rect 6546 26936 6552 26948
rect 6604 26936 6610 26988
rect 20898 26976 20904 26988
rect 20859 26948 20904 26976
rect 20898 26936 20904 26948
rect 20956 26936 20962 26988
rect 24210 26936 24216 26988
rect 24268 26976 24274 26988
rect 29089 26979 29147 26985
rect 29089 26976 29101 26979
rect 24268 26948 29101 26976
rect 24268 26936 24274 26948
rect 29089 26945 29101 26948
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 6641 26775 6699 26781
rect 6641 26741 6653 26775
rect 6687 26772 6699 26775
rect 8846 26772 8852 26784
rect 6687 26744 8852 26772
rect 6687 26741 6699 26744
rect 6641 26735 6699 26741
rect 8846 26732 8852 26744
rect 8904 26732 8910 26784
rect 20530 26732 20536 26784
rect 20588 26772 20594 26784
rect 20717 26775 20775 26781
rect 20717 26772 20729 26775
rect 20588 26744 20729 26772
rect 20588 26732 20594 26744
rect 20717 26741 20729 26744
rect 20763 26741 20775 26775
rect 20717 26735 20775 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 12713 26503 12771 26509
rect 12713 26469 12725 26503
rect 12759 26469 12771 26503
rect 12713 26463 12771 26469
rect 13357 26503 13415 26509
rect 13357 26469 13369 26503
rect 13403 26500 13415 26503
rect 14458 26500 14464 26512
rect 13403 26472 14464 26500
rect 13403 26469 13415 26472
rect 13357 26463 13415 26469
rect 12728 26432 12756 26463
rect 14458 26460 14464 26472
rect 14516 26460 14522 26512
rect 15933 26503 15991 26509
rect 15933 26469 15945 26503
rect 15979 26500 15991 26503
rect 17218 26500 17224 26512
rect 15979 26472 17224 26500
rect 15979 26469 15991 26472
rect 15933 26463 15991 26469
rect 17218 26460 17224 26472
rect 17276 26460 17282 26512
rect 12728 26404 13584 26432
rect 11790 26324 11796 26376
rect 11848 26364 11854 26376
rect 12253 26367 12311 26373
rect 12253 26364 12265 26367
rect 11848 26336 12265 26364
rect 11848 26324 11854 26336
rect 12253 26333 12265 26336
rect 12299 26364 12311 26367
rect 12299 26336 12434 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 12406 26296 12434 26336
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 13556 26373 13584 26404
rect 12897 26367 12955 26373
rect 12897 26364 12909 26367
rect 12584 26336 12909 26364
rect 12584 26324 12590 26336
rect 12897 26333 12909 26336
rect 12943 26333 12955 26367
rect 12897 26327 12955 26333
rect 13541 26367 13599 26373
rect 13541 26333 13553 26367
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 15286 26324 15292 26376
rect 15344 26364 15350 26376
rect 16117 26367 16175 26373
rect 16117 26364 16129 26367
rect 15344 26336 16129 26364
rect 15344 26324 15350 26336
rect 16117 26333 16129 26336
rect 16163 26333 16175 26367
rect 16117 26327 16175 26333
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26333 17279 26367
rect 17221 26327 17279 26333
rect 16850 26296 16856 26308
rect 12406 26268 16856 26296
rect 16850 26256 16856 26268
rect 16908 26296 16914 26308
rect 17236 26296 17264 26327
rect 20622 26324 20628 26376
rect 20680 26364 20686 26376
rect 20993 26367 21051 26373
rect 20993 26364 21005 26367
rect 20680 26336 21005 26364
rect 20680 26324 20686 26336
rect 20993 26333 21005 26336
rect 21039 26333 21051 26367
rect 20993 26327 21051 26333
rect 16908 26268 17264 26296
rect 16908 26256 16914 26268
rect 20438 26256 20444 26308
rect 20496 26296 20502 26308
rect 21085 26299 21143 26305
rect 21085 26296 21097 26299
rect 20496 26268 21097 26296
rect 20496 26256 20502 26268
rect 21085 26265 21097 26268
rect 21131 26265 21143 26299
rect 21085 26259 21143 26265
rect 11974 26188 11980 26240
rect 12032 26228 12038 26240
rect 12069 26231 12127 26237
rect 12069 26228 12081 26231
rect 12032 26200 12081 26228
rect 12032 26188 12038 26200
rect 12069 26197 12081 26200
rect 12115 26197 12127 26231
rect 12069 26191 12127 26197
rect 17037 26231 17095 26237
rect 17037 26197 17049 26231
rect 17083 26228 17095 26231
rect 17678 26228 17684 26240
rect 17083 26200 17684 26228
rect 17083 26197 17095 26200
rect 17037 26191 17095 26197
rect 17678 26188 17684 26200
rect 17736 26188 17742 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 33594 26024 33600 26036
rect 33555 25996 33600 26024
rect 33594 25984 33600 25996
rect 33652 25984 33658 26036
rect 36722 26024 36728 26036
rect 36683 25996 36728 26024
rect 36722 25984 36728 25996
rect 36780 25984 36786 26036
rect 12526 25916 12532 25968
rect 12584 25956 12590 25968
rect 12584 25928 14228 25956
rect 12584 25916 12590 25928
rect 5442 25848 5448 25900
rect 5500 25888 5506 25900
rect 10597 25891 10655 25897
rect 10597 25888 10609 25891
rect 5500 25860 10609 25888
rect 5500 25848 5506 25860
rect 10597 25857 10609 25860
rect 10643 25888 10655 25891
rect 11790 25888 11796 25900
rect 10643 25860 11796 25888
rect 10643 25857 10655 25860
rect 10597 25851 10655 25857
rect 11790 25848 11796 25860
rect 11848 25848 11854 25900
rect 11974 25888 11980 25900
rect 11935 25860 11980 25888
rect 11974 25848 11980 25860
rect 12032 25848 12038 25900
rect 12618 25888 12624 25900
rect 12579 25860 12624 25888
rect 12618 25848 12624 25860
rect 12676 25848 12682 25900
rect 14200 25897 14228 25928
rect 14185 25891 14243 25897
rect 14185 25857 14197 25891
rect 14231 25857 14243 25891
rect 15286 25888 15292 25900
rect 15247 25860 15292 25888
rect 14185 25851 14243 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 16850 25888 16856 25900
rect 16811 25860 16856 25888
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17678 25888 17684 25900
rect 17639 25860 17684 25888
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 23569 25891 23627 25897
rect 23569 25888 23581 25891
rect 23532 25860 23581 25888
rect 23532 25848 23538 25860
rect 23569 25857 23581 25860
rect 23615 25857 23627 25891
rect 23569 25851 23627 25857
rect 31754 25848 31760 25900
rect 31812 25888 31818 25900
rect 33781 25891 33839 25897
rect 33781 25888 33793 25891
rect 31812 25860 33793 25888
rect 31812 25848 31818 25860
rect 33781 25857 33793 25860
rect 33827 25857 33839 25891
rect 36906 25888 36912 25900
rect 36867 25860 36912 25888
rect 33781 25851 33839 25857
rect 36906 25848 36912 25860
rect 36964 25848 36970 25900
rect 13538 25820 13544 25832
rect 13499 25792 13544 25820
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 15930 25820 15936 25832
rect 15891 25792 15936 25820
rect 15930 25780 15936 25792
rect 15988 25780 15994 25832
rect 10594 25644 10600 25696
rect 10652 25684 10658 25696
rect 10689 25687 10747 25693
rect 10689 25684 10701 25687
rect 10652 25656 10701 25684
rect 10652 25644 10658 25656
rect 10689 25653 10701 25656
rect 10735 25653 10747 25687
rect 11790 25684 11796 25696
rect 11751 25656 11796 25684
rect 10689 25647 10747 25653
rect 11790 25644 11796 25656
rect 11848 25644 11854 25696
rect 12437 25687 12495 25693
rect 12437 25653 12449 25687
rect 12483 25684 12495 25687
rect 13998 25684 14004 25696
rect 12483 25656 14004 25684
rect 12483 25653 12495 25656
rect 12437 25647 12495 25653
rect 13998 25644 14004 25656
rect 14056 25644 14062 25696
rect 14274 25684 14280 25696
rect 14235 25656 14280 25684
rect 14274 25644 14280 25656
rect 14332 25644 14338 25696
rect 15194 25644 15200 25696
rect 15252 25684 15258 25696
rect 15381 25687 15439 25693
rect 15381 25684 15393 25687
rect 15252 25656 15393 25684
rect 15252 25644 15258 25656
rect 15381 25653 15393 25656
rect 15427 25653 15439 25687
rect 16942 25684 16948 25696
rect 16903 25656 16948 25684
rect 15381 25647 15439 25653
rect 16942 25644 16948 25656
rect 17000 25644 17006 25696
rect 17494 25684 17500 25696
rect 17455 25656 17500 25684
rect 17494 25644 17500 25656
rect 17552 25644 17558 25696
rect 23385 25687 23443 25693
rect 23385 25653 23397 25687
rect 23431 25684 23443 25687
rect 23566 25684 23572 25696
rect 23431 25656 23572 25684
rect 23431 25653 23443 25656
rect 23385 25647 23443 25653
rect 23566 25644 23572 25656
rect 23624 25644 23630 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 9769 25483 9827 25489
rect 9769 25449 9781 25483
rect 9815 25480 9827 25483
rect 12618 25480 12624 25492
rect 9815 25452 12624 25480
rect 9815 25449 9827 25452
rect 9769 25443 9827 25449
rect 12618 25440 12624 25452
rect 12676 25440 12682 25492
rect 14734 25480 14740 25492
rect 14695 25452 14740 25480
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 1581 25415 1639 25421
rect 1581 25381 1593 25415
rect 1627 25412 1639 25415
rect 5810 25412 5816 25424
rect 1627 25384 5816 25412
rect 1627 25381 1639 25384
rect 1581 25375 1639 25381
rect 5810 25372 5816 25384
rect 5868 25372 5874 25424
rect 11057 25415 11115 25421
rect 11057 25381 11069 25415
rect 11103 25412 11115 25415
rect 13354 25412 13360 25424
rect 11103 25384 13360 25412
rect 11103 25381 11115 25384
rect 11057 25375 11115 25381
rect 13354 25372 13360 25384
rect 13412 25372 13418 25424
rect 8110 25304 8116 25356
rect 8168 25344 8174 25356
rect 10413 25347 10471 25353
rect 10413 25344 10425 25347
rect 8168 25316 10425 25344
rect 8168 25304 8174 25316
rect 10413 25313 10425 25316
rect 10459 25313 10471 25347
rect 10594 25344 10600 25356
rect 10555 25316 10600 25344
rect 10413 25307 10471 25313
rect 10594 25304 10600 25316
rect 10652 25304 10658 25356
rect 11790 25304 11796 25356
rect 11848 25344 11854 25356
rect 12713 25347 12771 25353
rect 12713 25344 12725 25347
rect 11848 25316 12725 25344
rect 11848 25304 11854 25316
rect 12713 25313 12725 25316
rect 12759 25313 12771 25347
rect 12713 25307 12771 25313
rect 13538 25304 13544 25356
rect 13596 25344 13602 25356
rect 14277 25347 14335 25353
rect 14277 25344 14289 25347
rect 13596 25316 14289 25344
rect 13596 25304 13602 25316
rect 14277 25313 14289 25316
rect 14323 25313 14335 25347
rect 14458 25344 14464 25356
rect 14419 25316 14464 25344
rect 14277 25307 14335 25313
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 15930 25344 15936 25356
rect 15891 25316 15936 25344
rect 15930 25304 15936 25316
rect 15988 25304 15994 25356
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25344 16175 25347
rect 17494 25344 17500 25356
rect 16163 25316 17500 25344
rect 16163 25313 16175 25316
rect 16117 25307 16175 25313
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 1762 25276 1768 25288
rect 1723 25248 1768 25276
rect 1762 25236 1768 25248
rect 1820 25236 1826 25288
rect 5169 25279 5227 25285
rect 5169 25245 5181 25279
rect 5215 25276 5227 25279
rect 7190 25276 7196 25288
rect 5215 25248 7196 25276
rect 5215 25245 5227 25248
rect 5169 25239 5227 25245
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 9953 25279 10011 25285
rect 9953 25276 9965 25279
rect 9916 25248 9965 25276
rect 9916 25236 9922 25248
rect 9953 25245 9965 25248
rect 9999 25245 10011 25279
rect 9953 25239 10011 25245
rect 11514 25236 11520 25288
rect 11572 25276 11578 25288
rect 12529 25279 12587 25285
rect 12529 25276 12541 25279
rect 11572 25248 12541 25276
rect 11572 25236 11578 25248
rect 12529 25245 12541 25248
rect 12575 25276 12587 25279
rect 14182 25276 14188 25288
rect 12575 25248 14188 25276
rect 12575 25245 12587 25248
rect 12529 25239 12587 25245
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 17218 25276 17224 25288
rect 17179 25248 17224 25276
rect 17218 25236 17224 25248
rect 17276 25236 17282 25288
rect 23566 25276 23572 25288
rect 23527 25248 23572 25276
rect 23566 25236 23572 25248
rect 23624 25236 23630 25288
rect 38286 25276 38292 25288
rect 38247 25248 38292 25276
rect 38286 25236 38292 25248
rect 38344 25236 38350 25288
rect 4985 25143 5043 25149
rect 4985 25109 4997 25143
rect 5031 25140 5043 25143
rect 5166 25140 5172 25152
rect 5031 25112 5172 25140
rect 5031 25109 5043 25112
rect 4985 25103 5043 25109
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 13173 25143 13231 25149
rect 13173 25109 13185 25143
rect 13219 25140 13231 25143
rect 13354 25140 13360 25152
rect 13219 25112 13360 25140
rect 13219 25109 13231 25112
rect 13173 25103 13231 25109
rect 13354 25100 13360 25112
rect 13412 25100 13418 25152
rect 16574 25140 16580 25152
rect 16535 25112 16580 25140
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 17034 25140 17040 25152
rect 16995 25112 17040 25140
rect 17034 25100 17040 25112
rect 17092 25100 17098 25152
rect 20346 25140 20352 25152
rect 20307 25112 20352 25140
rect 20346 25100 20352 25112
rect 20404 25100 20410 25152
rect 23382 25140 23388 25152
rect 23343 25112 23388 25140
rect 23382 25100 23388 25112
rect 23440 25100 23446 25152
rect 33962 25100 33968 25152
rect 34020 25140 34026 25152
rect 38105 25143 38163 25149
rect 38105 25140 38117 25143
rect 34020 25112 38117 25140
rect 34020 25100 34026 25112
rect 38105 25109 38117 25112
rect 38151 25109 38163 25143
rect 38105 25103 38163 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 14369 24939 14427 24945
rect 14369 24905 14381 24939
rect 14415 24936 14427 24939
rect 14734 24936 14740 24948
rect 14415 24908 14740 24936
rect 14415 24905 14427 24908
rect 14369 24899 14427 24905
rect 14734 24896 14740 24908
rect 14792 24896 14798 24948
rect 15194 24868 15200 24880
rect 15155 24840 15200 24868
rect 15194 24828 15200 24840
rect 15252 24828 15258 24880
rect 17034 24868 17040 24880
rect 16995 24840 17040 24868
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 5166 24800 5172 24812
rect 5127 24772 5172 24800
rect 5166 24760 5172 24772
rect 5224 24760 5230 24812
rect 7282 24800 7288 24812
rect 7243 24772 7288 24800
rect 7282 24760 7288 24772
rect 7340 24760 7346 24812
rect 8846 24800 8852 24812
rect 8807 24772 8852 24800
rect 8846 24760 8852 24772
rect 8904 24760 8910 24812
rect 9858 24760 9864 24812
rect 9916 24800 9922 24812
rect 9953 24803 10011 24809
rect 9953 24800 9965 24803
rect 9916 24772 9965 24800
rect 9916 24760 9922 24772
rect 9953 24769 9965 24772
rect 9999 24769 10011 24803
rect 9953 24763 10011 24769
rect 11238 24760 11244 24812
rect 11296 24800 11302 24812
rect 11977 24803 12035 24809
rect 11977 24800 11989 24803
rect 11296 24772 11989 24800
rect 11296 24760 11302 24772
rect 11977 24769 11989 24772
rect 12023 24769 12035 24803
rect 11977 24763 12035 24769
rect 12342 24760 12348 24812
rect 12400 24800 12406 24812
rect 12621 24803 12679 24809
rect 12621 24800 12633 24803
rect 12400 24772 12633 24800
rect 12400 24760 12406 24772
rect 12621 24769 12633 24772
rect 12667 24769 12679 24803
rect 12621 24763 12679 24769
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24769 13323 24803
rect 13265 24763 13323 24769
rect 9033 24735 9091 24741
rect 9033 24701 9045 24735
rect 9079 24732 9091 24735
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9079 24704 10057 24732
rect 9079 24701 9091 24704
rect 9033 24695 9091 24701
rect 10045 24701 10057 24704
rect 10091 24701 10103 24735
rect 13280 24732 13308 24763
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13909 24803 13967 24809
rect 13412 24772 13860 24800
rect 13412 24760 13418 24772
rect 13722 24732 13728 24744
rect 10045 24695 10103 24701
rect 12452 24704 13308 24732
rect 13683 24704 13728 24732
rect 12452 24673 12480 24704
rect 13722 24692 13728 24704
rect 13780 24692 13786 24744
rect 13832 24732 13860 24772
rect 13909 24769 13921 24803
rect 13955 24800 13967 24803
rect 14274 24800 14280 24812
rect 13955 24772 14280 24800
rect 13955 24769 13967 24772
rect 13909 24763 13967 24769
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 20346 24800 20352 24812
rect 20307 24772 20352 24800
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 20530 24800 20536 24812
rect 20491 24772 20536 24800
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 22002 24760 22008 24812
rect 22060 24800 22066 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 22060 24772 22201 24800
rect 22060 24760 22066 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 22554 24760 22560 24812
rect 22612 24800 22618 24812
rect 23293 24803 23351 24809
rect 23293 24800 23305 24803
rect 22612 24772 23305 24800
rect 22612 24760 22618 24772
rect 23293 24769 23305 24772
rect 23339 24800 23351 24803
rect 23474 24800 23480 24812
rect 23339 24772 23480 24800
rect 23339 24769 23351 24772
rect 23293 24763 23351 24769
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 33318 24800 33324 24812
rect 33279 24772 33324 24800
rect 33318 24760 33324 24772
rect 33376 24760 33382 24812
rect 35526 24800 35532 24812
rect 35487 24772 35532 24800
rect 35526 24760 35532 24772
rect 35584 24760 35590 24812
rect 35621 24803 35679 24809
rect 35621 24769 35633 24803
rect 35667 24800 35679 24803
rect 36906 24800 36912 24812
rect 35667 24772 36912 24800
rect 35667 24769 35679 24772
rect 35621 24763 35679 24769
rect 36906 24760 36912 24772
rect 36964 24760 36970 24812
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 13832 24704 15117 24732
rect 15105 24701 15117 24704
rect 15151 24701 15163 24735
rect 15105 24695 15163 24701
rect 16574 24692 16580 24744
rect 16632 24732 16638 24744
rect 16945 24735 17003 24741
rect 16945 24732 16957 24735
rect 16632 24704 16957 24732
rect 16632 24692 16638 24704
rect 16945 24701 16957 24704
rect 16991 24701 17003 24735
rect 22646 24732 22652 24744
rect 22607 24704 22652 24732
rect 16945 24695 17003 24701
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 9493 24667 9551 24673
rect 9493 24633 9505 24667
rect 9539 24664 9551 24667
rect 12437 24667 12495 24673
rect 9539 24636 11928 24664
rect 9539 24633 9551 24636
rect 9493 24627 9551 24633
rect 4982 24596 4988 24608
rect 4943 24568 4988 24596
rect 4982 24556 4988 24568
rect 5040 24556 5046 24608
rect 7101 24599 7159 24605
rect 7101 24565 7113 24599
rect 7147 24596 7159 24599
rect 7558 24596 7564 24608
rect 7147 24568 7564 24596
rect 7147 24565 7159 24568
rect 7101 24559 7159 24565
rect 7558 24556 7564 24568
rect 7616 24556 7622 24608
rect 11790 24596 11796 24608
rect 11751 24568 11796 24596
rect 11790 24556 11796 24568
rect 11848 24556 11854 24608
rect 11900 24596 11928 24636
rect 12437 24633 12449 24667
rect 12483 24633 12495 24667
rect 13740 24664 13768 24692
rect 12437 24627 12495 24633
rect 13004 24636 13768 24664
rect 15657 24667 15715 24673
rect 13004 24596 13032 24636
rect 15657 24633 15669 24667
rect 15703 24664 15715 24667
rect 17497 24667 17555 24673
rect 17497 24664 17509 24667
rect 15703 24636 17509 24664
rect 15703 24633 15715 24636
rect 15657 24627 15715 24633
rect 17497 24633 17509 24636
rect 17543 24664 17555 24667
rect 32766 24664 32772 24676
rect 17543 24636 32772 24664
rect 17543 24633 17555 24636
rect 17497 24627 17555 24633
rect 32766 24624 32772 24636
rect 32824 24624 32830 24676
rect 11900 24568 13032 24596
rect 13081 24599 13139 24605
rect 13081 24565 13093 24599
rect 13127 24596 13139 24599
rect 13170 24596 13176 24608
rect 13127 24568 13176 24596
rect 13127 24565 13139 24568
rect 13081 24559 13139 24565
rect 13170 24556 13176 24568
rect 13228 24556 13234 24608
rect 20806 24596 20812 24608
rect 20767 24568 20812 24596
rect 20806 24556 20812 24568
rect 20864 24556 20870 24608
rect 21450 24556 21456 24608
rect 21508 24596 21514 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21508 24568 22017 24596
rect 21508 24556 21514 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22005 24559 22063 24565
rect 22738 24556 22744 24608
rect 22796 24596 22802 24608
rect 23385 24599 23443 24605
rect 23385 24596 23397 24599
rect 22796 24568 23397 24596
rect 22796 24556 22802 24568
rect 23385 24565 23397 24568
rect 23431 24565 23443 24599
rect 33410 24596 33416 24608
rect 33371 24568 33416 24596
rect 23385 24559 23443 24565
rect 33410 24556 33416 24568
rect 33468 24556 33474 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 13722 24352 13728 24404
rect 13780 24392 13786 24404
rect 15197 24395 15255 24401
rect 15197 24392 15209 24395
rect 13780 24364 15209 24392
rect 13780 24352 13786 24364
rect 15197 24361 15209 24364
rect 15243 24361 15255 24395
rect 16574 24392 16580 24404
rect 16535 24364 16580 24392
rect 15197 24355 15255 24361
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 20806 24392 20812 24404
rect 20767 24364 20812 24392
rect 20806 24352 20812 24364
rect 20864 24352 20870 24404
rect 12618 24256 12624 24268
rect 11624 24228 12624 24256
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 2314 24188 2320 24200
rect 2275 24160 2320 24188
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 4154 24188 4160 24200
rect 4115 24160 4160 24188
rect 4154 24148 4160 24160
rect 4212 24148 4218 24200
rect 7558 24188 7564 24200
rect 7519 24160 7564 24188
rect 7558 24148 7564 24160
rect 7616 24148 7622 24200
rect 11624 24197 11652 24228
rect 12618 24216 12624 24228
rect 12676 24216 12682 24268
rect 13998 24216 14004 24268
rect 14056 24256 14062 24268
rect 15013 24259 15071 24265
rect 15013 24256 15025 24259
rect 14056 24228 15025 24256
rect 14056 24216 14062 24228
rect 15013 24225 15025 24228
rect 15059 24225 15071 24259
rect 16206 24256 16212 24268
rect 16167 24228 16212 24256
rect 15013 24219 15071 24225
rect 16206 24216 16212 24228
rect 16264 24216 16270 24268
rect 16393 24259 16451 24265
rect 16393 24225 16405 24259
rect 16439 24256 16451 24259
rect 16942 24256 16948 24268
rect 16439 24228 16948 24256
rect 16439 24225 16451 24228
rect 16393 24219 16451 24225
rect 16942 24216 16948 24228
rect 17000 24216 17006 24268
rect 20162 24256 20168 24268
rect 20123 24228 20168 24256
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 20349 24259 20407 24265
rect 20349 24225 20361 24259
rect 20395 24256 20407 24259
rect 20438 24256 20444 24268
rect 20395 24228 20444 24256
rect 20395 24225 20407 24228
rect 20349 24219 20407 24225
rect 20438 24216 20444 24228
rect 20496 24216 20502 24268
rect 20824 24256 20852 24352
rect 21634 24284 21640 24336
rect 21692 24324 21698 24336
rect 21910 24324 21916 24336
rect 21692 24296 21916 24324
rect 21692 24284 21698 24296
rect 21910 24284 21916 24296
rect 21968 24284 21974 24336
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 20824 24228 21373 24256
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 22738 24256 22744 24268
rect 22699 24228 22744 24256
rect 21361 24219 21419 24225
rect 22738 24216 22744 24228
rect 22796 24216 22802 24268
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24157 11667 24191
rect 11609 24151 11667 24157
rect 11790 24148 11796 24200
rect 11848 24188 11854 24200
rect 12437 24191 12495 24197
rect 12437 24188 12449 24191
rect 11848 24160 12449 24188
rect 11848 24148 11854 24160
rect 12437 24157 12449 24160
rect 12483 24157 12495 24191
rect 12437 24151 12495 24157
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 11514 24080 11520 24132
rect 11572 24120 11578 24132
rect 12342 24120 12348 24132
rect 11572 24092 12348 24120
rect 11572 24080 11578 24092
rect 12342 24080 12348 24092
rect 12400 24120 12406 24132
rect 12912 24120 12940 24151
rect 13078 24148 13084 24200
rect 13136 24188 13142 24200
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 13136 24160 13737 24188
rect 13136 24148 13142 24160
rect 13725 24157 13737 24160
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 14829 24191 14887 24197
rect 14829 24157 14841 24191
rect 14875 24157 14887 24191
rect 16224 24188 16252 24216
rect 17954 24188 17960 24200
rect 16224 24160 17960 24188
rect 14829 24151 14887 24157
rect 12400 24092 12940 24120
rect 14844 24120 14872 24151
rect 17954 24148 17960 24160
rect 18012 24148 18018 24200
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 24762 24188 24768 24200
rect 24723 24160 24768 24188
rect 22557 24151 22615 24157
rect 17862 24120 17868 24132
rect 14844 24092 17868 24120
rect 12400 24080 12406 24092
rect 17862 24080 17868 24092
rect 17920 24080 17926 24132
rect 21450 24080 21456 24132
rect 21508 24120 21514 24132
rect 22572 24120 22600 24151
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 38286 24188 38292 24200
rect 38247 24160 38292 24188
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 33686 24120 33692 24132
rect 21508 24092 21553 24120
rect 22572 24092 33692 24120
rect 21508 24080 21514 24092
rect 33686 24080 33692 24092
rect 33744 24080 33750 24132
rect 1762 24052 1768 24064
rect 1723 24024 1768 24052
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 1946 24012 1952 24064
rect 2004 24052 2010 24064
rect 2409 24055 2467 24061
rect 2409 24052 2421 24055
rect 2004 24024 2421 24052
rect 2004 24012 2010 24024
rect 2409 24021 2421 24024
rect 2455 24021 2467 24055
rect 2409 24015 2467 24021
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 5074 24052 5080 24064
rect 4019 24024 5080 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 5074 24012 5080 24024
rect 5132 24012 5138 24064
rect 6730 24052 6736 24064
rect 6691 24024 6736 24052
rect 6730 24012 6736 24024
rect 6788 24012 6794 24064
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7377 24055 7435 24061
rect 7377 24052 7389 24055
rect 6972 24024 7389 24052
rect 6972 24012 6978 24024
rect 7377 24021 7389 24024
rect 7423 24021 7435 24055
rect 7377 24015 7435 24021
rect 11701 24055 11759 24061
rect 11701 24021 11713 24055
rect 11747 24052 11759 24055
rect 12066 24052 12072 24064
rect 11747 24024 12072 24052
rect 11747 24021 11759 24024
rect 11701 24015 11759 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 12253 24055 12311 24061
rect 12253 24021 12265 24055
rect 12299 24052 12311 24055
rect 12802 24052 12808 24064
rect 12299 24024 12808 24052
rect 12299 24021 12311 24024
rect 12253 24015 12311 24021
rect 12802 24012 12808 24024
rect 12860 24012 12866 24064
rect 12986 24052 12992 24064
rect 12947 24024 12992 24052
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 13541 24055 13599 24061
rect 13541 24021 13553 24055
rect 13587 24052 13599 24055
rect 14458 24052 14464 24064
rect 13587 24024 14464 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 23198 24052 23204 24064
rect 23159 24024 23204 24052
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 24581 24055 24639 24061
rect 24581 24021 24593 24055
rect 24627 24052 24639 24055
rect 25222 24052 25228 24064
rect 24627 24024 25228 24052
rect 24627 24021 24639 24024
rect 24581 24015 24639 24021
rect 25222 24012 25228 24024
rect 25280 24012 25286 24064
rect 36998 24012 37004 24064
rect 37056 24052 37062 24064
rect 38105 24055 38163 24061
rect 38105 24052 38117 24055
rect 37056 24024 38117 24052
rect 37056 24012 37062 24024
rect 38105 24021 38117 24024
rect 38151 24021 38163 24055
rect 38105 24015 38163 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 1765 23851 1823 23857
rect 1765 23848 1777 23851
rect 1636 23820 1777 23848
rect 1636 23808 1642 23820
rect 1765 23817 1777 23820
rect 1811 23817 1823 23851
rect 1765 23811 1823 23817
rect 10321 23851 10379 23857
rect 10321 23817 10333 23851
rect 10367 23817 10379 23851
rect 10321 23811 10379 23817
rect 10336 23780 10364 23811
rect 10870 23808 10876 23860
rect 10928 23848 10934 23860
rect 12529 23851 12587 23857
rect 10928 23820 12434 23848
rect 10928 23808 10934 23820
rect 12406 23780 12434 23820
rect 12529 23817 12541 23851
rect 12575 23848 12587 23851
rect 13078 23848 13084 23860
rect 12575 23820 13084 23848
rect 12575 23817 12587 23820
rect 12529 23811 12587 23817
rect 13078 23808 13084 23820
rect 13136 23808 13142 23860
rect 13173 23851 13231 23857
rect 13173 23817 13185 23851
rect 13219 23848 13231 23851
rect 14461 23851 14519 23857
rect 13219 23820 13952 23848
rect 13219 23817 13231 23820
rect 13173 23811 13231 23817
rect 10336 23752 11192 23780
rect 12406 23752 13400 23780
rect 1946 23712 1952 23724
rect 1907 23684 1952 23712
rect 1946 23672 1952 23684
rect 2004 23672 2010 23724
rect 2130 23672 2136 23724
rect 2188 23712 2194 23724
rect 2501 23715 2559 23721
rect 2501 23712 2513 23715
rect 2188 23684 2513 23712
rect 2188 23672 2194 23684
rect 2501 23681 2513 23684
rect 2547 23712 2559 23715
rect 2682 23712 2688 23724
rect 2547 23684 2688 23712
rect 2547 23681 2559 23684
rect 2501 23675 2559 23681
rect 2682 23672 2688 23684
rect 2740 23712 2746 23724
rect 3145 23715 3203 23721
rect 3145 23712 3157 23715
rect 2740 23684 3157 23712
rect 2740 23672 2746 23684
rect 3145 23681 3157 23684
rect 3191 23681 3203 23715
rect 3878 23712 3884 23724
rect 3839 23684 3884 23712
rect 3145 23675 3203 23681
rect 3878 23672 3884 23684
rect 3936 23672 3942 23724
rect 4525 23715 4583 23721
rect 4525 23681 4537 23715
rect 4571 23681 4583 23715
rect 5350 23712 5356 23724
rect 5311 23684 5356 23712
rect 4525 23675 4583 23681
rect 2590 23604 2596 23656
rect 2648 23644 2654 23656
rect 4154 23644 4160 23656
rect 2648 23616 4160 23644
rect 2648 23604 2654 23616
rect 4154 23604 4160 23616
rect 4212 23644 4218 23656
rect 4540 23644 4568 23675
rect 5350 23672 5356 23684
rect 5408 23672 5414 23724
rect 5718 23672 5724 23724
rect 5776 23712 5782 23724
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 5776 23684 7021 23712
rect 5776 23672 5782 23684
rect 7009 23681 7021 23684
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 7190 23672 7196 23724
rect 7248 23712 7254 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7248 23684 7665 23712
rect 7248 23672 7254 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 9398 23712 9404 23724
rect 9359 23684 9404 23712
rect 7653 23675 7711 23681
rect 9398 23672 9404 23684
rect 9456 23672 9462 23724
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23712 10563 23715
rect 10962 23712 10968 23724
rect 10551 23684 10968 23712
rect 10551 23681 10563 23684
rect 10505 23675 10563 23681
rect 10962 23672 10968 23684
rect 11020 23672 11026 23724
rect 11164 23721 11192 23752
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 13372 23721 13400 23752
rect 12713 23715 12771 23721
rect 12713 23712 12725 23715
rect 12676 23684 12725 23712
rect 12676 23672 12682 23684
rect 12713 23681 12725 23684
rect 12759 23681 12771 23715
rect 12713 23675 12771 23681
rect 13357 23715 13415 23721
rect 13357 23681 13369 23715
rect 13403 23712 13415 23715
rect 13817 23715 13875 23721
rect 13817 23712 13829 23715
rect 13403 23684 13829 23712
rect 13403 23681 13415 23684
rect 13357 23675 13415 23681
rect 13817 23681 13829 23684
rect 13863 23681 13875 23715
rect 13924 23712 13952 23820
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 20349 23851 20407 23857
rect 14507 23820 15332 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 15304 23789 15332 23820
rect 20349 23817 20361 23851
rect 20395 23817 20407 23851
rect 22002 23848 22008 23860
rect 21963 23820 22008 23848
rect 20349 23811 20407 23817
rect 15289 23783 15347 23789
rect 15289 23749 15301 23783
rect 15335 23749 15347 23783
rect 15838 23780 15844 23792
rect 15799 23752 15844 23780
rect 15289 23743 15347 23749
rect 15838 23740 15844 23752
rect 15896 23740 15902 23792
rect 20364 23780 20392 23811
rect 22002 23808 22008 23820
rect 22060 23808 22066 23860
rect 23198 23808 23204 23860
rect 23256 23848 23262 23860
rect 23293 23851 23351 23857
rect 23293 23848 23305 23851
rect 23256 23820 23305 23848
rect 23256 23808 23262 23820
rect 23293 23817 23305 23820
rect 23339 23817 23351 23851
rect 23293 23811 23351 23817
rect 24762 23780 24768 23792
rect 20364 23752 21220 23780
rect 14645 23715 14703 23721
rect 14645 23712 14657 23715
rect 13924 23684 14657 23712
rect 13817 23675 13875 23681
rect 14645 23681 14657 23684
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23681 17647 23715
rect 18414 23712 18420 23724
rect 18375 23684 18420 23712
rect 17589 23675 17647 23681
rect 4212 23616 4568 23644
rect 4212 23604 4218 23616
rect 6822 23604 6828 23656
rect 6880 23644 6886 23656
rect 11885 23647 11943 23653
rect 6880 23616 9720 23644
rect 6880 23604 6886 23616
rect 3973 23579 4031 23585
rect 3973 23545 3985 23579
rect 4019 23576 4031 23579
rect 4890 23576 4896 23588
rect 4019 23548 4896 23576
rect 4019 23545 4031 23548
rect 3973 23539 4031 23545
rect 4890 23536 4896 23548
rect 4948 23536 4954 23588
rect 7101 23579 7159 23585
rect 7101 23545 7113 23579
rect 7147 23576 7159 23579
rect 9582 23576 9588 23588
rect 7147 23548 9588 23576
rect 7147 23545 7159 23548
rect 7101 23539 7159 23545
rect 9582 23536 9588 23548
rect 9640 23536 9646 23588
rect 9692 23576 9720 23616
rect 11885 23613 11897 23647
rect 11931 23644 11943 23647
rect 13078 23644 13084 23656
rect 11931 23616 13084 23644
rect 11931 23613 11943 23616
rect 11885 23607 11943 23613
rect 13078 23604 13084 23616
rect 13136 23604 13142 23656
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23644 15255 23647
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 15243 23616 16865 23644
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 16853 23613 16865 23616
rect 16899 23613 16911 23647
rect 16853 23607 16911 23613
rect 17604 23644 17632 23675
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23712 19303 23715
rect 20070 23712 20076 23724
rect 19291 23684 20076 23712
rect 19291 23681 19303 23684
rect 19245 23675 19303 23681
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 21192 23721 21220 23752
rect 22066 23752 24768 23780
rect 20533 23715 20591 23721
rect 20533 23681 20545 23715
rect 20579 23681 20591 23715
rect 20533 23675 20591 23681
rect 21177 23715 21235 23721
rect 21177 23681 21189 23715
rect 21223 23681 21235 23715
rect 21177 23675 21235 23681
rect 20548 23644 20576 23675
rect 22066 23644 22094 23752
rect 24762 23740 24768 23752
rect 24820 23740 24826 23792
rect 22186 23712 22192 23724
rect 22147 23684 22192 23712
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 22646 23712 22652 23724
rect 22607 23684 22652 23712
rect 22646 23672 22652 23684
rect 22704 23672 22710 23724
rect 22833 23715 22891 23721
rect 22833 23681 22845 23715
rect 22879 23712 22891 23715
rect 23382 23712 23388 23724
rect 22879 23684 23388 23712
rect 22879 23681 22891 23684
rect 22833 23675 22891 23681
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 23937 23715 23995 23721
rect 23937 23681 23949 23715
rect 23983 23712 23995 23715
rect 25222 23712 25228 23724
rect 23983 23684 25084 23712
rect 25183 23684 25228 23712
rect 23983 23681 23995 23684
rect 23937 23675 23995 23681
rect 24394 23644 24400 23656
rect 17604 23616 22094 23644
rect 24355 23616 24400 23644
rect 17604 23576 17632 23616
rect 24394 23604 24400 23616
rect 24452 23604 24458 23656
rect 25056 23644 25084 23684
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 25498 23644 25504 23656
rect 25056 23616 25504 23644
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 9692 23548 12434 23576
rect 2593 23511 2651 23517
rect 2593 23477 2605 23511
rect 2639 23508 2651 23511
rect 2866 23508 2872 23520
rect 2639 23480 2872 23508
rect 2639 23477 2651 23480
rect 2593 23471 2651 23477
rect 2866 23468 2872 23480
rect 2924 23468 2930 23520
rect 3142 23468 3148 23520
rect 3200 23508 3206 23520
rect 3237 23511 3295 23517
rect 3237 23508 3249 23511
rect 3200 23480 3249 23508
rect 3200 23468 3206 23480
rect 3237 23477 3249 23480
rect 3283 23477 3295 23511
rect 4614 23508 4620 23520
rect 4575 23480 4620 23508
rect 3237 23471 3295 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 5169 23511 5227 23517
rect 5169 23477 5181 23511
rect 5215 23508 5227 23511
rect 6638 23508 6644 23520
rect 5215 23480 6644 23508
rect 5215 23477 5227 23480
rect 5169 23471 5227 23477
rect 6638 23468 6644 23480
rect 6696 23468 6702 23520
rect 7745 23511 7803 23517
rect 7745 23477 7757 23511
rect 7791 23508 7803 23511
rect 8018 23508 8024 23520
rect 7791 23480 8024 23508
rect 7791 23477 7803 23480
rect 7745 23471 7803 23477
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 9217 23511 9275 23517
rect 9217 23477 9229 23511
rect 9263 23508 9275 23511
rect 9674 23508 9680 23520
rect 9263 23480 9680 23508
rect 9263 23477 9275 23480
rect 9217 23471 9275 23477
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 10965 23511 11023 23517
rect 10965 23477 10977 23511
rect 11011 23508 11023 23511
rect 12250 23508 12256 23520
rect 11011 23480 12256 23508
rect 11011 23477 11023 23480
rect 10965 23471 11023 23477
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 12406 23508 12434 23548
rect 13832 23548 17632 23576
rect 13832 23508 13860 23548
rect 12406 23480 13860 23508
rect 13909 23511 13967 23517
rect 13909 23477 13921 23511
rect 13955 23508 13967 23511
rect 14826 23508 14832 23520
rect 13955 23480 14832 23508
rect 13955 23477 13967 23480
rect 13909 23471 13967 23477
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 17678 23508 17684 23520
rect 17639 23480 17684 23508
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18506 23508 18512 23520
rect 18467 23480 18512 23508
rect 18506 23468 18512 23480
rect 18564 23468 18570 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 19061 23511 19119 23517
rect 19061 23508 19073 23511
rect 18748 23480 19073 23508
rect 18748 23468 18754 23480
rect 19061 23477 19073 23480
rect 19107 23477 19119 23511
rect 20990 23508 20996 23520
rect 20951 23480 20996 23508
rect 19061 23471 19119 23477
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 23750 23508 23756 23520
rect 23711 23480 23756 23508
rect 23750 23468 23756 23480
rect 23808 23468 23814 23520
rect 25038 23508 25044 23520
rect 24999 23480 25044 23508
rect 25038 23468 25044 23480
rect 25096 23468 25102 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 8389 23307 8447 23313
rect 3988 23276 7420 23304
rect 1581 23239 1639 23245
rect 1581 23205 1593 23239
rect 1627 23236 1639 23239
rect 3878 23236 3884 23248
rect 1627 23208 3884 23236
rect 1627 23205 1639 23208
rect 1581 23199 1639 23205
rect 3878 23196 3884 23208
rect 3936 23196 3942 23248
rect 3988 23168 4016 23276
rect 4065 23239 4123 23245
rect 4065 23205 4077 23239
rect 4111 23236 4123 23239
rect 5534 23236 5540 23248
rect 4111 23208 5540 23236
rect 4111 23205 4123 23208
rect 4065 23199 4123 23205
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 7282 23236 7288 23248
rect 6012 23208 7288 23236
rect 4890 23168 4896 23180
rect 2608 23140 4016 23168
rect 4851 23140 4896 23168
rect 2608 23109 2636 23140
rect 4890 23128 4896 23140
rect 4948 23128 4954 23180
rect 4982 23128 4988 23180
rect 5040 23168 5046 23180
rect 5077 23171 5135 23177
rect 5077 23168 5089 23171
rect 5040 23140 5089 23168
rect 5040 23128 5046 23140
rect 5077 23137 5089 23140
rect 5123 23137 5135 23171
rect 5077 23131 5135 23137
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 2593 23103 2651 23109
rect 1811 23072 2544 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 2409 22967 2467 22973
rect 2409 22964 2421 22967
rect 1728 22936 2421 22964
rect 1728 22924 1734 22936
rect 2409 22933 2421 22936
rect 2455 22933 2467 22967
rect 2516 22964 2544 23072
rect 2593 23069 2605 23103
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 2682 23060 2688 23112
rect 2740 23100 2746 23112
rect 3145 23103 3203 23109
rect 3145 23100 3157 23103
rect 2740 23072 3157 23100
rect 2740 23060 2746 23072
rect 3145 23069 3157 23072
rect 3191 23100 3203 23103
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 3191 23072 3985 23100
rect 3191 23069 3203 23072
rect 3145 23063 3203 23069
rect 3973 23069 3985 23072
rect 4019 23100 4031 23103
rect 4154 23100 4160 23112
rect 4019 23072 4160 23100
rect 4019 23069 4031 23072
rect 3973 23063 4031 23069
rect 4154 23060 4160 23072
rect 4212 23060 4218 23112
rect 5166 23060 5172 23112
rect 5224 23100 5230 23112
rect 6012 23109 6040 23208
rect 7282 23196 7288 23208
rect 7340 23196 7346 23248
rect 7392 23236 7420 23276
rect 8389 23273 8401 23307
rect 8435 23304 8447 23307
rect 9398 23304 9404 23316
rect 8435 23276 9404 23304
rect 8435 23273 8447 23276
rect 8389 23267 8447 23273
rect 9398 23264 9404 23276
rect 9456 23264 9462 23316
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 20070 23304 20076 23316
rect 12492 23276 16620 23304
rect 20031 23276 20076 23304
rect 12492 23264 12498 23276
rect 9306 23236 9312 23248
rect 7392 23208 9312 23236
rect 9306 23196 9312 23208
rect 9364 23196 9370 23248
rect 12529 23239 12587 23245
rect 12529 23205 12541 23239
rect 12575 23236 12587 23239
rect 14645 23239 14703 23245
rect 14645 23236 14657 23239
rect 12575 23208 14657 23236
rect 12575 23205 12587 23208
rect 12529 23199 12587 23205
rect 14645 23205 14657 23208
rect 14691 23236 14703 23239
rect 15010 23236 15016 23248
rect 14691 23208 15016 23236
rect 14691 23205 14703 23208
rect 14645 23199 14703 23205
rect 15010 23196 15016 23208
rect 15068 23196 15074 23248
rect 6730 23168 6736 23180
rect 6691 23140 6736 23168
rect 6730 23128 6736 23140
rect 6788 23128 6794 23180
rect 7374 23168 7380 23180
rect 7335 23140 7380 23168
rect 7374 23128 7380 23140
rect 7432 23128 7438 23180
rect 9674 23168 9680 23180
rect 9635 23140 9680 23168
rect 9674 23128 9680 23140
rect 9732 23128 9738 23180
rect 11882 23168 11888 23180
rect 11843 23140 11888 23168
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 12066 23168 12072 23180
rect 12027 23140 12072 23168
rect 12066 23128 12072 23140
rect 12124 23128 12130 23180
rect 13078 23168 13084 23180
rect 13039 23140 13084 23168
rect 13078 23128 13084 23140
rect 13136 23128 13142 23180
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23168 13783 23171
rect 14090 23168 14096 23180
rect 13771 23140 14096 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 14090 23128 14096 23140
rect 14148 23128 14154 23180
rect 14458 23168 14464 23180
rect 14419 23140 14464 23168
rect 14458 23128 14464 23140
rect 14516 23128 14522 23180
rect 16592 23168 16620 23276
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 20640 23276 20944 23304
rect 17773 23239 17831 23245
rect 17773 23205 17785 23239
rect 17819 23236 17831 23239
rect 20530 23236 20536 23248
rect 17819 23208 20536 23236
rect 17819 23205 17831 23208
rect 17773 23199 17831 23205
rect 20530 23196 20536 23208
rect 20588 23196 20594 23248
rect 17129 23171 17187 23177
rect 17129 23168 17141 23171
rect 16592 23140 17141 23168
rect 17129 23137 17141 23140
rect 17175 23137 17187 23171
rect 17129 23131 17187 23137
rect 17313 23171 17371 23177
rect 17313 23137 17325 23171
rect 17359 23168 17371 23171
rect 17678 23168 17684 23180
rect 17359 23140 17684 23168
rect 17359 23137 17371 23140
rect 17313 23131 17371 23137
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23168 18475 23171
rect 18506 23168 18512 23180
rect 18463 23140 18512 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 20640 23168 20668 23276
rect 20916 23236 20944 23276
rect 21358 23264 21364 23316
rect 21416 23304 21422 23316
rect 29822 23304 29828 23316
rect 21416 23276 29828 23304
rect 21416 23264 21422 23276
rect 29822 23264 29828 23276
rect 29880 23264 29886 23316
rect 28074 23236 28080 23248
rect 20916 23208 28080 23236
rect 28074 23196 28080 23208
rect 28132 23196 28138 23248
rect 20990 23168 20996 23180
rect 19536 23140 20668 23168
rect 20951 23140 20996 23168
rect 5997 23103 6055 23109
rect 5997 23100 6009 23103
rect 5224 23072 6009 23100
rect 5224 23060 5230 23072
rect 5997 23069 6009 23072
rect 6043 23069 6055 23103
rect 5997 23063 6055 23069
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23069 8631 23103
rect 8573 23063 8631 23069
rect 5537 23035 5595 23041
rect 5537 23001 5549 23035
rect 5583 23032 5595 23035
rect 6546 23032 6552 23044
rect 5583 23004 6552 23032
rect 5583 23001 5595 23004
rect 5537 22995 5595 23001
rect 6546 22992 6552 23004
rect 6604 22992 6610 23044
rect 6825 23035 6883 23041
rect 6825 23001 6837 23035
rect 6871 23032 6883 23035
rect 6914 23032 6920 23044
rect 6871 23004 6920 23032
rect 6871 23001 6883 23004
rect 6825 22995 6883 23001
rect 6914 22992 6920 23004
rect 6972 22992 6978 23044
rect 7558 22992 7564 23044
rect 7616 23032 7622 23044
rect 8588 23032 8616 23063
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 9456 23072 9505 23100
rect 9456 23060 9462 23072
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 11238 23100 11244 23112
rect 11199 23072 11244 23100
rect 9493 23063 9551 23069
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 14274 23100 14280 23112
rect 14235 23072 14280 23100
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 15378 23100 15384 23112
rect 15339 23072 15384 23100
rect 15378 23060 15384 23072
rect 15436 23100 15442 23112
rect 16209 23103 16267 23109
rect 16209 23100 16221 23103
rect 15436 23072 16221 23100
rect 15436 23060 15442 23072
rect 16209 23069 16221 23072
rect 16255 23069 16267 23103
rect 16209 23063 16267 23069
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 19536 23100 19564 23140
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 22373 23171 22431 23177
rect 22373 23137 22385 23171
rect 22419 23168 22431 23171
rect 23198 23168 23204 23180
rect 22419 23140 23204 23168
rect 22419 23137 22431 23140
rect 22373 23131 22431 23137
rect 23198 23128 23204 23140
rect 23256 23128 23262 23180
rect 24394 23128 24400 23180
rect 24452 23168 24458 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 24452 23140 24593 23168
rect 24452 23128 24458 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 24765 23171 24823 23177
rect 24765 23137 24777 23171
rect 24811 23168 24823 23171
rect 25038 23168 25044 23180
rect 24811 23140 25044 23168
rect 24811 23137 24823 23140
rect 24765 23131 24823 23137
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 18279 23072 19564 23100
rect 19613 23103 19671 23109
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 19613 23069 19625 23103
rect 19659 23100 19671 23103
rect 20162 23100 20168 23112
rect 19659 23072 20168 23100
rect 19659 23069 19671 23072
rect 19613 23063 19671 23069
rect 20162 23060 20168 23072
rect 20220 23060 20226 23112
rect 20257 23103 20315 23109
rect 20257 23069 20269 23103
rect 20303 23069 20315 23103
rect 20806 23100 20812 23112
rect 20767 23072 20812 23100
rect 20257 23063 20315 23069
rect 7616 23004 13124 23032
rect 7616 22992 7622 23004
rect 2774 22964 2780 22976
rect 2516 22936 2780 22964
rect 2409 22927 2467 22933
rect 2774 22924 2780 22936
rect 2832 22924 2838 22976
rect 3234 22964 3240 22976
rect 3195 22936 3240 22964
rect 3234 22924 3240 22936
rect 3292 22924 3298 22976
rect 6086 22964 6092 22976
rect 6047 22936 6092 22964
rect 6086 22924 6092 22936
rect 6144 22924 6150 22976
rect 9674 22924 9680 22976
rect 9732 22964 9738 22976
rect 10137 22967 10195 22973
rect 10137 22964 10149 22967
rect 9732 22936 10149 22964
rect 9732 22924 9738 22936
rect 10137 22933 10149 22936
rect 10183 22933 10195 22967
rect 10594 22964 10600 22976
rect 10555 22936 10600 22964
rect 10137 22927 10195 22933
rect 10594 22924 10600 22936
rect 10652 22924 10658 22976
rect 11333 22967 11391 22973
rect 11333 22933 11345 22967
rect 11379 22964 11391 22967
rect 12342 22964 12348 22976
rect 11379 22936 12348 22964
rect 11379 22933 11391 22936
rect 11333 22927 11391 22933
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 13096 22964 13124 23004
rect 13170 22992 13176 23044
rect 13228 23032 13234 23044
rect 16114 23032 16120 23044
rect 13228 23004 13273 23032
rect 15028 23004 16120 23032
rect 13228 22992 13234 23004
rect 15028 22964 15056 23004
rect 16114 22992 16120 23004
rect 16172 22992 16178 23044
rect 18414 22992 18420 23044
rect 18472 23032 18478 23044
rect 20272 23032 20300 23063
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 23566 23060 23572 23112
rect 23624 23100 23630 23112
rect 24029 23103 24087 23109
rect 24029 23100 24041 23103
rect 23624 23072 24041 23100
rect 23624 23060 23630 23072
rect 24029 23069 24041 23072
rect 24075 23069 24087 23103
rect 33962 23100 33968 23112
rect 33923 23072 33968 23100
rect 24029 23063 24087 23069
rect 33962 23060 33968 23072
rect 34020 23060 34026 23112
rect 18472 23004 20300 23032
rect 18472 22992 18478 23004
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 21453 23035 21511 23041
rect 21453 23032 21465 23035
rect 20588 23004 21465 23032
rect 20588 22992 20594 23004
rect 21453 23001 21465 23004
rect 21499 23032 21511 23035
rect 22094 23032 22100 23044
rect 21499 23004 22100 23032
rect 21499 23001 21511 23004
rect 21453 22995 21511 23001
rect 22094 22992 22100 23004
rect 22152 22992 22158 23044
rect 22462 22992 22468 23044
rect 22520 23032 22526 23044
rect 22520 23004 22565 23032
rect 22520 22992 22526 23004
rect 22646 22992 22652 23044
rect 22704 23032 22710 23044
rect 23385 23035 23443 23041
rect 23385 23032 23397 23035
rect 22704 23004 23397 23032
rect 22704 22992 22710 23004
rect 23385 23001 23397 23004
rect 23431 23032 23443 23035
rect 34790 23032 34796 23044
rect 23431 23004 34796 23032
rect 23431 23001 23443 23004
rect 23385 22995 23443 23001
rect 34790 22992 34796 23004
rect 34848 22992 34854 23044
rect 13096 22936 15056 22964
rect 15102 22924 15108 22976
rect 15160 22964 15166 22976
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 15160 22936 15485 22964
rect 15160 22924 15166 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 16022 22964 16028 22976
rect 15983 22936 16028 22964
rect 15473 22927 15531 22933
rect 16022 22924 16028 22936
rect 16080 22924 16086 22976
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 18877 22967 18935 22973
rect 18877 22964 18889 22967
rect 18656 22936 18889 22964
rect 18656 22924 18662 22936
rect 18877 22933 18889 22936
rect 18923 22933 18935 22967
rect 18877 22927 18935 22933
rect 19242 22924 19248 22976
rect 19300 22964 19306 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 19300 22936 19441 22964
rect 19300 22924 19306 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 19429 22927 19487 22933
rect 20806 22924 20812 22976
rect 20864 22964 20870 22976
rect 21358 22964 21364 22976
rect 20864 22936 21364 22964
rect 20864 22924 20870 22936
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23845 22967 23903 22973
rect 23845 22964 23857 22967
rect 23532 22936 23857 22964
rect 23532 22924 23538 22936
rect 23845 22933 23857 22936
rect 23891 22933 23903 22967
rect 23845 22927 23903 22933
rect 25038 22924 25044 22976
rect 25096 22964 25102 22976
rect 25225 22967 25283 22973
rect 25225 22964 25237 22967
rect 25096 22936 25237 22964
rect 25096 22924 25102 22936
rect 25225 22933 25237 22936
rect 25271 22933 25283 22967
rect 34054 22964 34060 22976
rect 34015 22936 34060 22964
rect 25225 22927 25283 22933
rect 34054 22924 34060 22936
rect 34112 22924 34118 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 9398 22760 9404 22772
rect 1627 22732 6592 22760
rect 9359 22732 9404 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 3878 22652 3884 22704
rect 3936 22652 3942 22704
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 4154 22584 4160 22636
rect 4212 22624 4218 22636
rect 4893 22627 4951 22633
rect 4893 22624 4905 22627
rect 4212 22596 4905 22624
rect 4212 22584 4218 22596
rect 4893 22593 4905 22596
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 5350 22584 5356 22636
rect 5408 22624 5414 22636
rect 5537 22627 5595 22633
rect 5537 22624 5549 22627
rect 5408 22596 5549 22624
rect 5408 22584 5414 22596
rect 5537 22593 5549 22596
rect 5583 22624 5595 22627
rect 6270 22624 6276 22636
rect 5583 22596 6276 22624
rect 5583 22593 5595 22596
rect 5537 22587 5595 22593
rect 6270 22584 6276 22596
rect 6328 22584 6334 22636
rect 6564 22633 6592 22732
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 15378 22760 15384 22772
rect 9646 22732 15384 22760
rect 8570 22652 8576 22704
rect 8628 22692 8634 22704
rect 9646 22692 9674 22732
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 18230 22720 18236 22772
rect 18288 22760 18294 22772
rect 18598 22760 18604 22772
rect 18288 22732 18604 22760
rect 18288 22720 18294 22732
rect 18598 22720 18604 22732
rect 18656 22720 18662 22772
rect 20162 22760 20168 22772
rect 20123 22732 20168 22760
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 25038 22760 25044 22772
rect 23308 22732 25044 22760
rect 8628 22664 9674 22692
rect 8628 22652 8634 22664
rect 10594 22652 10600 22704
rect 10652 22692 10658 22704
rect 12161 22695 12219 22701
rect 12161 22692 12173 22695
rect 10652 22664 12173 22692
rect 10652 22652 10658 22664
rect 12161 22661 12173 22664
rect 12207 22661 12219 22695
rect 12161 22655 12219 22661
rect 12250 22652 12256 22704
rect 12308 22692 12314 22704
rect 12805 22695 12863 22701
rect 12308 22664 12353 22692
rect 12308 22652 12314 22664
rect 12805 22661 12817 22695
rect 12851 22692 12863 22695
rect 12894 22692 12900 22704
rect 12851 22664 12900 22692
rect 12851 22661 12863 22664
rect 12805 22655 12863 22661
rect 12894 22652 12900 22664
rect 12952 22692 12958 22704
rect 13446 22692 13452 22704
rect 12952 22664 13452 22692
rect 12952 22652 12958 22664
rect 13446 22652 13452 22664
rect 13504 22652 13510 22704
rect 15102 22692 15108 22704
rect 15063 22664 15108 22692
rect 15102 22652 15108 22664
rect 15160 22652 15166 22704
rect 15654 22692 15660 22704
rect 15615 22664 15660 22692
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 23308 22701 23336 22732
rect 25038 22720 25044 22732
rect 25096 22720 25102 22772
rect 25498 22760 25504 22772
rect 25459 22732 25504 22760
rect 25498 22720 25504 22732
rect 25556 22720 25562 22772
rect 21361 22695 21419 22701
rect 21361 22661 21373 22695
rect 21407 22692 21419 22695
rect 22189 22695 22247 22701
rect 22189 22692 22201 22695
rect 21407 22664 22201 22692
rect 21407 22661 21419 22664
rect 21361 22655 21419 22661
rect 22189 22661 22201 22664
rect 22235 22661 22247 22695
rect 22189 22655 22247 22661
rect 23293 22695 23351 22701
rect 23293 22661 23305 22695
rect 23339 22661 23351 22695
rect 23293 22655 23351 22661
rect 23385 22695 23443 22701
rect 23385 22661 23397 22695
rect 23431 22692 23443 22695
rect 23474 22692 23480 22704
rect 23431 22664 23480 22692
rect 23431 22661 23443 22664
rect 23385 22655 23443 22661
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7285 22627 7343 22633
rect 7285 22624 7297 22627
rect 7248 22596 7297 22624
rect 7248 22584 7254 22596
rect 7285 22593 7297 22596
rect 7331 22624 7343 22627
rect 7558 22624 7564 22636
rect 7331 22596 7564 22624
rect 7331 22593 7343 22596
rect 7285 22587 7343 22593
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 8478 22624 8484 22636
rect 8439 22596 8484 22624
rect 8478 22584 8484 22596
rect 8536 22584 8542 22636
rect 9582 22584 9588 22636
rect 9640 22624 9646 22636
rect 10045 22627 10103 22633
rect 10045 22624 10057 22627
rect 9640 22596 10057 22624
rect 9640 22584 9646 22596
rect 10045 22593 10057 22596
rect 10091 22593 10103 22627
rect 10045 22587 10103 22593
rect 13817 22627 13875 22633
rect 13817 22593 13829 22627
rect 13863 22624 13875 22627
rect 14550 22624 14556 22636
rect 13863 22596 14556 22624
rect 13863 22593 13875 22596
rect 13817 22587 13875 22593
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 15930 22584 15936 22636
rect 15988 22624 15994 22636
rect 16114 22624 16120 22636
rect 15988 22596 16120 22624
rect 15988 22584 15994 22596
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 17037 22627 17095 22633
rect 17037 22624 17049 22627
rect 16540 22596 17049 22624
rect 16540 22584 16546 22596
rect 17037 22593 17049 22596
rect 17083 22593 17095 22627
rect 17954 22624 17960 22636
rect 17915 22596 17960 22624
rect 17037 22587 17095 22593
rect 17954 22584 17960 22596
rect 18012 22584 18018 22636
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22624 18199 22627
rect 18690 22624 18696 22636
rect 18187 22596 18696 22624
rect 18187 22593 18199 22596
rect 18141 22587 18199 22593
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 19242 22624 19248 22636
rect 19203 22596 19248 22624
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 20162 22584 20168 22636
rect 20220 22624 20226 22636
rect 20349 22627 20407 22633
rect 20349 22624 20361 22627
rect 20220 22596 20361 22624
rect 20220 22584 20226 22596
rect 20349 22593 20361 22596
rect 20395 22593 20407 22627
rect 21266 22624 21272 22636
rect 21227 22596 21272 22624
rect 20349 22587 20407 22593
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 25222 22584 25228 22636
rect 25280 22624 25286 22636
rect 25685 22627 25743 22633
rect 25685 22624 25697 22627
rect 25280 22596 25697 22624
rect 25280 22584 25286 22596
rect 25685 22593 25697 22596
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22624 32367 22627
rect 36998 22624 37004 22636
rect 32355 22596 37004 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 36998 22584 37004 22596
rect 37056 22584 37062 22636
rect 1578 22516 1584 22568
rect 1636 22556 1642 22568
rect 2593 22559 2651 22565
rect 2593 22556 2605 22559
rect 1636 22528 2605 22556
rect 1636 22516 1642 22528
rect 2593 22525 2605 22528
rect 2639 22525 2651 22559
rect 2593 22519 2651 22525
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 3510 22556 3516 22568
rect 2915 22528 3516 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 3510 22516 3516 22528
rect 3568 22516 3574 22568
rect 10226 22556 10232 22568
rect 10187 22528 10232 22556
rect 10226 22516 10232 22528
rect 10284 22516 10290 22568
rect 12802 22516 12808 22568
rect 12860 22556 12866 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 12860 22528 14013 22556
rect 12860 22516 12866 22528
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 15010 22556 15016 22568
rect 14971 22528 15016 22556
rect 14001 22519 14059 22525
rect 15010 22516 15016 22528
rect 15068 22516 15074 22568
rect 19058 22556 19064 22568
rect 19019 22528 19064 22556
rect 19058 22516 19064 22528
rect 19116 22516 19122 22568
rect 22094 22556 22100 22568
rect 22055 22528 22100 22556
rect 22094 22516 22100 22528
rect 22152 22516 22158 22568
rect 24394 22556 24400 22568
rect 24355 22528 24400 22556
rect 24394 22516 24400 22528
rect 24452 22516 24458 22568
rect 24581 22559 24639 22565
rect 24581 22525 24593 22559
rect 24627 22556 24639 22559
rect 25406 22556 25412 22568
rect 24627 22528 25412 22556
rect 24627 22525 24639 22528
rect 24581 22519 24639 22525
rect 25406 22516 25412 22528
rect 25464 22516 25470 22568
rect 7377 22491 7435 22497
rect 7377 22457 7389 22491
rect 7423 22488 7435 22491
rect 9214 22488 9220 22500
rect 7423 22460 9220 22488
rect 7423 22457 7435 22460
rect 7377 22451 7435 22457
rect 9214 22448 9220 22460
rect 9272 22448 9278 22500
rect 22649 22491 22707 22497
rect 22649 22457 22661 22491
rect 22695 22488 22707 22491
rect 23845 22491 23903 22497
rect 23845 22488 23857 22491
rect 22695 22460 23857 22488
rect 22695 22457 22707 22460
rect 22649 22451 22707 22457
rect 23845 22457 23857 22460
rect 23891 22488 23903 22491
rect 29730 22488 29736 22500
rect 23891 22460 29736 22488
rect 23891 22457 23903 22460
rect 23845 22451 23903 22457
rect 29730 22448 29736 22460
rect 29788 22448 29794 22500
rect 4341 22423 4399 22429
rect 4341 22389 4353 22423
rect 4387 22420 4399 22423
rect 4706 22420 4712 22432
rect 4387 22392 4712 22420
rect 4387 22389 4399 22392
rect 4341 22383 4399 22389
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 4982 22420 4988 22432
rect 4943 22392 4988 22420
rect 4982 22380 4988 22392
rect 5040 22380 5046 22432
rect 5629 22423 5687 22429
rect 5629 22389 5641 22423
rect 5675 22420 5687 22423
rect 5994 22420 6000 22432
rect 5675 22392 6000 22420
rect 5675 22389 5687 22392
rect 5629 22383 5687 22389
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 6362 22380 6368 22432
rect 6420 22420 6426 22432
rect 6641 22423 6699 22429
rect 6641 22420 6653 22423
rect 6420 22392 6653 22420
rect 6420 22380 6426 22392
rect 6641 22389 6653 22392
rect 6687 22389 6699 22423
rect 6641 22383 6699 22389
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 8297 22423 8355 22429
rect 8297 22420 8309 22423
rect 6972 22392 8309 22420
rect 6972 22380 6978 22392
rect 8297 22389 8309 22392
rect 8343 22389 8355 22423
rect 8297 22383 8355 22389
rect 10689 22423 10747 22429
rect 10689 22389 10701 22423
rect 10735 22420 10747 22423
rect 13906 22420 13912 22432
rect 10735 22392 13912 22420
rect 10735 22389 10747 22392
rect 10689 22383 10747 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 14185 22423 14243 22429
rect 14185 22420 14197 22423
rect 14056 22392 14197 22420
rect 14056 22380 14062 22392
rect 14185 22389 14197 22392
rect 14231 22389 14243 22423
rect 16206 22420 16212 22432
rect 16167 22392 16212 22420
rect 14185 22383 14243 22389
rect 16206 22380 16212 22392
rect 16264 22380 16270 22432
rect 16850 22420 16856 22432
rect 16811 22392 16856 22420
rect 16850 22380 16856 22392
rect 16908 22380 16914 22432
rect 19426 22420 19432 22432
rect 19387 22392 19432 22420
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 19518 22380 19524 22432
rect 19576 22420 19582 22432
rect 24946 22420 24952 22432
rect 19576 22392 24952 22420
rect 19576 22380 19582 22392
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 32398 22420 32404 22432
rect 32359 22392 32404 22420
rect 32398 22380 32404 22392
rect 32456 22380 32462 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1936 22219 1994 22225
rect 1936 22185 1948 22219
rect 1982 22216 1994 22219
rect 4065 22219 4123 22225
rect 4065 22216 4077 22219
rect 1982 22188 4077 22216
rect 1982 22185 1994 22188
rect 1936 22179 1994 22185
rect 4065 22185 4077 22188
rect 4111 22216 4123 22219
rect 4111 22188 6500 22216
rect 4111 22185 4123 22188
rect 4065 22179 4123 22185
rect 6472 22148 6500 22188
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 8205 22219 8263 22225
rect 8205 22216 8217 22219
rect 6696 22188 8217 22216
rect 6696 22176 6702 22188
rect 8205 22185 8217 22188
rect 8251 22185 8263 22219
rect 8205 22179 8263 22185
rect 9677 22219 9735 22225
rect 9677 22185 9689 22219
rect 9723 22216 9735 22219
rect 10226 22216 10232 22228
rect 9723 22188 10232 22216
rect 9723 22185 9735 22188
rect 9677 22179 9735 22185
rect 10226 22176 10232 22188
rect 10284 22176 10290 22228
rect 10584 22219 10642 22225
rect 10584 22185 10596 22219
rect 10630 22216 10642 22219
rect 11146 22216 11152 22228
rect 10630 22188 11152 22216
rect 10630 22185 10642 22188
rect 10584 22179 10642 22185
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 12268 22188 12848 22216
rect 6822 22148 6828 22160
rect 6472 22120 6828 22148
rect 6822 22108 6828 22120
rect 6880 22108 6886 22160
rect 12069 22151 12127 22157
rect 12069 22148 12081 22151
rect 11808 22120 12081 22148
rect 4157 22083 4215 22089
rect 4157 22080 4169 22083
rect 1688 22052 4169 22080
rect 1578 21972 1584 22024
rect 1636 22012 1642 22024
rect 1688 22021 1716 22052
rect 4157 22049 4169 22052
rect 4203 22049 4215 22083
rect 5626 22080 5632 22092
rect 4157 22043 4215 22049
rect 5552 22052 5632 22080
rect 1673 22015 1731 22021
rect 1673 22012 1685 22015
rect 1636 21984 1685 22012
rect 1636 21972 1642 21984
rect 1673 21981 1685 21984
rect 1719 21981 1731 22015
rect 5552 21998 5580 22052
rect 5626 22040 5632 22052
rect 5684 22040 5690 22092
rect 5902 22080 5908 22092
rect 5815 22052 5908 22080
rect 5902 22040 5908 22052
rect 5960 22080 5966 22092
rect 5960 22052 7972 22080
rect 5960 22040 5966 22052
rect 6365 22015 6423 22021
rect 1673 21975 1731 21981
rect 6365 21981 6377 22015
rect 6411 22012 6423 22015
rect 6730 22012 6736 22024
rect 6411 21984 6736 22012
rect 6411 21981 6423 21984
rect 6365 21975 6423 21981
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 7193 22015 7251 22021
rect 7193 22012 7205 22015
rect 7064 21984 7205 22012
rect 7064 21972 7070 21984
rect 7193 21981 7205 21984
rect 7239 22012 7251 22015
rect 7650 22012 7656 22024
rect 7239 21984 7656 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 7834 22012 7840 22024
rect 7795 21984 7840 22012
rect 7834 21972 7840 21984
rect 7892 21972 7898 22024
rect 2958 21904 2964 21956
rect 3016 21904 3022 21956
rect 4430 21944 4436 21956
rect 4391 21916 4436 21944
rect 4430 21904 4436 21916
rect 4488 21904 4494 21956
rect 7944 21944 7972 22052
rect 8018 22040 8024 22092
rect 8076 22080 8082 22092
rect 8478 22080 8484 22092
rect 8076 22052 8121 22080
rect 8312 22052 8484 22080
rect 8076 22040 8082 22052
rect 8110 21972 8116 22024
rect 8168 22012 8174 22024
rect 8312 22012 8340 22052
rect 8478 22040 8484 22052
rect 8536 22040 8542 22092
rect 10962 22040 10968 22092
rect 11020 22080 11026 22092
rect 11808 22080 11836 22120
rect 12069 22117 12081 22120
rect 12115 22117 12127 22151
rect 12069 22111 12127 22117
rect 11020 22052 11836 22080
rect 11020 22040 11026 22052
rect 8168 21984 8340 22012
rect 8168 21972 8174 21984
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9861 22015 9919 22021
rect 9861 22012 9873 22015
rect 8444 21984 9873 22012
rect 8444 21972 8450 21984
rect 9861 21981 9873 21984
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10321 22015 10379 22021
rect 10321 22012 10333 22015
rect 10008 21984 10333 22012
rect 10008 21972 10014 21984
rect 10321 21981 10333 21984
rect 10367 21981 10379 22015
rect 10321 21975 10379 21981
rect 10502 21944 10508 21956
rect 6012 21916 7788 21944
rect 7944 21916 10508 21944
rect 2682 21836 2688 21888
rect 2740 21876 2746 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 2740 21848 3433 21876
rect 2740 21836 2746 21848
rect 3421 21845 3433 21848
rect 3467 21876 3479 21879
rect 6012 21876 6040 21916
rect 6178 21876 6184 21888
rect 3467 21848 6040 21876
rect 6139 21848 6184 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 7098 21836 7104 21888
rect 7156 21876 7162 21888
rect 7285 21879 7343 21885
rect 7285 21876 7297 21879
rect 7156 21848 7297 21876
rect 7156 21836 7162 21848
rect 7285 21845 7297 21848
rect 7331 21845 7343 21879
rect 7760 21876 7788 21916
rect 10502 21904 10508 21916
rect 10560 21904 10566 21956
rect 11330 21904 11336 21956
rect 11388 21904 11394 21956
rect 12268 21876 12296 22188
rect 12342 22108 12348 22160
rect 12400 22148 12406 22160
rect 12820 22148 12848 22188
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 23290 22216 23296 22228
rect 14332 22188 23296 22216
rect 14332 22176 14338 22188
rect 23290 22176 23296 22188
rect 23348 22176 23354 22228
rect 24394 22176 24400 22228
rect 24452 22216 24458 22228
rect 33778 22216 33784 22228
rect 24452 22188 33784 22216
rect 24452 22176 24458 22188
rect 33778 22176 33784 22188
rect 33836 22176 33842 22228
rect 12400 22120 12756 22148
rect 12820 22120 18276 22148
rect 12400 22108 12406 22120
rect 12728 22089 12756 22120
rect 12714 22083 12772 22089
rect 12714 22049 12726 22083
rect 12760 22049 12772 22083
rect 16850 22080 16856 22092
rect 12714 22043 12772 22049
rect 16040 22052 16856 22080
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 21981 12587 22015
rect 12529 21975 12587 21981
rect 7760 21848 12296 21876
rect 7285 21839 7343 21845
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12544 21876 12572 21975
rect 12894 21972 12900 22024
rect 12952 22012 12958 22024
rect 14550 22012 14556 22024
rect 12952 21984 14556 22012
rect 12952 21972 12958 21984
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 15381 22015 15439 22021
rect 15381 21981 15393 22015
rect 15427 22012 15439 22015
rect 15746 22012 15752 22024
rect 15427 21984 15752 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 15746 21972 15752 21984
rect 15804 21972 15810 22024
rect 16040 22021 16068 22052
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16482 22012 16488 22024
rect 16443 21984 16488 22012
rect 16025 21975 16083 21981
rect 16482 21972 16488 21984
rect 16540 21972 16546 22024
rect 18248 22012 18276 22120
rect 19334 22108 19340 22160
rect 19392 22148 19398 22160
rect 24949 22151 25007 22157
rect 24949 22148 24961 22151
rect 19392 22120 19656 22148
rect 19392 22108 19398 22120
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 19058 22080 19064 22092
rect 18739 22052 19064 22080
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 19429 22083 19487 22089
rect 19429 22049 19441 22083
rect 19475 22080 19487 22083
rect 19518 22080 19524 22092
rect 19475 22052 19524 22080
rect 19475 22049 19487 22052
rect 19429 22043 19487 22049
rect 19518 22040 19524 22052
rect 19576 22040 19582 22092
rect 19628 22089 19656 22120
rect 23676 22120 24961 22148
rect 19613 22083 19671 22089
rect 19613 22049 19625 22083
rect 19659 22049 19671 22083
rect 21266 22080 21272 22092
rect 19613 22043 19671 22049
rect 20640 22052 21272 22080
rect 20640 22012 20668 22052
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 23106 22040 23112 22092
rect 23164 22080 23170 22092
rect 23676 22080 23704 22120
rect 24949 22117 24961 22120
rect 24995 22117 25007 22151
rect 24949 22111 25007 22117
rect 23164 22052 23704 22080
rect 23164 22040 23170 22052
rect 23750 22040 23756 22092
rect 23808 22080 23814 22092
rect 24765 22083 24823 22089
rect 24765 22080 24777 22083
rect 23808 22052 24777 22080
rect 23808 22040 23814 22052
rect 24765 22049 24777 22052
rect 24811 22049 24823 22083
rect 24765 22043 24823 22049
rect 25406 22040 25412 22092
rect 25464 22080 25470 22092
rect 26421 22083 26479 22089
rect 26421 22080 26433 22083
rect 25464 22052 26433 22080
rect 25464 22040 25470 22052
rect 26421 22049 26433 22052
rect 26467 22049 26479 22083
rect 26421 22043 26479 22049
rect 18248 21984 19334 22012
rect 13906 21904 13912 21956
rect 13964 21944 13970 21956
rect 14737 21947 14795 21953
rect 14737 21944 14749 21947
rect 13964 21916 14749 21944
rect 13964 21904 13970 21916
rect 14737 21913 14749 21916
rect 14783 21913 14795 21947
rect 14737 21907 14795 21913
rect 14826 21904 14832 21956
rect 14884 21944 14890 21956
rect 17589 21947 17647 21953
rect 14884 21916 14929 21944
rect 14884 21904 14890 21916
rect 17589 21913 17601 21947
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 12802 21876 12808 21888
rect 12492 21848 12808 21876
rect 12492 21836 12498 21848
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 13173 21879 13231 21885
rect 13173 21845 13185 21879
rect 13219 21876 13231 21879
rect 13998 21876 14004 21888
rect 13219 21848 14004 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13998 21836 14004 21848
rect 14056 21836 14062 21888
rect 15838 21876 15844 21888
rect 15799 21848 15844 21876
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 16577 21879 16635 21885
rect 16577 21845 16589 21879
rect 16623 21876 16635 21879
rect 16666 21876 16672 21888
rect 16623 21848 16672 21876
rect 16623 21845 16635 21848
rect 16577 21839 16635 21845
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 17604 21876 17632 21907
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 18233 21947 18291 21953
rect 17736 21916 17781 21944
rect 17736 21904 17742 21916
rect 18233 21913 18245 21947
rect 18279 21944 18291 21947
rect 18322 21944 18328 21956
rect 18279 21916 18328 21944
rect 18279 21913 18291 21916
rect 18233 21907 18291 21913
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 19306 21944 19334 21984
rect 19720 21984 20668 22012
rect 19720 21944 19748 21984
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 21177 22015 21235 22021
rect 20772 21984 20817 22012
rect 20772 21972 20778 21984
rect 21177 21981 21189 22015
rect 21223 21981 21235 22015
rect 21177 21975 21235 21981
rect 19306 21916 19748 21944
rect 20622 21904 20628 21956
rect 20680 21944 20686 21956
rect 21192 21944 21220 21975
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22097 22015 22155 22021
rect 22097 22012 22109 22015
rect 22060 21984 22109 22012
rect 22060 21972 22066 21984
rect 22097 21981 22109 21984
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 24486 22012 24492 22024
rect 23063 21984 24492 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 22186 21944 22192 21956
rect 20680 21916 22192 21944
rect 20680 21904 20686 21916
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 22848 21944 22876 21975
rect 24486 21972 24492 21984
rect 24544 21972 24550 22024
rect 24578 21972 24584 22024
rect 24636 22012 24642 22024
rect 24636 21984 24681 22012
rect 24636 21972 24642 21984
rect 24854 21972 24860 22024
rect 24912 22012 24918 22024
rect 26329 22015 26387 22021
rect 26329 22012 26341 22015
rect 24912 21984 26341 22012
rect 24912 21972 24918 21984
rect 26329 21981 26341 21984
rect 26375 21981 26387 22015
rect 26329 21975 26387 21981
rect 31665 22015 31723 22021
rect 31665 21981 31677 22015
rect 31711 22012 31723 22015
rect 38286 22012 38292 22024
rect 31711 21984 35894 22012
rect 38247 21984 38292 22012
rect 31711 21981 31723 21984
rect 31665 21975 31723 21981
rect 22848 21916 23612 21944
rect 19426 21876 19432 21888
rect 17604 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21876 19490 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 19484 21848 20085 21876
rect 19484 21836 19490 21848
rect 20073 21845 20085 21848
rect 20119 21845 20131 21879
rect 20530 21876 20536 21888
rect 20491 21848 20536 21876
rect 20073 21839 20131 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 20898 21836 20904 21888
rect 20956 21876 20962 21888
rect 21269 21879 21327 21885
rect 21269 21876 21281 21879
rect 20956 21848 21281 21876
rect 20956 21836 20962 21848
rect 21269 21845 21281 21848
rect 21315 21845 21327 21879
rect 21269 21839 21327 21845
rect 21913 21879 21971 21885
rect 21913 21845 21925 21879
rect 21959 21876 21971 21879
rect 22462 21876 22468 21888
rect 21959 21848 22468 21876
rect 21959 21845 21971 21848
rect 21913 21839 21971 21845
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 23106 21836 23112 21888
rect 23164 21876 23170 21888
rect 23477 21879 23535 21885
rect 23477 21876 23489 21879
rect 23164 21848 23489 21876
rect 23164 21836 23170 21848
rect 23477 21845 23489 21848
rect 23523 21845 23535 21879
rect 23584 21876 23612 21916
rect 23658 21904 23664 21956
rect 23716 21944 23722 21956
rect 25685 21947 25743 21953
rect 25685 21944 25697 21947
rect 23716 21916 25697 21944
rect 23716 21904 23722 21916
rect 25685 21913 25697 21916
rect 25731 21913 25743 21947
rect 31846 21944 31852 21956
rect 31807 21916 31852 21944
rect 25685 21907 25743 21913
rect 31846 21904 31852 21916
rect 31904 21904 31910 21956
rect 25130 21876 25136 21888
rect 23584 21848 25136 21876
rect 23477 21839 23535 21845
rect 25130 21836 25136 21848
rect 25188 21836 25194 21888
rect 35866 21876 35894 21984
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 35866 21848 38117 21876
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1360 21644 3096 21672
rect 1360 21632 1366 21644
rect 2682 21604 2688 21616
rect 2643 21576 2688 21604
rect 2682 21564 2688 21576
rect 2740 21564 2746 21616
rect 3068 21604 3096 21644
rect 3694 21632 3700 21684
rect 3752 21672 3758 21684
rect 3752 21644 5304 21672
rect 3752 21632 3758 21644
rect 5276 21604 5304 21644
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 6178 21672 6184 21684
rect 5408 21644 6184 21672
rect 5408 21632 5414 21644
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 6549 21675 6607 21681
rect 6549 21641 6561 21675
rect 6595 21672 6607 21675
rect 7742 21672 7748 21684
rect 6595 21644 7748 21672
rect 6595 21641 6607 21644
rect 6549 21635 6607 21641
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 7834 21632 7840 21684
rect 7892 21672 7898 21684
rect 12069 21675 12127 21681
rect 7892 21644 11100 21672
rect 7892 21632 7898 21644
rect 8754 21604 8760 21616
rect 3068 21576 3174 21604
rect 5276 21576 8760 21604
rect 8754 21564 8760 21576
rect 8812 21564 8818 21616
rect 10410 21604 10416 21616
rect 9982 21576 10416 21604
rect 10410 21564 10416 21576
rect 10468 21564 10474 21616
rect 11072 21604 11100 21644
rect 12069 21641 12081 21675
rect 12115 21672 12127 21675
rect 12115 21644 14596 21672
rect 12115 21641 12127 21644
rect 12069 21635 12127 21641
rect 12434 21604 12440 21616
rect 11072 21576 12440 21604
rect 12434 21564 12440 21576
rect 12492 21564 12498 21616
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 13541 21607 13599 21613
rect 13541 21604 13553 21607
rect 13044 21576 13553 21604
rect 13044 21564 13050 21576
rect 13541 21573 13553 21576
rect 13587 21573 13599 21607
rect 14090 21604 14096 21616
rect 14051 21576 14096 21604
rect 13541 21567 13599 21573
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 1762 21536 1768 21548
rect 1723 21508 1768 21536
rect 1762 21496 1768 21508
rect 1820 21496 1826 21548
rect 5074 21536 5080 21548
rect 5035 21508 5080 21536
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 5718 21496 5724 21548
rect 5776 21536 5782 21548
rect 5813 21539 5871 21545
rect 5813 21536 5825 21539
rect 5776 21508 5825 21536
rect 5776 21496 5782 21508
rect 5813 21505 5825 21508
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21536 6791 21539
rect 6914 21536 6920 21548
rect 6779 21508 6920 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7377 21539 7435 21545
rect 7377 21505 7389 21539
rect 7423 21536 7435 21539
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7423 21508 7849 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 7837 21505 7849 21508
rect 7883 21536 7895 21539
rect 8110 21536 8116 21548
rect 7883 21508 8116 21536
rect 7883 21505 7895 21508
rect 7837 21499 7895 21505
rect 8110 21496 8116 21508
rect 8168 21496 8174 21548
rect 10962 21536 10968 21548
rect 10923 21508 10968 21536
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 14568 21545 14596 21644
rect 14642 21632 14648 21684
rect 14700 21672 14706 21684
rect 14700 21644 17356 21672
rect 14700 21632 14706 21644
rect 15010 21564 15016 21616
rect 15068 21604 15074 21616
rect 17218 21604 17224 21616
rect 15068 21576 15976 21604
rect 17179 21576 17224 21604
rect 15068 21564 15074 21576
rect 12897 21539 12955 21545
rect 12897 21536 12909 21539
rect 12676 21508 12909 21536
rect 12676 21496 12682 21508
rect 12897 21505 12909 21508
rect 12943 21505 12955 21539
rect 12897 21499 12955 21505
rect 14553 21539 14611 21545
rect 14553 21505 14565 21539
rect 14599 21505 14611 21539
rect 15838 21536 15844 21548
rect 15799 21508 15844 21536
rect 14553 21499 14611 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 1578 21428 1584 21480
rect 1636 21468 1642 21480
rect 2409 21471 2467 21477
rect 2409 21468 2421 21471
rect 1636 21440 2421 21468
rect 1636 21428 1642 21440
rect 2409 21437 2421 21440
rect 2455 21437 2467 21471
rect 4430 21468 4436 21480
rect 4343 21440 4436 21468
rect 2409 21431 2467 21437
rect 4430 21428 4436 21440
rect 4488 21468 4494 21480
rect 4890 21468 4896 21480
rect 4488 21440 4896 21468
rect 4488 21428 4494 21440
rect 4890 21428 4896 21440
rect 4948 21428 4954 21480
rect 8481 21471 8539 21477
rect 8481 21468 8493 21471
rect 6748 21440 8493 21468
rect 6748 21412 6776 21440
rect 8481 21437 8493 21440
rect 8527 21437 8539 21471
rect 8481 21431 8539 21437
rect 4614 21360 4620 21412
rect 4672 21400 4678 21412
rect 4672 21372 6684 21400
rect 4672 21360 4678 21372
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 1946 21332 1952 21344
rect 1627 21304 1952 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 1946 21292 1952 21304
rect 2004 21292 2010 21344
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 4893 21335 4951 21341
rect 4893 21332 4905 21335
rect 3108 21304 4905 21332
rect 3108 21292 3114 21304
rect 4893 21301 4905 21304
rect 4939 21301 4951 21335
rect 4893 21295 4951 21301
rect 5905 21335 5963 21341
rect 5905 21301 5917 21335
rect 5951 21332 5963 21335
rect 6362 21332 6368 21344
rect 5951 21304 6368 21332
rect 5951 21301 5963 21304
rect 5905 21295 5963 21301
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 6656 21332 6684 21372
rect 6730 21360 6736 21412
rect 6788 21360 6794 21412
rect 7193 21335 7251 21341
rect 7193 21332 7205 21335
rect 6656 21304 7205 21332
rect 7193 21301 7205 21304
rect 7239 21301 7251 21335
rect 7193 21295 7251 21301
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 7929 21335 7987 21341
rect 7929 21332 7941 21335
rect 7892 21304 7941 21332
rect 7892 21292 7898 21304
rect 7929 21301 7941 21304
rect 7975 21301 7987 21335
rect 8496 21332 8524 21431
rect 8754 21428 8760 21480
rect 8812 21468 8818 21480
rect 9766 21468 9772 21480
rect 8812 21440 9772 21468
rect 8812 21428 8818 21440
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 10502 21428 10508 21480
rect 10560 21468 10566 21480
rect 13449 21471 13507 21477
rect 10560 21440 13400 21468
rect 10560 21428 10566 21440
rect 11057 21403 11115 21409
rect 11057 21369 11069 21403
rect 11103 21400 11115 21403
rect 12894 21400 12900 21412
rect 11103 21372 12900 21400
rect 11103 21369 11115 21372
rect 11057 21363 11115 21369
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 13372 21400 13400 21440
rect 13449 21437 13461 21471
rect 13495 21468 13507 21471
rect 14182 21468 14188 21480
rect 13495 21440 14188 21468
rect 13495 21437 13507 21440
rect 13449 21431 13507 21437
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 14734 21468 14740 21480
rect 14695 21440 14740 21468
rect 14734 21428 14740 21440
rect 14792 21428 14798 21480
rect 15657 21471 15715 21477
rect 15657 21437 15669 21471
rect 15703 21468 15715 21471
rect 15746 21468 15752 21480
rect 15703 21440 15752 21468
rect 15703 21437 15715 21440
rect 15657 21431 15715 21437
rect 15746 21428 15752 21440
rect 15804 21428 15810 21480
rect 15948 21468 15976 21576
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 17328 21604 17356 21644
rect 17678 21632 17684 21684
rect 17736 21672 17742 21684
rect 18509 21675 18567 21681
rect 18509 21672 18521 21675
rect 17736 21644 18521 21672
rect 17736 21632 17742 21644
rect 18509 21641 18521 21644
rect 18555 21641 18567 21675
rect 22002 21672 22008 21684
rect 18509 21635 18567 21641
rect 18616 21644 21772 21672
rect 21963 21644 22008 21672
rect 18616 21604 18644 21644
rect 20530 21604 20536 21616
rect 17328 21576 18644 21604
rect 18708 21576 20536 21604
rect 18708 21545 18736 21576
rect 20530 21564 20536 21576
rect 20588 21564 20594 21616
rect 20898 21604 20904 21616
rect 20859 21576 20904 21604
rect 20898 21564 20904 21576
rect 20956 21564 20962 21616
rect 21453 21607 21511 21613
rect 21453 21573 21465 21607
rect 21499 21604 21511 21607
rect 21634 21604 21640 21616
rect 21499 21576 21640 21604
rect 21499 21573 21511 21576
rect 21453 21567 21511 21573
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 21744 21604 21772 21644
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22649 21675 22707 21681
rect 22649 21641 22661 21675
rect 22695 21672 22707 21675
rect 23474 21672 23480 21684
rect 22695 21644 23480 21672
rect 22695 21641 22707 21644
rect 22649 21635 22707 21641
rect 23474 21632 23480 21644
rect 23532 21632 23538 21684
rect 25317 21675 25375 21681
rect 25317 21672 25329 21675
rect 23676 21644 25329 21672
rect 23676 21613 23704 21644
rect 25317 21641 25329 21644
rect 25363 21641 25375 21675
rect 33778 21672 33784 21684
rect 33739 21644 33784 21672
rect 25317 21635 25375 21641
rect 33778 21632 33784 21644
rect 33836 21632 33842 21684
rect 23661 21607 23719 21613
rect 21744 21576 22094 21604
rect 22066 21548 22094 21576
rect 23661 21573 23673 21607
rect 23707 21573 23719 21607
rect 24210 21604 24216 21616
rect 24171 21576 24216 21604
rect 23661 21567 23719 21573
rect 24210 21564 24216 21576
rect 24268 21564 24274 21616
rect 24486 21564 24492 21616
rect 24544 21604 24550 21616
rect 24765 21607 24823 21613
rect 24765 21604 24777 21607
rect 24544 21576 24777 21604
rect 24544 21564 24550 21576
rect 24765 21573 24777 21576
rect 24811 21573 24823 21607
rect 24765 21567 24823 21573
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 19245 21539 19303 21545
rect 19245 21505 19257 21539
rect 19291 21536 19303 21539
rect 19334 21536 19340 21548
rect 19291 21508 19340 21536
rect 19291 21505 19303 21508
rect 19245 21499 19303 21505
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 19978 21496 19984 21548
rect 20036 21536 20042 21548
rect 20073 21539 20131 21545
rect 20073 21536 20085 21539
rect 20036 21508 20085 21536
rect 20036 21496 20042 21508
rect 20073 21505 20085 21508
rect 20119 21536 20131 21539
rect 20438 21536 20444 21548
rect 20119 21508 20444 21536
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 22066 21536 22100 21548
rect 22007 21508 22100 21536
rect 22094 21496 22100 21508
rect 22152 21536 22158 21548
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 22152 21508 22201 21536
rect 22152 21496 22158 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 17129 21471 17187 21477
rect 17129 21468 17141 21471
rect 15948 21440 17141 21468
rect 17129 21437 17141 21440
rect 17175 21437 17187 21471
rect 20622 21468 20628 21480
rect 17129 21431 17187 21437
rect 17604 21440 20628 21468
rect 17604 21400 17632 21440
rect 20622 21428 20628 21440
rect 20680 21428 20686 21480
rect 20809 21471 20867 21477
rect 20809 21437 20821 21471
rect 20855 21468 20867 21471
rect 20898 21468 20904 21480
rect 20855 21440 20904 21468
rect 20855 21437 20867 21440
rect 20809 21431 20867 21437
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 22848 21468 22876 21499
rect 24578 21496 24584 21548
rect 24636 21536 24642 21548
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 24636 21508 24685 21536
rect 24636 21496 24642 21508
rect 24673 21505 24685 21508
rect 24719 21536 24731 21539
rect 25222 21536 25228 21548
rect 24719 21508 25228 21536
rect 24719 21505 24731 21508
rect 24673 21499 24731 21505
rect 25222 21496 25228 21508
rect 25280 21496 25286 21548
rect 25498 21536 25504 21548
rect 25459 21508 25504 21536
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 26145 21539 26203 21545
rect 26145 21505 26157 21539
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 33689 21539 33747 21545
rect 33689 21505 33701 21539
rect 33735 21536 33747 21539
rect 38102 21536 38108 21548
rect 33735 21508 38108 21536
rect 33735 21505 33747 21508
rect 33689 21499 33747 21505
rect 21324 21440 22876 21468
rect 23569 21471 23627 21477
rect 21324 21428 21330 21440
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 23658 21468 23664 21480
rect 23615 21440 23664 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 24854 21428 24860 21480
rect 24912 21468 24918 21480
rect 26160 21468 26188 21499
rect 38102 21496 38108 21508
rect 38160 21496 38166 21548
rect 24912 21440 26188 21468
rect 24912 21428 24918 21440
rect 13372 21372 17632 21400
rect 17681 21403 17739 21409
rect 17681 21369 17693 21403
rect 17727 21400 17739 21403
rect 18138 21400 18144 21412
rect 17727 21372 18144 21400
rect 17727 21369 17739 21372
rect 17681 21363 17739 21369
rect 18138 21360 18144 21372
rect 18196 21360 18202 21412
rect 19337 21403 19395 21409
rect 19337 21369 19349 21403
rect 19383 21400 19395 21403
rect 19426 21400 19432 21412
rect 19383 21372 19432 21400
rect 19383 21369 19395 21372
rect 19337 21363 19395 21369
rect 19426 21360 19432 21372
rect 19484 21360 19490 21412
rect 9766 21332 9772 21344
rect 8496 21304 9772 21332
rect 7929 21295 7987 21301
rect 9766 21292 9772 21304
rect 9824 21332 9830 21344
rect 9950 21332 9956 21344
rect 9824 21304 9956 21332
rect 9824 21292 9830 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10229 21335 10287 21341
rect 10229 21301 10241 21335
rect 10275 21332 10287 21335
rect 10502 21332 10508 21344
rect 10275 21304 10508 21332
rect 10275 21301 10287 21304
rect 10229 21295 10287 21301
rect 10502 21292 10508 21304
rect 10560 21292 10566 21344
rect 12713 21335 12771 21341
rect 12713 21301 12725 21335
rect 12759 21332 12771 21335
rect 14550 21332 14556 21344
rect 12759 21304 14556 21332
rect 12759 21301 12771 21304
rect 12713 21295 12771 21301
rect 14550 21292 14556 21304
rect 14608 21292 14614 21344
rect 14826 21292 14832 21344
rect 14884 21332 14890 21344
rect 14921 21335 14979 21341
rect 14921 21332 14933 21335
rect 14884 21304 14933 21332
rect 14884 21292 14890 21304
rect 14921 21301 14933 21304
rect 14967 21301 14979 21335
rect 14921 21295 14979 21301
rect 15194 21292 15200 21344
rect 15252 21332 15258 21344
rect 16025 21335 16083 21341
rect 16025 21332 16037 21335
rect 15252 21304 16037 21332
rect 15252 21292 15258 21304
rect 16025 21301 16037 21304
rect 16071 21332 16083 21335
rect 16390 21332 16396 21344
rect 16071 21304 16396 21332
rect 16071 21301 16083 21304
rect 16025 21295 16083 21301
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 20165 21335 20223 21341
rect 20165 21301 20177 21335
rect 20211 21332 20223 21335
rect 20438 21332 20444 21344
rect 20211 21304 20444 21332
rect 20211 21301 20223 21304
rect 20165 21295 20223 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 20530 21292 20536 21344
rect 20588 21332 20594 21344
rect 25590 21332 25596 21344
rect 20588 21304 25596 21332
rect 20588 21292 20594 21304
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 25958 21332 25964 21344
rect 25919 21304 25964 21332
rect 25958 21292 25964 21304
rect 26016 21292 26022 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 4236 21131 4294 21137
rect 4236 21097 4248 21131
rect 4282 21128 4294 21131
rect 5902 21128 5908 21140
rect 4282 21100 5908 21128
rect 4282 21097 4294 21100
rect 4236 21091 4294 21097
rect 5902 21088 5908 21100
rect 5960 21088 5966 21140
rect 9858 21128 9864 21140
rect 6932 21100 9864 21128
rect 3973 20995 4031 21001
rect 3973 20992 3985 20995
rect 1596 20964 3985 20992
rect 1596 20936 1624 20964
rect 3973 20961 3985 20964
rect 4019 20992 4031 20995
rect 4246 20992 4252 21004
rect 4019 20964 4252 20992
rect 4019 20961 4031 20964
rect 3973 20955 4031 20961
rect 4246 20952 4252 20964
rect 4304 20952 4310 21004
rect 5997 20995 6055 21001
rect 5997 20961 6009 20995
rect 6043 20992 6055 20995
rect 6932 20992 6960 21100
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 10318 21088 10324 21140
rect 10376 21128 10382 21140
rect 11977 21131 12035 21137
rect 11977 21128 11989 21131
rect 10376 21100 11989 21128
rect 10376 21088 10382 21100
rect 11977 21097 11989 21100
rect 12023 21097 12035 21131
rect 11977 21091 12035 21097
rect 16390 21088 16396 21140
rect 16448 21128 16454 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 16448 21100 16681 21128
rect 16448 21088 16454 21100
rect 16669 21097 16681 21100
rect 16715 21097 16727 21131
rect 16669 21091 16727 21097
rect 16758 21088 16764 21140
rect 16816 21128 16822 21140
rect 20530 21128 20536 21140
rect 16816 21100 20536 21128
rect 16816 21088 16822 21100
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 22741 21131 22799 21137
rect 22741 21097 22753 21131
rect 22787 21128 22799 21131
rect 25498 21128 25504 21140
rect 22787 21100 25504 21128
rect 22787 21097 22799 21100
rect 22741 21091 22799 21097
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 25590 21088 25596 21140
rect 25648 21128 25654 21140
rect 27893 21131 27951 21137
rect 25648 21100 26234 21128
rect 25648 21088 25654 21100
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 8573 21063 8631 21069
rect 8573 21060 8585 21063
rect 8536 21032 8585 21060
rect 8536 21020 8542 21032
rect 8573 21029 8585 21032
rect 8619 21029 8631 21063
rect 8573 21023 8631 21029
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 9585 21063 9643 21069
rect 9585 21060 9597 21063
rect 9364 21032 9597 21060
rect 9364 21020 9370 21032
rect 9585 21029 9597 21032
rect 9631 21029 9643 21063
rect 14826 21060 14832 21072
rect 14787 21032 14832 21060
rect 9585 21023 9643 21029
rect 14826 21020 14832 21032
rect 14884 21020 14890 21072
rect 15102 21020 15108 21072
rect 15160 21060 15166 21072
rect 19978 21060 19984 21072
rect 15160 21032 19984 21060
rect 15160 21020 15166 21032
rect 19978 21020 19984 21032
rect 20036 21020 20042 21072
rect 25958 21060 25964 21072
rect 23584 21032 25964 21060
rect 6043 20964 6960 20992
rect 7101 20995 7159 21001
rect 6043 20961 6055 20964
rect 5997 20955 6055 20961
rect 7101 20961 7113 20995
rect 7147 20992 7159 20995
rect 7190 20992 7196 21004
rect 7147 20964 7196 20992
rect 7147 20961 7159 20964
rect 7101 20955 7159 20961
rect 7190 20952 7196 20964
rect 7248 20952 7254 21004
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 9950 20992 9956 21004
rect 8168 20964 9956 20992
rect 8168 20952 8174 20964
rect 9950 20952 9956 20964
rect 10008 20952 10014 21004
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 10502 20992 10508 21004
rect 10284 20964 10329 20992
rect 10463 20964 10508 20992
rect 10284 20952 10290 20964
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 10594 20952 10600 21004
rect 10652 20992 10658 21004
rect 12805 20995 12863 21001
rect 10652 20964 12664 20992
rect 10652 20952 10658 20964
rect 1578 20924 1584 20936
rect 1539 20896 1584 20924
rect 1578 20884 1584 20896
rect 1636 20884 1642 20936
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6788 20896 6837 20924
rect 6788 20884 6794 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 8478 20884 8484 20936
rect 8536 20924 8542 20936
rect 9769 20927 9827 20933
rect 8536 20896 9720 20924
rect 8536 20884 8542 20896
rect 1857 20859 1915 20865
rect 1857 20825 1869 20859
rect 1903 20825 1915 20859
rect 1857 20819 1915 20825
rect 1872 20788 1900 20819
rect 2866 20816 2872 20868
rect 2924 20816 2930 20868
rect 3602 20856 3608 20868
rect 3160 20828 3608 20856
rect 3160 20788 3188 20828
rect 3602 20816 3608 20828
rect 3660 20816 3666 20868
rect 5258 20816 5264 20868
rect 5316 20816 5322 20868
rect 7558 20816 7564 20868
rect 7616 20816 7622 20868
rect 9692 20856 9720 20896
rect 9769 20893 9781 20927
rect 9815 20924 9827 20927
rect 10042 20924 10048 20936
rect 9815 20896 10048 20924
rect 9815 20893 9827 20896
rect 9769 20887 9827 20893
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 10594 20856 10600 20868
rect 8404 20828 9628 20856
rect 9692 20828 10600 20856
rect 1872 20760 3188 20788
rect 3329 20791 3387 20797
rect 3329 20757 3341 20791
rect 3375 20788 3387 20791
rect 4154 20788 4160 20800
rect 3375 20760 4160 20788
rect 3375 20757 3387 20760
rect 3329 20751 3387 20757
rect 4154 20748 4160 20760
rect 4212 20748 4218 20800
rect 4890 20748 4896 20800
rect 4948 20788 4954 20800
rect 8404 20788 8432 20828
rect 4948 20760 8432 20788
rect 9600 20788 9628 20828
rect 10594 20816 10600 20828
rect 10652 20816 10658 20868
rect 11054 20816 11060 20868
rect 11112 20816 11118 20868
rect 11790 20788 11796 20800
rect 9600 20760 11796 20788
rect 4948 20748 4954 20760
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 12636 20788 12664 20964
rect 12805 20961 12817 20995
rect 12851 20992 12863 20995
rect 13262 20992 13268 21004
rect 12851 20964 13268 20992
rect 12851 20961 12863 20964
rect 12805 20955 12863 20961
rect 13262 20952 13268 20964
rect 13320 20952 13326 21004
rect 13446 20992 13452 21004
rect 13407 20964 13452 20992
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 14461 20995 14519 21001
rect 14461 20961 14473 20995
rect 14507 20992 14519 20995
rect 14918 20992 14924 21004
rect 14507 20964 14924 20992
rect 14507 20961 14519 20964
rect 14461 20955 14519 20961
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20992 16543 20995
rect 16666 20992 16672 21004
rect 16531 20964 16672 20992
rect 16531 20961 16543 20964
rect 16485 20955 16543 20961
rect 16666 20952 16672 20964
rect 16724 20952 16730 21004
rect 19334 20992 19340 21004
rect 16776 20964 19340 20992
rect 14642 20924 14648 20936
rect 14603 20896 14648 20924
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20924 15899 20927
rect 15930 20924 15936 20936
rect 15887 20896 15936 20924
rect 15887 20893 15899 20896
rect 15841 20887 15899 20893
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16298 20924 16304 20936
rect 16259 20896 16304 20924
rect 16298 20884 16304 20896
rect 16356 20884 16362 20936
rect 12894 20816 12900 20868
rect 12952 20856 12958 20868
rect 16776 20856 16804 20964
rect 19334 20952 19340 20964
rect 19392 20992 19398 21004
rect 20070 20992 20076 21004
rect 19392 20964 20076 20992
rect 19392 20952 19398 20964
rect 20070 20952 20076 20964
rect 20128 20952 20134 21004
rect 20438 20992 20444 21004
rect 20399 20964 20444 20992
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 23584 21001 23612 21032
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 26206 21060 26234 21100
rect 27893 21097 27905 21131
rect 27939 21128 27951 21131
rect 31754 21128 31760 21140
rect 27939 21100 31760 21128
rect 27939 21097 27951 21100
rect 27893 21091 27951 21097
rect 31754 21088 31760 21100
rect 31812 21088 31818 21140
rect 38102 21128 38108 21140
rect 38063 21100 38108 21128
rect 38102 21088 38108 21100
rect 38160 21088 38166 21140
rect 30466 21060 30472 21072
rect 26206 21032 30472 21060
rect 30466 21020 30472 21032
rect 30524 21020 30530 21072
rect 23569 20995 23627 21001
rect 23569 20961 23581 20995
rect 23615 20961 23627 20995
rect 23569 20955 23627 20961
rect 24765 20995 24823 21001
rect 24765 20961 24777 20995
rect 24811 20992 24823 20995
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 24811 20964 27169 20992
rect 24811 20961 24823 20964
rect 24765 20955 24823 20961
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 18564 20896 19625 20924
rect 18564 20884 18570 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20924 20315 20927
rect 20806 20924 20812 20936
rect 20303 20896 20812 20924
rect 20303 20893 20315 20896
rect 20257 20887 20315 20893
rect 20806 20884 20812 20896
rect 20864 20884 20870 20936
rect 21542 20924 21548 20936
rect 21503 20896 21548 20924
rect 21542 20884 21548 20896
rect 21600 20884 21606 20936
rect 22278 20924 22284 20936
rect 22239 20896 22284 20924
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 22738 20884 22744 20936
rect 22796 20924 22802 20936
rect 22925 20927 22983 20933
rect 22925 20924 22937 20927
rect 22796 20896 22937 20924
rect 22796 20884 22802 20896
rect 22925 20893 22937 20896
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23385 20927 23443 20933
rect 23385 20893 23397 20927
rect 23431 20924 23443 20927
rect 24670 20924 24676 20936
rect 23431 20896 24676 20924
rect 23431 20893 23443 20896
rect 23385 20887 23443 20893
rect 24670 20884 24676 20896
rect 24728 20884 24734 20936
rect 24949 20927 25007 20933
rect 24949 20893 24961 20927
rect 24995 20924 25007 20927
rect 25774 20924 25780 20936
rect 24995 20896 25780 20924
rect 24995 20893 25007 20896
rect 24949 20887 25007 20893
rect 25774 20884 25780 20896
rect 25832 20884 25838 20936
rect 25866 20884 25872 20936
rect 25924 20924 25930 20936
rect 26697 20927 26755 20933
rect 26697 20924 26709 20927
rect 25924 20896 26709 20924
rect 25924 20884 25930 20896
rect 26697 20893 26709 20896
rect 26743 20893 26755 20927
rect 27798 20924 27804 20936
rect 27759 20896 27804 20924
rect 26697 20887 26755 20893
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 38286 20924 38292 20936
rect 38247 20896 38292 20924
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 17678 20856 17684 20868
rect 12952 20828 12997 20856
rect 13096 20828 16804 20856
rect 17639 20828 17684 20856
rect 12952 20816 12958 20828
rect 13096 20788 13124 20828
rect 17678 20816 17684 20828
rect 17736 20816 17742 20868
rect 17773 20859 17831 20865
rect 17773 20825 17785 20859
rect 17819 20856 17831 20859
rect 18046 20856 18052 20868
rect 17819 20828 18052 20856
rect 17819 20825 17831 20828
rect 17773 20819 17831 20825
rect 18046 20816 18052 20828
rect 18104 20816 18110 20868
rect 18138 20816 18144 20868
rect 18196 20856 18202 20868
rect 18325 20859 18383 20865
rect 18325 20856 18337 20859
rect 18196 20828 18337 20856
rect 18196 20816 18202 20828
rect 18325 20825 18337 20828
rect 18371 20825 18383 20859
rect 35526 20856 35532 20868
rect 18325 20819 18383 20825
rect 19306 20828 35532 20856
rect 12636 20760 13124 20788
rect 15286 20748 15292 20800
rect 15344 20788 15350 20800
rect 15657 20791 15715 20797
rect 15657 20788 15669 20791
rect 15344 20760 15669 20788
rect 15344 20748 15350 20760
rect 15657 20757 15669 20760
rect 15703 20757 15715 20791
rect 15657 20751 15715 20757
rect 15746 20748 15752 20800
rect 15804 20788 15810 20800
rect 16758 20788 16764 20800
rect 15804 20760 16764 20788
rect 15804 20748 15810 20760
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 18340 20788 18368 20819
rect 19306 20788 19334 20828
rect 35526 20816 35532 20828
rect 35584 20816 35590 20868
rect 19426 20788 19432 20800
rect 18340 20760 19334 20788
rect 19387 20760 19432 20788
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 20898 20788 20904 20800
rect 20859 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 21358 20788 21364 20800
rect 21319 20760 21364 20788
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20788 22155 20791
rect 22462 20788 22468 20800
rect 22143 20760 22468 20788
rect 22143 20757 22155 20760
rect 22097 20751 22155 20757
rect 22462 20748 22468 20760
rect 22520 20748 22526 20800
rect 24026 20788 24032 20800
rect 23987 20760 24032 20788
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 25406 20788 25412 20800
rect 25367 20760 25412 20788
rect 25406 20748 25412 20760
rect 25464 20748 25470 20800
rect 25958 20788 25964 20800
rect 25919 20760 25964 20788
rect 25958 20748 25964 20760
rect 26016 20748 26022 20800
rect 26510 20788 26516 20800
rect 26471 20760 26516 20788
rect 26510 20748 26516 20760
rect 26568 20748 26574 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 11146 20584 11152 20596
rect 1872 20556 3556 20584
rect 1872 20525 1900 20556
rect 1857 20519 1915 20525
rect 1857 20485 1869 20519
rect 1903 20485 1915 20519
rect 3234 20516 3240 20528
rect 3082 20488 3240 20516
rect 1857 20479 1915 20485
rect 3234 20476 3240 20488
rect 3292 20476 3298 20528
rect 1578 20380 1584 20392
rect 1539 20352 1584 20380
rect 1578 20340 1584 20352
rect 1636 20340 1642 20392
rect 3528 20380 3556 20556
rect 3712 20556 11008 20584
rect 11107 20556 11152 20584
rect 3602 20408 3608 20460
rect 3660 20448 3666 20460
rect 3712 20448 3740 20556
rect 4522 20516 4528 20528
rect 4483 20488 4528 20516
rect 4522 20476 4528 20488
rect 4580 20476 4586 20528
rect 5534 20476 5540 20528
rect 5592 20476 5598 20528
rect 7558 20476 7564 20528
rect 7616 20476 7622 20528
rect 9766 20516 9772 20528
rect 9416 20488 9772 20516
rect 4246 20448 4252 20460
rect 3660 20420 3753 20448
rect 4207 20420 4252 20448
rect 3660 20408 3666 20420
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 9416 20457 9444 20488
rect 9766 20476 9772 20488
rect 9824 20476 9830 20528
rect 10980 20516 11008 20556
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 11698 20584 11704 20596
rect 11388 20556 11704 20584
rect 11388 20544 11394 20556
rect 11698 20544 11704 20556
rect 11756 20584 11762 20596
rect 12526 20584 12532 20596
rect 11756 20556 12532 20584
rect 11756 20544 11762 20556
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 13909 20587 13967 20593
rect 13909 20553 13921 20587
rect 13955 20584 13967 20587
rect 16945 20587 17003 20593
rect 13955 20556 15424 20584
rect 13955 20553 13967 20556
rect 13909 20547 13967 20553
rect 10980 20488 12434 20516
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20417 9459 20451
rect 9401 20411 9459 20417
rect 10778 20408 10784 20460
rect 10836 20408 10842 20460
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 3528 20352 5580 20380
rect 5552 20312 5580 20352
rect 5902 20340 5908 20392
rect 5960 20380 5966 20392
rect 6730 20380 6736 20392
rect 5960 20352 6736 20380
rect 5960 20340 5966 20352
rect 6730 20340 6736 20352
rect 6788 20340 6794 20392
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7558 20380 7564 20392
rect 7055 20352 7564 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7558 20340 7564 20352
rect 7616 20340 7622 20392
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20380 8539 20383
rect 8570 20380 8576 20392
rect 8527 20352 8576 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9677 20383 9735 20389
rect 9677 20380 9689 20383
rect 9180 20352 9689 20380
rect 9180 20340 9186 20352
rect 9677 20349 9689 20352
rect 9723 20349 9735 20383
rect 9677 20343 9735 20349
rect 10042 20340 10048 20392
rect 10100 20380 10106 20392
rect 12176 20380 12204 20411
rect 10100 20352 12204 20380
rect 10100 20340 10106 20352
rect 12406 20324 12434 20488
rect 12618 20476 12624 20528
rect 12676 20516 12682 20528
rect 13357 20519 13415 20525
rect 12676 20488 13308 20516
rect 12676 20476 12682 20488
rect 13280 20457 13308 20488
rect 13357 20485 13369 20519
rect 13403 20516 13415 20519
rect 14642 20516 14648 20528
rect 13403 20488 14648 20516
rect 13403 20485 13415 20488
rect 13357 20479 13415 20485
rect 14642 20476 14648 20488
rect 14700 20476 14706 20528
rect 15286 20516 15292 20528
rect 14752 20488 15292 20516
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20448 13323 20451
rect 13538 20448 13544 20460
rect 13311 20420 13544 20448
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 12820 20380 12848 20411
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 14752 20457 14780 20488
rect 15286 20476 15292 20488
rect 15344 20476 15350 20528
rect 15396 20525 15424 20556
rect 16945 20553 16957 20587
rect 16991 20584 17003 20587
rect 17678 20584 17684 20596
rect 16991 20556 17684 20584
rect 16991 20553 17003 20556
rect 16945 20547 17003 20553
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 18046 20544 18052 20596
rect 18104 20584 18110 20596
rect 18785 20587 18843 20593
rect 18785 20584 18797 20587
rect 18104 20556 18797 20584
rect 18104 20544 18110 20556
rect 18785 20553 18797 20556
rect 18831 20553 18843 20587
rect 18785 20547 18843 20553
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 22278 20584 22284 20596
rect 22143 20556 22284 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 23661 20587 23719 20593
rect 23661 20553 23673 20587
rect 23707 20584 23719 20587
rect 24854 20584 24860 20596
rect 23707 20556 24860 20584
rect 23707 20553 23719 20556
rect 23661 20547 23719 20553
rect 24854 20544 24860 20556
rect 24912 20544 24918 20596
rect 25406 20584 25412 20596
rect 25367 20556 25412 20584
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 25869 20587 25927 20593
rect 25869 20584 25881 20587
rect 25832 20556 25881 20584
rect 25832 20544 25838 20556
rect 25869 20553 25881 20556
rect 25915 20553 25927 20587
rect 25869 20547 25927 20553
rect 15381 20519 15439 20525
rect 15381 20485 15393 20519
rect 15427 20485 15439 20519
rect 15381 20479 15439 20485
rect 17773 20519 17831 20525
rect 17773 20485 17785 20519
rect 17819 20516 17831 20519
rect 18138 20516 18144 20528
rect 17819 20488 18144 20516
rect 17819 20485 17831 20488
rect 17773 20479 17831 20485
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 18322 20516 18328 20528
rect 18283 20488 18328 20516
rect 18322 20476 18328 20488
rect 18380 20476 18386 20528
rect 20070 20476 20076 20528
rect 20128 20516 20134 20528
rect 20128 20488 23888 20516
rect 20128 20476 20134 20488
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14737 20451 14795 20457
rect 14139 20420 14688 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14366 20380 14372 20392
rect 12820 20352 14372 20380
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 12250 20312 12256 20324
rect 5552 20284 6040 20312
rect 4246 20204 4252 20256
rect 4304 20244 4310 20256
rect 5074 20244 5080 20256
rect 4304 20216 5080 20244
rect 4304 20204 4310 20216
rect 5074 20204 5080 20216
rect 5132 20244 5138 20256
rect 5902 20244 5908 20256
rect 5132 20216 5908 20244
rect 5132 20204 5138 20216
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 6012 20253 6040 20284
rect 8036 20284 8616 20312
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 8036 20244 8064 20284
rect 6043 20216 8064 20244
rect 8588 20244 8616 20284
rect 10704 20284 12256 20312
rect 10704 20244 10732 20284
rect 12250 20272 12256 20284
rect 12308 20272 12314 20324
rect 12406 20284 12440 20324
rect 12434 20272 12440 20284
rect 12492 20272 12498 20324
rect 13722 20312 13728 20324
rect 12544 20284 13728 20312
rect 8588 20216 10732 20244
rect 11977 20247 12035 20253
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 11977 20213 11989 20247
rect 12023 20244 12035 20247
rect 12544 20244 12572 20284
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 14660 20312 14688 20420
rect 14737 20417 14749 20451
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20448 19027 20451
rect 19426 20448 19432 20460
rect 19015 20420 19432 20448
rect 19015 20417 19027 20420
rect 18969 20411 19027 20417
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 19978 20408 19984 20460
rect 20036 20448 20042 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 20036 20420 20177 20448
rect 20036 20408 20042 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20809 20451 20867 20457
rect 20809 20417 20821 20451
rect 20855 20448 20867 20451
rect 21358 20448 21364 20460
rect 20855 20420 21364 20448
rect 20855 20417 20867 20420
rect 20809 20411 20867 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20448 22339 20451
rect 22370 20448 22376 20460
rect 22327 20420 22376 20448
rect 22327 20417 22339 20420
rect 22281 20411 22339 20417
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 22738 20448 22744 20460
rect 22699 20420 22744 20448
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 23860 20457 23888 20488
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20448 23903 20451
rect 24118 20448 24124 20460
rect 23891 20420 24124 20448
rect 23891 20417 23903 20420
rect 23845 20411 23903 20417
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24670 20408 24676 20460
rect 24728 20448 24734 20460
rect 24765 20451 24823 20457
rect 24765 20448 24777 20451
rect 24728 20420 24777 20448
rect 24728 20408 24734 20420
rect 24765 20417 24777 20420
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 24949 20451 25007 20457
rect 24949 20417 24961 20451
rect 24995 20448 25007 20451
rect 25958 20448 25964 20460
rect 24995 20420 25964 20448
rect 24995 20417 25007 20420
rect 24949 20411 25007 20417
rect 25958 20408 25964 20420
rect 26016 20408 26022 20460
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26510 20448 26516 20460
rect 26099 20420 26516 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26510 20408 26516 20420
rect 26568 20408 26574 20460
rect 15289 20383 15347 20389
rect 15289 20349 15301 20383
rect 15335 20380 15347 20383
rect 15470 20380 15476 20392
rect 15335 20352 15476 20380
rect 15335 20349 15347 20352
rect 15289 20343 15347 20349
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 15562 20340 15568 20392
rect 15620 20380 15626 20392
rect 17681 20383 17739 20389
rect 15620 20352 15665 20380
rect 15620 20340 15626 20352
rect 17681 20349 17693 20383
rect 17727 20349 17739 20383
rect 17681 20343 17739 20349
rect 16022 20312 16028 20324
rect 14660 20284 16028 20312
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 17696 20312 17724 20343
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 18012 20352 20637 20380
rect 18012 20340 18018 20352
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 24026 20312 24032 20324
rect 17696 20284 24032 20312
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 12023 20216 12572 20244
rect 12621 20247 12679 20253
rect 12023 20213 12035 20216
rect 11977 20207 12035 20213
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 14458 20244 14464 20256
rect 12667 20216 14464 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 14553 20247 14611 20253
rect 14553 20213 14565 20247
rect 14599 20244 14611 20247
rect 15378 20244 15384 20256
rect 14599 20216 15384 20244
rect 14599 20213 14611 20216
rect 14553 20207 14611 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 19981 20247 20039 20253
rect 19981 20213 19993 20247
rect 20027 20244 20039 20247
rect 20530 20244 20536 20256
rect 20027 20216 20536 20244
rect 20027 20213 20039 20216
rect 19981 20207 20039 20213
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 21269 20247 21327 20253
rect 21269 20213 21281 20247
rect 21315 20244 21327 20247
rect 22186 20244 22192 20256
rect 21315 20216 22192 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 22278 20204 22284 20256
rect 22336 20244 22342 20256
rect 22833 20247 22891 20253
rect 22833 20244 22845 20247
rect 22336 20216 22845 20244
rect 22336 20204 22342 20216
rect 22833 20213 22845 20216
rect 22879 20213 22891 20247
rect 22833 20207 22891 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 4522 20000 4528 20052
rect 4580 20040 4586 20052
rect 4890 20040 4896 20052
rect 4580 20012 4896 20040
rect 4580 20000 4586 20012
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 6825 20043 6883 20049
rect 6825 20009 6837 20043
rect 6871 20040 6883 20043
rect 7190 20040 7196 20052
rect 6871 20012 7196 20040
rect 6871 20009 6883 20012
rect 6825 20003 6883 20009
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 11974 20040 11980 20052
rect 9171 20012 11980 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 14553 20043 14611 20049
rect 12406 20012 13308 20040
rect 8294 19972 8300 19984
rect 8255 19944 8300 19972
rect 8294 19932 8300 19944
rect 8352 19932 8358 19984
rect 9766 19932 9772 19984
rect 9824 19932 9830 19984
rect 9861 19975 9919 19981
rect 9861 19941 9873 19975
rect 9907 19972 9919 19975
rect 12406 19972 12434 20012
rect 9907 19944 10548 19972
rect 9907 19941 9919 19944
rect 9861 19935 9919 19941
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19904 1915 19907
rect 3786 19904 3792 19916
rect 1903 19876 3792 19904
rect 1903 19873 1915 19876
rect 1857 19867 1915 19873
rect 3786 19864 3792 19876
rect 3844 19864 3850 19916
rect 5074 19904 5080 19916
rect 5035 19876 5080 19904
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 5442 19864 5448 19916
rect 5500 19904 5506 19916
rect 8386 19904 8392 19916
rect 5500 19876 8392 19904
rect 5500 19864 5506 19876
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 9784 19904 9812 19932
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 9784 19876 10425 19904
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 10520 19904 10548 19944
rect 11716 19944 12434 19972
rect 11716 19904 11744 19944
rect 13280 19913 13308 20012
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 14734 20040 14740 20052
rect 14599 20012 14740 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 17497 20043 17555 20049
rect 17497 20040 17509 20043
rect 17276 20012 17509 20040
rect 17276 20000 17282 20012
rect 17497 20009 17509 20012
rect 17543 20009 17555 20043
rect 18138 20040 18144 20052
rect 18099 20012 18144 20040
rect 17497 20003 17555 20009
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21542 20040 21548 20052
rect 21131 20012 21548 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 31846 20040 31852 20052
rect 23348 20012 31852 20040
rect 23348 20000 23354 20012
rect 31846 20000 31852 20012
rect 31904 20000 31910 20052
rect 15194 19972 15200 19984
rect 13556 19944 15200 19972
rect 13265 19907 13323 19913
rect 10520 19876 11744 19904
rect 11992 19876 13216 19904
rect 10413 19867 10471 19873
rect 1578 19836 1584 19848
rect 1539 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 4614 19836 4620 19848
rect 4575 19808 4620 19836
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 9306 19836 9312 19848
rect 9267 19808 9312 19836
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19836 9827 19839
rect 10134 19836 10140 19848
rect 9815 19808 10140 19836
rect 9815 19805 9827 19808
rect 9769 19799 9827 19805
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 3142 19768 3148 19780
rect 3082 19740 3148 19768
rect 3142 19728 3148 19740
rect 3200 19728 3206 19780
rect 5074 19768 5080 19780
rect 3344 19740 5080 19768
rect 3234 19660 3240 19712
rect 3292 19700 3298 19712
rect 3344 19709 3372 19740
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 5353 19771 5411 19777
rect 5353 19737 5365 19771
rect 5399 19768 5411 19771
rect 5626 19768 5632 19780
rect 5399 19740 5632 19768
rect 5399 19737 5411 19740
rect 5353 19731 5411 19737
rect 5626 19728 5632 19740
rect 5684 19728 5690 19780
rect 5902 19728 5908 19780
rect 5960 19728 5966 19780
rect 7745 19771 7803 19777
rect 7745 19737 7757 19771
rect 7791 19737 7803 19771
rect 7745 19731 7803 19737
rect 3329 19703 3387 19709
rect 3329 19700 3341 19703
rect 3292 19672 3341 19700
rect 3292 19660 3298 19672
rect 3329 19669 3341 19672
rect 3375 19669 3387 19703
rect 3329 19663 3387 19669
rect 4433 19703 4491 19709
rect 4433 19669 4445 19703
rect 4479 19700 4491 19703
rect 6730 19700 6736 19712
rect 4479 19672 6736 19700
rect 4479 19669 4491 19672
rect 4433 19663 4491 19669
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 7760 19700 7788 19731
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 7892 19740 7937 19768
rect 7892 19728 7898 19740
rect 8018 19728 8024 19780
rect 8076 19768 8082 19780
rect 10594 19768 10600 19780
rect 8076 19740 10600 19768
rect 8076 19728 8082 19740
rect 10594 19728 10600 19740
rect 10652 19728 10658 19780
rect 10689 19771 10747 19777
rect 10689 19737 10701 19771
rect 10735 19768 10747 19771
rect 10962 19768 10968 19780
rect 10735 19740 10968 19768
rect 10735 19737 10747 19740
rect 10689 19731 10747 19737
rect 10962 19728 10968 19740
rect 11020 19728 11026 19780
rect 11422 19728 11428 19780
rect 11480 19728 11486 19780
rect 11992 19700 12020 19876
rect 13078 19836 13084 19848
rect 13039 19808 13084 19836
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13188 19836 13216 19876
rect 13265 19873 13277 19907
rect 13311 19873 13323 19907
rect 13265 19867 13323 19873
rect 13556 19836 13584 19944
rect 15194 19932 15200 19944
rect 15252 19932 15258 19984
rect 15562 19972 15568 19984
rect 15523 19944 15568 19972
rect 15562 19932 15568 19944
rect 15620 19972 15626 19984
rect 16669 19975 16727 19981
rect 16669 19972 16681 19975
rect 15620 19944 16681 19972
rect 15620 19932 15626 19944
rect 16669 19941 16681 19944
rect 16715 19941 16727 19975
rect 18506 19972 18512 19984
rect 16669 19935 16727 19941
rect 17972 19944 18512 19972
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15436 19876 15481 19904
rect 15436 19864 15442 19876
rect 16206 19864 16212 19916
rect 16264 19904 16270 19916
rect 16485 19907 16543 19913
rect 16485 19904 16497 19907
rect 16264 19876 16497 19904
rect 16264 19864 16270 19876
rect 16485 19873 16497 19876
rect 16531 19873 16543 19907
rect 16485 19867 16543 19873
rect 13188 19808 13584 19836
rect 14550 19796 14556 19848
rect 14608 19836 14614 19848
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 14608 19808 14749 19836
rect 14608 19796 14614 19808
rect 14737 19805 14749 19808
rect 14783 19805 14795 19839
rect 14737 19799 14795 19805
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19836 15255 19839
rect 15746 19836 15752 19848
rect 15243 19808 15752 19836
rect 15243 19805 15255 19808
rect 15197 19799 15255 19805
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 16298 19836 16304 19848
rect 16259 19808 16304 19836
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 17402 19836 17408 19848
rect 17315 19808 17408 19836
rect 17402 19796 17408 19808
rect 17460 19836 17466 19848
rect 17972 19836 18000 19944
rect 18506 19932 18512 19944
rect 18564 19932 18570 19984
rect 22370 19972 22376 19984
rect 21284 19944 22376 19972
rect 19242 19864 19248 19916
rect 19300 19904 19306 19916
rect 20714 19904 20720 19916
rect 19300 19876 20720 19904
rect 19300 19864 19306 19876
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 17460 19808 18000 19836
rect 18049 19839 18107 19845
rect 17460 19796 17466 19808
rect 18049 19805 18061 19839
rect 18095 19832 18107 19839
rect 18138 19832 18144 19848
rect 18095 19805 18144 19832
rect 18049 19804 18144 19805
rect 18049 19799 18107 19804
rect 18138 19796 18144 19804
rect 18196 19796 18202 19848
rect 18874 19836 18880 19848
rect 18787 19808 18880 19836
rect 18874 19796 18880 19808
rect 18932 19836 18938 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 18932 19808 19441 19836
rect 18932 19796 18938 19808
rect 19429 19805 19441 19808
rect 19475 19836 19487 19839
rect 19978 19836 19984 19848
rect 19475 19808 19984 19836
rect 19475 19805 19487 19808
rect 19429 19799 19487 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20530 19836 20536 19848
rect 20491 19808 20536 19836
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 21284 19845 21312 19944
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 22922 19932 22928 19984
rect 22980 19972 22986 19984
rect 23661 19975 23719 19981
rect 23661 19972 23673 19975
rect 22980 19944 23673 19972
rect 22980 19932 22986 19944
rect 23661 19941 23673 19944
rect 23707 19941 23719 19975
rect 23661 19935 23719 19941
rect 24394 19932 24400 19984
rect 24452 19972 24458 19984
rect 25593 19975 25651 19981
rect 25593 19972 25605 19975
rect 24452 19944 25605 19972
rect 24452 19932 24458 19944
rect 25593 19941 25605 19944
rect 25639 19941 25651 19975
rect 25593 19935 25651 19941
rect 22833 19907 22891 19913
rect 22833 19873 22845 19907
rect 22879 19904 22891 19907
rect 24210 19904 24216 19916
rect 22879 19876 24216 19904
rect 22879 19873 22891 19876
rect 22833 19867 22891 19873
rect 24210 19864 24216 19876
rect 24268 19864 24274 19916
rect 25041 19907 25099 19913
rect 25041 19873 25053 19907
rect 25087 19904 25099 19907
rect 25406 19904 25412 19916
rect 25087 19876 25412 19904
rect 25087 19873 25099 19876
rect 25041 19867 25099 19873
rect 25406 19864 25412 19876
rect 25464 19864 25470 19916
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 23290 19836 23296 19848
rect 23251 19808 23296 19836
rect 21269 19799 21327 19805
rect 12434 19728 12440 19780
rect 12492 19768 12498 19780
rect 21284 19768 21312 19799
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19836 23535 19839
rect 24670 19836 24676 19848
rect 23523 19808 24676 19836
rect 23523 19805 23535 19808
rect 23477 19799 23535 19805
rect 24670 19796 24676 19808
rect 24728 19796 24734 19848
rect 26326 19836 26332 19848
rect 26287 19808 26332 19836
rect 26326 19796 26332 19808
rect 26384 19796 26390 19848
rect 12492 19740 21312 19768
rect 12492 19728 12498 19740
rect 21542 19728 21548 19780
rect 21600 19768 21606 19780
rect 22189 19771 22247 19777
rect 22189 19768 22201 19771
rect 21600 19740 22201 19768
rect 21600 19728 21606 19740
rect 22189 19737 22201 19740
rect 22235 19737 22247 19771
rect 22189 19731 22247 19737
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 25130 19768 25136 19780
rect 22336 19740 22381 19768
rect 25091 19740 25136 19768
rect 22336 19728 22342 19740
rect 25130 19728 25136 19740
rect 25188 19728 25194 19780
rect 7760 19672 12020 19700
rect 12161 19703 12219 19709
rect 12161 19669 12173 19703
rect 12207 19700 12219 19703
rect 12250 19700 12256 19712
rect 12207 19672 12256 19700
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 13814 19700 13820 19712
rect 13771 19672 13820 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 13814 19660 13820 19672
rect 13872 19700 13878 19712
rect 15010 19700 15016 19712
rect 13872 19672 15016 19700
rect 13872 19660 13878 19672
rect 15010 19660 15016 19672
rect 15068 19660 15074 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 18414 19700 18420 19712
rect 15160 19672 18420 19700
rect 15160 19660 15166 19672
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 18690 19700 18696 19712
rect 18651 19672 18696 19700
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19334 19660 19340 19712
rect 19392 19700 19398 19712
rect 19521 19703 19579 19709
rect 19521 19700 19533 19703
rect 19392 19672 19533 19700
rect 19392 19660 19398 19672
rect 19521 19669 19533 19672
rect 19567 19669 19579 19703
rect 20346 19700 20352 19712
rect 20307 19672 20352 19700
rect 19521 19663 19579 19669
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 26050 19660 26056 19712
rect 26108 19700 26114 19712
rect 26145 19703 26203 19709
rect 26145 19700 26157 19703
rect 26108 19672 26157 19700
rect 26108 19660 26114 19672
rect 26145 19669 26157 19672
rect 26191 19669 26203 19703
rect 26145 19663 26203 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 4709 19499 4767 19505
rect 4709 19465 4721 19499
rect 4755 19496 4767 19499
rect 5442 19496 5448 19508
rect 4755 19468 5448 19496
rect 4755 19465 4767 19468
rect 4709 19459 4767 19465
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 5994 19456 6000 19508
rect 6052 19496 6058 19508
rect 8757 19499 8815 19505
rect 6052 19468 6592 19496
rect 6052 19456 6058 19468
rect 3786 19428 3792 19440
rect 3747 19400 3792 19428
rect 3786 19388 3792 19400
rect 3844 19388 3850 19440
rect 6564 19428 6592 19468
rect 8757 19465 8769 19499
rect 8803 19496 8815 19499
rect 11882 19496 11888 19508
rect 8803 19468 11888 19496
rect 8803 19465 8815 19468
rect 8757 19459 8815 19465
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 13814 19496 13820 19508
rect 12483 19468 13820 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 16390 19496 16396 19508
rect 14108 19468 16396 19496
rect 6733 19431 6791 19437
rect 6733 19428 6745 19431
rect 6564 19400 6745 19428
rect 6733 19397 6745 19400
rect 6779 19397 6791 19431
rect 6733 19391 6791 19397
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 8113 19431 8171 19437
rect 6972 19400 7328 19428
rect 6972 19388 6978 19400
rect 3142 19320 3148 19372
rect 3200 19320 3206 19372
rect 4890 19320 4896 19372
rect 4948 19360 4954 19372
rect 5997 19363 6055 19369
rect 4948 19332 4993 19360
rect 4948 19320 4954 19332
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 6270 19360 6276 19372
rect 6043 19332 6276 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 7300 19360 7328 19400
rect 8113 19397 8125 19431
rect 8159 19428 8171 19431
rect 9306 19428 9312 19440
rect 8159 19400 9312 19428
rect 8159 19397 8171 19400
rect 8113 19391 8171 19397
rect 9306 19388 9312 19400
rect 9364 19388 9370 19440
rect 9766 19428 9772 19440
rect 9416 19400 9772 19428
rect 9416 19369 9444 19400
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 14108 19428 14136 19468
rect 16390 19456 16396 19468
rect 16448 19496 16454 19508
rect 17954 19496 17960 19508
rect 16448 19468 17960 19496
rect 16448 19456 16454 19468
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 20349 19499 20407 19505
rect 20349 19465 20361 19499
rect 20395 19496 20407 19499
rect 20898 19496 20904 19508
rect 20395 19468 20904 19496
rect 20395 19465 20407 19468
rect 20349 19459 20407 19465
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 22922 19496 22928 19508
rect 22883 19468 22928 19496
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 24670 19496 24676 19508
rect 23400 19468 23704 19496
rect 24631 19468 24676 19496
rect 12676 19400 14136 19428
rect 12676 19388 12682 19400
rect 14182 19388 14188 19440
rect 14240 19428 14246 19440
rect 14369 19431 14427 19437
rect 14369 19428 14381 19431
rect 14240 19400 14381 19428
rect 14240 19388 14246 19400
rect 14369 19397 14381 19400
rect 14415 19397 14427 19431
rect 14369 19391 14427 19397
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 21453 19431 21511 19437
rect 16356 19400 18552 19428
rect 16356 19388 16362 19400
rect 8941 19363 8999 19369
rect 8941 19360 8953 19363
rect 7300 19332 8953 19360
rect 8941 19329 8953 19332
rect 8987 19329 8999 19363
rect 8941 19323 8999 19329
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19329 9459 19363
rect 9401 19323 9459 19329
rect 10778 19320 10784 19372
rect 10836 19320 10842 19372
rect 11790 19360 11796 19372
rect 11751 19332 11796 19360
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12308 19332 12664 19360
rect 12308 19320 12314 19332
rect 1578 19252 1584 19304
rect 1636 19292 1642 19304
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1636 19264 1777 19292
rect 1636 19252 1642 19264
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 3326 19292 3332 19304
rect 2087 19264 3332 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 3326 19252 3332 19264
rect 3384 19252 3390 19304
rect 4706 19252 4712 19304
rect 4764 19252 4770 19304
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19292 5411 19295
rect 5442 19292 5448 19304
rect 5399 19264 5448 19292
rect 5399 19261 5411 19264
rect 5353 19255 5411 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 5537 19295 5595 19301
rect 5537 19261 5549 19295
rect 5583 19261 5595 19295
rect 5537 19255 5595 19261
rect 4724 19224 4752 19252
rect 5552 19224 5580 19255
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6696 19264 6741 19292
rect 6696 19252 6702 19264
rect 7558 19252 7564 19304
rect 7616 19292 7622 19304
rect 7616 19264 10732 19292
rect 7616 19252 7622 19264
rect 4724 19196 5580 19224
rect 6546 19184 6552 19236
rect 6604 19224 6610 19236
rect 7193 19227 7251 19233
rect 7193 19224 7205 19227
rect 6604 19196 7205 19224
rect 6604 19184 6610 19196
rect 7193 19193 7205 19196
rect 7239 19193 7251 19227
rect 7193 19187 7251 19193
rect 7926 19184 7932 19236
rect 7984 19224 7990 19236
rect 9030 19224 9036 19236
rect 7984 19196 9036 19224
rect 7984 19184 7990 19196
rect 9030 19184 9036 19196
rect 9088 19224 9094 19236
rect 10704 19224 10732 19264
rect 10870 19252 10876 19304
rect 10928 19292 10934 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 10928 19264 11161 19292
rect 10928 19252 10934 19264
rect 11149 19261 11161 19264
rect 11195 19261 11207 19295
rect 11974 19292 11980 19304
rect 11935 19264 11980 19292
rect 11149 19255 11207 19261
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12342 19224 12348 19236
rect 9088 19196 9536 19224
rect 10704 19196 12348 19224
rect 9088 19184 9094 19196
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4890 19156 4896 19168
rect 4212 19128 4896 19156
rect 4212 19116 4218 19128
rect 4890 19116 4896 19128
rect 4948 19156 4954 19168
rect 9122 19156 9128 19168
rect 4948 19128 9128 19156
rect 4948 19116 4954 19128
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 9508 19156 9536 19196
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 12636 19224 12664 19332
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12768 19332 13093 19360
rect 12768 19320 12774 19332
rect 13081 19329 13093 19332
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19360 13231 19363
rect 15194 19360 15200 19372
rect 13219 19332 15200 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13096 19292 13124 19323
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 17862 19360 17868 19372
rect 16899 19332 17868 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 18524 19369 18552 19400
rect 21453 19397 21465 19431
rect 21499 19428 21511 19431
rect 21542 19428 21548 19440
rect 21499 19400 21548 19428
rect 21499 19397 21511 19400
rect 21453 19391 21511 19397
rect 21542 19388 21548 19400
rect 21600 19388 21606 19440
rect 23400 19428 23428 19468
rect 23566 19428 23572 19440
rect 22066 19400 23428 19428
rect 23527 19400 23572 19428
rect 18509 19363 18567 19369
rect 18509 19329 18521 19363
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20346 19360 20352 19372
rect 19935 19332 20352 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 13354 19292 13360 19304
rect 13096 19264 13360 19292
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13630 19252 13636 19304
rect 13688 19292 13694 19304
rect 13725 19295 13783 19301
rect 13725 19292 13737 19295
rect 13688 19264 13737 19292
rect 13688 19252 13694 19264
rect 13725 19261 13737 19264
rect 13771 19261 13783 19295
rect 13725 19255 13783 19261
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 13909 19295 13967 19301
rect 13909 19292 13921 19295
rect 13872 19264 13921 19292
rect 13872 19252 13878 19264
rect 13909 19261 13921 19264
rect 13955 19261 13967 19295
rect 13909 19255 13967 19261
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14516 19264 15056 19292
rect 14516 19252 14522 19264
rect 14918 19224 14924 19236
rect 12636 19196 14924 19224
rect 14918 19184 14924 19196
rect 14976 19184 14982 19236
rect 15028 19224 15056 19264
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15289 19295 15347 19301
rect 15160 19264 15205 19292
rect 15160 19252 15166 19264
rect 15289 19261 15301 19295
rect 15335 19261 15347 19295
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 15289 19255 15347 19261
rect 15304 19224 15332 19255
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 17368 19264 17509 19292
rect 17368 19252 17374 19264
rect 17497 19261 17509 19264
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19292 18751 19295
rect 19334 19292 19340 19304
rect 18739 19264 19340 19292
rect 18739 19261 18751 19264
rect 18693 19255 18751 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19720 19292 19748 19323
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 22066 19360 22094 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 23676 19428 23704 19468
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 25130 19456 25136 19508
rect 25188 19496 25194 19508
rect 25869 19499 25927 19505
rect 25869 19496 25881 19499
rect 25188 19468 25881 19496
rect 25188 19456 25194 19468
rect 25869 19465 25881 19468
rect 25915 19465 25927 19499
rect 25869 19459 25927 19465
rect 34054 19428 34060 19440
rect 23676 19400 34060 19428
rect 34054 19388 34060 19400
rect 34112 19388 34118 19440
rect 20855 19332 22094 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 22186 19320 22192 19372
rect 22244 19360 22250 19372
rect 22830 19360 22836 19372
rect 22244 19332 22836 19360
rect 22244 19320 22250 19332
rect 22830 19320 22836 19332
rect 22888 19360 22894 19372
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 22888 19332 23336 19360
rect 22888 19320 22894 19332
rect 20254 19292 20260 19304
rect 19720 19264 20260 19292
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19292 21051 19295
rect 21266 19292 21272 19304
rect 21039 19264 21272 19292
rect 21039 19261 21051 19264
rect 20993 19255 21051 19261
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 22278 19292 22284 19304
rect 22239 19264 22284 19292
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 22462 19292 22468 19304
rect 22423 19264 22468 19292
rect 22462 19252 22468 19264
rect 22520 19252 22526 19304
rect 23308 19292 23336 19332
rect 24136 19332 24593 19360
rect 23477 19295 23535 19301
rect 23477 19292 23489 19295
rect 23308 19264 23489 19292
rect 23477 19261 23489 19264
rect 23523 19261 23535 19295
rect 24136 19292 24164 19332
rect 24581 19329 24593 19332
rect 24627 19329 24639 19363
rect 25406 19360 25412 19372
rect 25367 19332 25412 19360
rect 24581 19323 24639 19329
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 26050 19360 26056 19372
rect 26011 19332 26056 19360
rect 26050 19320 26056 19332
rect 26108 19320 26114 19372
rect 23477 19255 23535 19261
rect 23860 19264 24164 19292
rect 15470 19224 15476 19236
rect 15028 19196 15332 19224
rect 15431 19196 15476 19224
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 22738 19224 22744 19236
rect 15580 19196 22744 19224
rect 9658 19159 9716 19165
rect 9658 19156 9670 19159
rect 9508 19128 9670 19156
rect 9658 19125 9670 19128
rect 9704 19125 9716 19159
rect 9658 19119 9716 19125
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 12066 19156 12072 19168
rect 11112 19128 12072 19156
rect 11112 19116 11118 19128
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 15580 19156 15608 19196
rect 22738 19184 22744 19196
rect 22796 19184 22802 19236
rect 23860 19224 23888 19264
rect 23400 19196 23888 19224
rect 12216 19128 15608 19156
rect 12216 19116 12222 19128
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 19058 19156 19064 19168
rect 16356 19128 19064 19156
rect 16356 19116 16362 19128
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 19153 19159 19211 19165
rect 19153 19125 19165 19159
rect 19199 19156 19211 19159
rect 19242 19156 19248 19168
rect 19199 19128 19248 19156
rect 19199 19125 19211 19128
rect 19153 19119 19211 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 23400 19156 23428 19196
rect 23934 19184 23940 19236
rect 23992 19224 23998 19236
rect 24029 19227 24087 19233
rect 24029 19224 24041 19227
rect 23992 19196 24041 19224
rect 23992 19184 23998 19196
rect 24029 19193 24041 19196
rect 24075 19224 24087 19227
rect 27522 19224 27528 19236
rect 24075 19196 27528 19224
rect 24075 19193 24087 19196
rect 24029 19187 24087 19193
rect 27522 19184 27528 19196
rect 27580 19184 27586 19236
rect 25222 19156 25228 19168
rect 22428 19128 23428 19156
rect 25183 19128 25228 19156
rect 22428 19116 22434 19128
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 3326 18952 3332 18964
rect 3239 18924 3332 18952
rect 3326 18912 3332 18924
rect 3384 18952 3390 18964
rect 9677 18955 9735 18961
rect 3384 18924 8432 18952
rect 3384 18912 3390 18924
rect 5721 18887 5779 18893
rect 5721 18853 5733 18887
rect 5767 18884 5779 18887
rect 7558 18884 7564 18896
rect 5767 18856 7564 18884
rect 5767 18853 5779 18856
rect 5721 18847 5779 18853
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 8205 18887 8263 18893
rect 8205 18853 8217 18887
rect 8251 18884 8263 18887
rect 8294 18884 8300 18896
rect 8251 18856 8300 18884
rect 8251 18853 8263 18856
rect 8205 18847 8263 18853
rect 8294 18844 8300 18856
rect 8352 18844 8358 18896
rect 8404 18884 8432 18924
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 10042 18952 10048 18964
rect 9723 18924 10048 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 10042 18912 10048 18924
rect 10100 18912 10106 18964
rect 13725 18955 13783 18961
rect 13725 18921 13737 18955
rect 13771 18952 13783 18955
rect 13906 18952 13912 18964
rect 13771 18924 13912 18952
rect 13771 18921 13783 18924
rect 13725 18915 13783 18921
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14424 18924 14473 18952
rect 14424 18912 14430 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 14461 18915 14519 18921
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15654 18912 15660 18964
rect 15712 18952 15718 18964
rect 18046 18952 18052 18964
rect 15712 18924 18052 18952
rect 15712 18912 15718 18924
rect 18046 18912 18052 18924
rect 18104 18952 18110 18964
rect 30006 18952 30012 18964
rect 18104 18924 30012 18952
rect 18104 18912 18110 18924
rect 30006 18912 30012 18924
rect 30064 18912 30070 18964
rect 12066 18884 12072 18896
rect 8404 18856 10456 18884
rect 12027 18856 12072 18884
rect 3973 18819 4031 18825
rect 3973 18816 3985 18819
rect 1596 18788 3985 18816
rect 1596 18760 1624 18788
rect 3973 18785 3985 18788
rect 4019 18785 4031 18819
rect 3973 18779 4031 18785
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18816 4307 18819
rect 4890 18816 4896 18828
rect 4295 18788 4896 18816
rect 4295 18785 4307 18788
rect 4249 18779 4307 18785
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18816 7711 18819
rect 8938 18816 8944 18828
rect 7699 18788 8944 18816
rect 7699 18785 7711 18788
rect 7653 18779 7711 18785
rect 8938 18776 8944 18788
rect 8996 18776 9002 18828
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 9824 18788 10333 18816
rect 9824 18776 9830 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10428 18816 10456 18856
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 23934 18884 23940 18896
rect 13004 18856 23796 18884
rect 23895 18856 23940 18884
rect 10428 18788 11928 18816
rect 10321 18779 10379 18785
rect 1578 18748 1584 18760
rect 1539 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 6914 18748 6920 18760
rect 5868 18720 6920 18748
rect 5868 18708 5874 18720
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7190 18748 7196 18760
rect 7147 18720 7196 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 8352 18720 9873 18748
rect 8352 18708 8358 18720
rect 9861 18717 9873 18720
rect 9907 18748 9919 18751
rect 10134 18748 10140 18760
rect 9907 18720 10140 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 1964 18652 2346 18680
rect 1210 18572 1216 18624
rect 1268 18612 1274 18624
rect 1964 18612 1992 18652
rect 4982 18640 4988 18692
rect 5040 18640 5046 18692
rect 6273 18683 6331 18689
rect 6273 18649 6285 18683
rect 6319 18680 6331 18683
rect 6638 18680 6644 18692
rect 6319 18652 6644 18680
rect 6319 18649 6331 18652
rect 6273 18643 6331 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 6730 18640 6736 18692
rect 6788 18680 6794 18692
rect 7738 18683 7796 18689
rect 6788 18652 7604 18680
rect 6788 18640 6794 18652
rect 6914 18612 6920 18624
rect 1268 18584 1992 18612
rect 6875 18584 6920 18612
rect 1268 18572 1274 18584
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7576 18612 7604 18652
rect 7738 18649 7750 18683
rect 7784 18649 7796 18683
rect 7738 18643 7796 18649
rect 7760 18612 7788 18643
rect 8570 18640 8576 18692
rect 8628 18680 8634 18692
rect 10318 18680 10324 18692
rect 8628 18652 10324 18680
rect 8628 18640 8634 18652
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 10594 18680 10600 18692
rect 10555 18652 10600 18680
rect 10594 18640 10600 18652
rect 10652 18640 10658 18692
rect 11606 18640 11612 18692
rect 11664 18640 11670 18692
rect 11900 18680 11928 18788
rect 13004 18748 13032 18856
rect 13081 18819 13139 18825
rect 13081 18785 13093 18819
rect 13127 18816 13139 18819
rect 13127 18788 15240 18816
rect 13127 18785 13139 18788
rect 13081 18779 13139 18785
rect 13265 18751 13323 18757
rect 13004 18720 13124 18748
rect 13096 18680 13124 18720
rect 13265 18717 13277 18751
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 11900 18652 13124 18680
rect 7576 18584 7788 18612
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 13280 18612 13308 18711
rect 13354 18708 13360 18760
rect 13412 18748 13418 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 13412 18720 14657 18748
rect 13412 18708 13418 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 15010 18708 15016 18760
rect 15068 18750 15074 18760
rect 15105 18751 15163 18757
rect 15105 18750 15117 18751
rect 15068 18722 15117 18750
rect 15068 18708 15074 18722
rect 15105 18717 15117 18722
rect 15151 18717 15163 18751
rect 15212 18748 15240 18788
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 17681 18819 17739 18825
rect 15344 18788 15389 18816
rect 15344 18776 15350 18788
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17727 18788 18429 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19116 18788 19441 18816
rect 19116 18776 19122 18788
rect 19429 18785 19441 18788
rect 19475 18816 19487 18819
rect 20070 18816 20076 18828
rect 19475 18788 20076 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 22278 18776 22284 18828
rect 22336 18816 22342 18828
rect 22373 18819 22431 18825
rect 22373 18816 22385 18819
rect 22336 18788 22385 18816
rect 22336 18776 22342 18788
rect 22373 18785 22385 18788
rect 22419 18785 22431 18819
rect 22373 18779 22431 18785
rect 22922 18776 22928 18828
rect 22980 18816 22986 18828
rect 23385 18819 23443 18825
rect 23385 18816 23397 18819
rect 22980 18788 23397 18816
rect 22980 18776 22986 18788
rect 23385 18785 23397 18788
rect 23431 18785 23443 18819
rect 23768 18816 23796 18856
rect 23934 18844 23940 18856
rect 23992 18844 23998 18896
rect 23768 18788 25268 18816
rect 23385 18779 23443 18785
rect 16298 18748 16304 18760
rect 15212 18720 16304 18748
rect 15105 18711 15163 18717
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17586 18748 17592 18760
rect 17547 18720 17592 18748
rect 17129 18711 17187 18717
rect 14274 18640 14280 18692
rect 14332 18680 14338 18692
rect 16850 18680 16856 18692
rect 14332 18652 16856 18680
rect 14332 18640 14338 18652
rect 16850 18640 16856 18652
rect 16908 18640 16914 18692
rect 17144 18680 17172 18711
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 18012 18720 18245 18748
rect 18012 18708 18018 18720
rect 18233 18717 18245 18720
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 19518 18708 19524 18760
rect 19576 18748 19582 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19576 18720 19625 18748
rect 19576 18708 19582 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18748 20591 18751
rect 22094 18748 22100 18760
rect 20579 18720 22100 18748
rect 20579 18717 20591 18720
rect 20533 18711 20591 18717
rect 22094 18708 22100 18720
rect 22152 18708 22158 18760
rect 24118 18708 24124 18760
rect 24176 18748 24182 18760
rect 25240 18757 25268 18788
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24176 18720 24593 18748
rect 24176 18708 24182 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18748 25283 18751
rect 26326 18748 26332 18760
rect 25271 18720 26332 18748
rect 25271 18717 25283 18720
rect 25225 18711 25283 18717
rect 26326 18708 26332 18720
rect 26384 18708 26390 18760
rect 18690 18680 18696 18692
rect 17144 18652 18696 18680
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 23474 18640 23480 18692
rect 23532 18680 23538 18692
rect 23532 18652 23577 18680
rect 23532 18640 23538 18652
rect 8904 18584 13308 18612
rect 8904 18572 8910 18584
rect 13354 18572 13360 18624
rect 13412 18612 13418 18624
rect 15654 18612 15660 18624
rect 13412 18584 15660 18612
rect 13412 18572 13418 18584
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 16298 18612 16304 18624
rect 16259 18584 16304 18612
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 16945 18615 17003 18621
rect 16945 18581 16957 18615
rect 16991 18612 17003 18615
rect 18138 18612 18144 18624
rect 16991 18584 18144 18612
rect 16991 18581 17003 18584
rect 16945 18575 17003 18581
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19150 18612 19156 18624
rect 18923 18584 19156 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 19150 18572 19156 18584
rect 19208 18612 19214 18624
rect 20073 18615 20131 18621
rect 20073 18612 20085 18615
rect 19208 18584 20085 18612
rect 19208 18572 19214 18584
rect 20073 18581 20085 18584
rect 20119 18581 20131 18615
rect 20622 18612 20628 18624
rect 20583 18584 20628 18612
rect 20073 18575 20131 18581
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 22922 18572 22928 18624
rect 22980 18612 22986 18624
rect 24673 18615 24731 18621
rect 24673 18612 24685 18615
rect 22980 18584 24685 18612
rect 22980 18572 22986 18584
rect 24673 18581 24685 18584
rect 24719 18581 24731 18615
rect 25314 18612 25320 18624
rect 25275 18584 25320 18612
rect 24673 18575 24731 18581
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1762 18408 1768 18420
rect 1723 18380 1768 18408
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 4798 18408 4804 18420
rect 2924 18380 4804 18408
rect 2924 18368 2930 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 6825 18411 6883 18417
rect 6825 18377 6837 18411
rect 6871 18408 6883 18411
rect 9122 18408 9128 18420
rect 6871 18380 9128 18408
rect 6871 18377 6883 18380
rect 6825 18371 6883 18377
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 9398 18368 9404 18420
rect 9456 18408 9462 18420
rect 9769 18411 9827 18417
rect 9769 18408 9781 18411
rect 9456 18380 9781 18408
rect 9456 18368 9462 18380
rect 9769 18377 9781 18380
rect 9815 18377 9827 18411
rect 9769 18371 9827 18377
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 16117 18411 16175 18417
rect 12216 18380 13308 18408
rect 12216 18368 12222 18380
rect 3329 18343 3387 18349
rect 3329 18309 3341 18343
rect 3375 18340 3387 18343
rect 6638 18340 6644 18352
rect 3375 18312 6644 18340
rect 3375 18309 3387 18312
rect 3329 18303 3387 18309
rect 6638 18300 6644 18312
rect 6696 18300 6702 18352
rect 7653 18343 7711 18349
rect 7653 18340 7665 18343
rect 7392 18312 7665 18340
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 2498 18272 2504 18284
rect 1627 18244 2504 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2498 18232 2504 18244
rect 2556 18232 2562 18284
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18272 3295 18275
rect 3602 18272 3608 18284
rect 3283 18244 3608 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 3602 18232 3608 18244
rect 3660 18232 3666 18284
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18241 3939 18275
rect 3881 18235 3939 18241
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18272 4767 18275
rect 4890 18272 4896 18284
rect 4755 18244 4896 18272
rect 4755 18241 4767 18244
rect 4709 18235 4767 18241
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18204 2651 18207
rect 3786 18204 3792 18216
rect 2639 18176 3792 18204
rect 2639 18173 2651 18176
rect 2593 18167 2651 18173
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 3896 18204 3924 18235
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 5626 18272 5632 18284
rect 5399 18244 5632 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 5368 18204 5396 18235
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 3896 18176 5396 18204
rect 3973 18139 4031 18145
rect 3973 18105 3985 18139
rect 4019 18136 4031 18139
rect 4982 18136 4988 18148
rect 4019 18108 4988 18136
rect 4019 18105 4031 18108
rect 3973 18099 4031 18105
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 5074 18096 5080 18148
rect 5132 18136 5138 18148
rect 5169 18139 5227 18145
rect 5169 18136 5181 18139
rect 5132 18108 5181 18136
rect 5132 18096 5138 18108
rect 5169 18105 5181 18108
rect 5215 18105 5227 18139
rect 5810 18136 5816 18148
rect 5771 18108 5816 18136
rect 5169 18099 5227 18105
rect 5810 18096 5816 18108
rect 5868 18096 5874 18148
rect 6012 18136 6040 18235
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6788 18244 7021 18272
rect 6788 18232 6794 18244
rect 7009 18241 7021 18244
rect 7055 18272 7067 18275
rect 7190 18272 7196 18284
rect 7055 18244 7196 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 7098 18164 7104 18216
rect 7156 18204 7162 18216
rect 7392 18204 7420 18312
rect 7653 18309 7665 18312
rect 7699 18309 7711 18343
rect 7653 18303 7711 18309
rect 7834 18300 7840 18352
rect 7892 18340 7898 18352
rect 7892 18312 9904 18340
rect 7892 18300 7898 18312
rect 9122 18232 9128 18284
rect 9180 18272 9186 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 9180 18244 9229 18272
rect 9180 18232 9186 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18272 9735 18275
rect 9766 18272 9772 18284
rect 9723 18244 9772 18272
rect 9723 18241 9735 18244
rect 9677 18235 9735 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 9876 18272 9904 18312
rect 10134 18300 10140 18352
rect 10192 18340 10198 18352
rect 10870 18340 10876 18352
rect 10192 18312 10876 18340
rect 10192 18300 10198 18312
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 11882 18340 11888 18352
rect 10980 18312 11284 18340
rect 11843 18312 11888 18340
rect 10321 18275 10379 18281
rect 10321 18272 10333 18275
rect 9876 18244 10333 18272
rect 10321 18241 10333 18244
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 10502 18232 10508 18284
rect 10560 18272 10566 18284
rect 10980 18272 11008 18312
rect 11146 18272 11152 18284
rect 10560 18244 11008 18272
rect 11107 18244 11152 18272
rect 10560 18232 10566 18244
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 11256 18272 11284 18312
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 13280 18281 13308 18380
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 17034 18408 17040 18420
rect 16163 18380 17040 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 21266 18408 21272 18420
rect 17184 18380 20760 18408
rect 21227 18380 21272 18408
rect 17184 18368 17190 18380
rect 14277 18343 14335 18349
rect 14277 18309 14289 18343
rect 14323 18340 14335 18343
rect 17678 18340 17684 18352
rect 14323 18312 17684 18340
rect 14323 18309 14335 18312
rect 14277 18303 14335 18309
rect 17678 18300 17684 18312
rect 17736 18300 17742 18352
rect 18046 18340 18052 18352
rect 17972 18312 18052 18340
rect 13265 18275 13323 18281
rect 11256 18244 11652 18272
rect 7156 18176 7420 18204
rect 7561 18207 7619 18213
rect 7156 18164 7162 18176
rect 7561 18173 7573 18207
rect 7607 18204 7619 18207
rect 10042 18204 10048 18216
rect 7607 18176 10048 18204
rect 7607 18173 7619 18176
rect 7561 18167 7619 18173
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 11624 18204 11652 18244
rect 13265 18241 13277 18275
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 13906 18232 13912 18284
rect 13964 18272 13970 18284
rect 15105 18275 15163 18281
rect 13964 18270 14964 18272
rect 15105 18270 15117 18275
rect 13964 18244 15117 18270
rect 13964 18232 13970 18244
rect 14936 18242 15117 18244
rect 15105 18241 15117 18242
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 15194 18232 15200 18284
rect 15252 18272 15258 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 15252 18244 15577 18272
rect 15252 18232 15258 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 16298 18272 16304 18284
rect 16259 18244 16304 18272
rect 15565 18235 15623 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 17972 18281 18000 18312
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 19150 18340 19156 18352
rect 19111 18312 19156 18340
rect 19150 18300 19156 18312
rect 19208 18300 19214 18352
rect 19245 18343 19303 18349
rect 19245 18309 19257 18343
rect 19291 18340 19303 18343
rect 20622 18340 20628 18352
rect 19291 18312 20628 18340
rect 19291 18309 19303 18312
rect 19245 18303 19303 18309
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 20732 18340 20760 18380
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 23566 18368 23572 18420
rect 23624 18408 23630 18420
rect 23937 18411 23995 18417
rect 23937 18408 23949 18411
rect 23624 18380 23949 18408
rect 23624 18368 23630 18380
rect 23937 18377 23949 18380
rect 23983 18377 23995 18411
rect 23937 18371 23995 18377
rect 24489 18411 24547 18417
rect 24489 18377 24501 18411
rect 24535 18377 24547 18411
rect 24489 18371 24547 18377
rect 20732 18312 23060 18340
rect 17957 18275 18015 18281
rect 16408 18244 17172 18272
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 10459 18176 11560 18204
rect 11624 18176 11805 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 8113 18139 8171 18145
rect 6012 18108 8064 18136
rect 4525 18071 4583 18077
rect 4525 18037 4537 18071
rect 4571 18068 4583 18071
rect 7650 18068 7656 18080
rect 4571 18040 7656 18068
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 8036 18068 8064 18108
rect 8113 18105 8125 18139
rect 8159 18136 8171 18139
rect 8202 18136 8208 18148
rect 8159 18108 8208 18136
rect 8159 18105 8171 18108
rect 8113 18099 8171 18105
rect 8202 18096 8208 18108
rect 8260 18096 8266 18148
rect 9033 18139 9091 18145
rect 9033 18105 9045 18139
rect 9079 18136 9091 18139
rect 11532 18136 11560 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 13078 18204 13084 18216
rect 13039 18176 13084 18204
rect 11793 18167 11851 18173
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13722 18164 13728 18216
rect 13780 18204 13786 18216
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 13780 18176 14933 18204
rect 13780 18164 13786 18176
rect 14921 18173 14933 18176
rect 14967 18204 14979 18207
rect 16408 18204 16436 18244
rect 16850 18204 16856 18216
rect 14967 18176 16436 18204
rect 16811 18176 16856 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 16850 18164 16856 18176
rect 16908 18164 16914 18216
rect 17034 18204 17040 18216
rect 16995 18176 17040 18204
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 17144 18204 17172 18244
rect 17957 18241 17969 18275
rect 18003 18241 18015 18275
rect 18138 18272 18144 18284
rect 18099 18244 18144 18272
rect 17957 18235 18015 18241
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 20956 18244 21189 18272
rect 20956 18232 20962 18244
rect 21177 18241 21189 18244
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18272 22155 18275
rect 22370 18272 22376 18284
rect 22143 18244 22376 18272
rect 22143 18241 22155 18244
rect 22097 18235 22155 18241
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 22922 18272 22928 18284
rect 22883 18244 22928 18272
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 23032 18272 23060 18312
rect 23474 18300 23480 18352
rect 23532 18340 23538 18352
rect 24504 18340 24532 18371
rect 25406 18340 25412 18352
rect 23532 18312 24532 18340
rect 24596 18312 25412 18340
rect 23532 18300 23538 18312
rect 23845 18275 23903 18281
rect 23845 18272 23857 18275
rect 23032 18244 23857 18272
rect 23845 18241 23857 18244
rect 23891 18272 23903 18275
rect 24596 18272 24624 18312
rect 25406 18300 25412 18312
rect 25464 18300 25470 18352
rect 23891 18244 24624 18272
rect 24673 18275 24731 18281
rect 23891 18241 23903 18244
rect 23845 18235 23903 18241
rect 24673 18241 24685 18275
rect 24719 18272 24731 18275
rect 25222 18272 25228 18284
rect 24719 18244 25228 18272
rect 24719 18241 24731 18244
rect 24673 18235 24731 18241
rect 25222 18232 25228 18244
rect 25280 18232 25286 18284
rect 20165 18207 20223 18213
rect 17144 18176 19334 18204
rect 12158 18136 12164 18148
rect 9079 18108 11468 18136
rect 11532 18108 12164 18136
rect 9079 18105 9091 18108
rect 9033 18099 9091 18105
rect 10502 18068 10508 18080
rect 8036 18040 10508 18068
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 10965 18071 11023 18077
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 11330 18068 11336 18080
rect 11011 18040 11336 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11440 18068 11468 18108
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 17126 18136 17132 18148
rect 12400 18108 17132 18136
rect 12400 18096 12406 18108
rect 17126 18096 17132 18108
rect 17184 18096 17190 18148
rect 19306 18136 19334 18176
rect 20165 18173 20177 18207
rect 20211 18204 20223 18207
rect 22646 18204 22652 18216
rect 20211 18176 22652 18204
rect 20211 18173 20223 18176
rect 20165 18167 20223 18173
rect 22646 18164 22652 18176
rect 22704 18164 22710 18216
rect 22741 18207 22799 18213
rect 22741 18173 22753 18207
rect 22787 18204 22799 18207
rect 23290 18204 23296 18216
rect 22787 18176 23296 18204
rect 22787 18173 22799 18176
rect 22741 18167 22799 18173
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 23385 18207 23443 18213
rect 23385 18173 23397 18207
rect 23431 18204 23443 18207
rect 24026 18204 24032 18216
rect 23431 18176 24032 18204
rect 23431 18173 23443 18176
rect 23385 18167 23443 18173
rect 24026 18164 24032 18176
rect 24084 18164 24090 18216
rect 20254 18136 20260 18148
rect 19306 18108 20260 18136
rect 20254 18096 20260 18108
rect 20312 18136 20318 18148
rect 20622 18136 20628 18148
rect 20312 18108 20628 18136
rect 20312 18096 20318 18108
rect 20622 18096 20628 18108
rect 20680 18096 20686 18148
rect 12618 18068 12624 18080
rect 11440 18040 12624 18068
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 13136 18040 13461 18068
rect 13136 18028 13142 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 13449 18031 13507 18037
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 18046 18068 18052 18080
rect 17543 18040 18052 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18601 18071 18659 18077
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 19242 18068 19248 18080
rect 18647 18040 19248 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 22189 18071 22247 18077
rect 22189 18037 22201 18071
rect 22235 18068 22247 18071
rect 22370 18068 22376 18080
rect 22235 18040 22376 18068
rect 22235 18037 22247 18040
rect 22189 18031 22247 18037
rect 22370 18028 22376 18040
rect 22428 18028 22434 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 7098 17864 7104 17876
rect 4724 17836 7104 17864
rect 2041 17799 2099 17805
rect 2041 17765 2053 17799
rect 2087 17796 2099 17799
rect 4430 17796 4436 17808
rect 2087 17768 4436 17796
rect 2087 17765 2099 17768
rect 2041 17759 2099 17765
rect 4430 17756 4436 17768
rect 4488 17756 4494 17808
rect 4525 17799 4583 17805
rect 4525 17765 4537 17799
rect 4571 17765 4583 17799
rect 4525 17759 4583 17765
rect 3694 17728 3700 17740
rect 2792 17700 3700 17728
rect 2792 17672 2820 17700
rect 3694 17688 3700 17700
rect 3752 17688 3758 17740
rect 1946 17660 1952 17672
rect 1907 17632 1952 17660
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2774 17660 2780 17672
rect 2735 17632 2780 17660
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 4540 17660 4568 17759
rect 4724 17669 4752 17836
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 9674 17864 9680 17876
rect 7668 17836 9680 17864
rect 5166 17756 5172 17808
rect 5224 17796 5230 17808
rect 5442 17796 5448 17808
rect 5224 17768 5448 17796
rect 5224 17756 5230 17768
rect 5442 17756 5448 17768
rect 5500 17756 5506 17808
rect 5813 17799 5871 17805
rect 5813 17765 5825 17799
rect 5859 17796 5871 17799
rect 6546 17796 6552 17808
rect 5859 17768 6552 17796
rect 5859 17765 5871 17768
rect 5813 17759 5871 17765
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 6454 17728 6460 17740
rect 5092 17700 6316 17728
rect 6415 17700 6460 17728
rect 3467 17632 4568 17660
rect 4709 17663 4767 17669
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 4709 17629 4721 17663
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 3970 17592 3976 17604
rect 2746 17564 3976 17592
rect 2593 17527 2651 17533
rect 2593 17493 2605 17527
rect 2639 17524 2651 17527
rect 2746 17524 2774 17564
rect 3970 17552 3976 17564
rect 4028 17552 4034 17604
rect 4062 17552 4068 17604
rect 4120 17592 4126 17604
rect 5092 17592 5120 17700
rect 6288 17660 6316 17700
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6638 17728 6644 17740
rect 6599 17700 6644 17728
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 7668 17737 7696 17836
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 11790 17864 11796 17876
rect 10704 17836 11796 17864
rect 8202 17796 8208 17808
rect 8163 17768 8208 17796
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 8662 17756 8668 17808
rect 8720 17796 8726 17808
rect 10594 17796 10600 17808
rect 8720 17768 10600 17796
rect 8720 17756 8726 17768
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 7653 17731 7711 17737
rect 7653 17697 7665 17731
rect 7699 17697 7711 17731
rect 9122 17728 9128 17740
rect 9083 17700 9128 17728
rect 7653 17691 7711 17697
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 9214 17688 9220 17740
rect 9272 17728 9278 17740
rect 9309 17731 9367 17737
rect 9309 17728 9321 17731
rect 9272 17700 9321 17728
rect 9272 17688 9278 17700
rect 9309 17697 9321 17700
rect 9355 17697 9367 17731
rect 9309 17691 9367 17697
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 10704 17728 10732 17836
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 11885 17867 11943 17873
rect 11885 17833 11897 17867
rect 11931 17864 11943 17867
rect 18874 17864 18880 17876
rect 11931 17836 15608 17864
rect 11931 17833 11943 17836
rect 11885 17827 11943 17833
rect 11149 17799 11207 17805
rect 11149 17765 11161 17799
rect 11195 17796 11207 17799
rect 11195 17768 14504 17796
rect 11195 17765 11207 17768
rect 11149 17759 11207 17765
rect 9456 17700 10732 17728
rect 9456 17688 9462 17700
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 12618 17728 12624 17740
rect 11296 17700 11836 17728
rect 12579 17700 12624 17728
rect 11296 17688 11302 17700
rect 7190 17660 7196 17672
rect 6288 17632 7196 17660
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 10502 17660 10508 17672
rect 10463 17632 10508 17660
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 11330 17660 11336 17672
rect 11291 17632 11336 17660
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11808 17669 11836 17700
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 13078 17728 13084 17740
rect 13039 17700 13084 17728
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 14476 17737 14504 17768
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 14461 17731 14519 17737
rect 13587 17700 14412 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12526 17660 12532 17672
rect 12483 17632 12532 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 14274 17660 14280 17672
rect 14235 17632 14280 17660
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 14384 17660 14412 17700
rect 14461 17697 14473 17731
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 14918 17688 14924 17740
rect 14976 17728 14982 17740
rect 15580 17737 15608 17836
rect 15672 17836 18880 17864
rect 15565 17731 15623 17737
rect 14976 17700 15516 17728
rect 14976 17688 14982 17700
rect 15102 17660 15108 17672
rect 14384 17632 15108 17660
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 15378 17660 15384 17672
rect 15339 17632 15384 17660
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 15488 17660 15516 17700
rect 15565 17697 15577 17731
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 15672 17660 15700 17836
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 19426 17864 19432 17876
rect 19387 17836 19432 17864
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 17126 17796 17132 17808
rect 17087 17768 17132 17796
rect 17126 17756 17132 17768
rect 17184 17756 17190 17808
rect 20073 17799 20131 17805
rect 20073 17796 20085 17799
rect 17880 17768 20085 17796
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 17678 17728 17684 17740
rect 16623 17700 17540 17728
rect 17639 17700 17684 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 15488 17632 15700 17660
rect 17512 17660 17540 17700
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 17880 17737 17908 17768
rect 20073 17765 20085 17768
rect 20119 17765 20131 17799
rect 20073 17759 20131 17765
rect 23937 17799 23995 17805
rect 23937 17765 23949 17799
rect 23983 17796 23995 17799
rect 24394 17796 24400 17808
rect 23983 17768 24400 17796
rect 23983 17765 23995 17768
rect 23937 17759 23995 17765
rect 24394 17756 24400 17768
rect 24452 17756 24458 17808
rect 17865 17731 17923 17737
rect 17865 17697 17877 17731
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 18138 17660 18144 17672
rect 17512 17632 18144 17660
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 18782 17620 18788 17672
rect 18840 17660 18846 17672
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 18840 17632 19625 17660
rect 18840 17620 18846 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 20254 17660 20260 17672
rect 20215 17632 20260 17660
rect 19613 17623 19671 17629
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20956 17632 21373 17660
rect 20956 17620 20962 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 24394 17620 24400 17672
rect 24452 17660 24458 17672
rect 24581 17663 24639 17669
rect 24581 17660 24593 17663
rect 24452 17632 24593 17660
rect 24452 17620 24458 17632
rect 24581 17629 24593 17632
rect 24627 17660 24639 17663
rect 25866 17660 25872 17672
rect 24627 17632 25872 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 4120 17564 5120 17592
rect 5261 17595 5319 17601
rect 4120 17552 4126 17564
rect 5261 17561 5273 17595
rect 5307 17561 5319 17595
rect 5261 17555 5319 17561
rect 2639 17496 2774 17524
rect 3237 17527 3295 17533
rect 2639 17493 2651 17496
rect 2593 17487 2651 17493
rect 3237 17493 3249 17527
rect 3283 17524 3295 17527
rect 4798 17524 4804 17536
rect 3283 17496 4804 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 5166 17484 5172 17536
rect 5224 17524 5230 17536
rect 5276 17524 5304 17555
rect 5350 17552 5356 17604
rect 5408 17592 5414 17604
rect 5408 17564 5453 17592
rect 5552 17564 7236 17592
rect 5408 17552 5414 17564
rect 5224 17496 5304 17524
rect 5224 17484 5230 17496
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 5552 17524 5580 17564
rect 7098 17524 7104 17536
rect 5500 17496 5580 17524
rect 7059 17496 7104 17524
rect 5500 17484 5506 17496
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 7208 17524 7236 17564
rect 7742 17552 7748 17604
rect 7800 17592 7806 17604
rect 7800 17564 7845 17592
rect 7800 17552 7806 17564
rect 8018 17552 8024 17604
rect 8076 17592 8082 17604
rect 10597 17595 10655 17601
rect 8076 17564 9996 17592
rect 8076 17552 8082 17564
rect 9398 17524 9404 17536
rect 7208 17496 9404 17524
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9968 17524 9996 17564
rect 10597 17561 10609 17595
rect 10643 17592 10655 17595
rect 16669 17595 16727 17601
rect 10643 17564 16160 17592
rect 10643 17561 10655 17564
rect 10597 17555 10655 17561
rect 13078 17524 13084 17536
rect 9968 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 13504 17496 14933 17524
rect 13504 17484 13510 17496
rect 14921 17493 14933 17496
rect 14967 17524 14979 17527
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 14967 17496 16037 17524
rect 14967 17493 14979 17496
rect 14921 17487 14979 17493
rect 16025 17493 16037 17496
rect 16071 17493 16083 17527
rect 16132 17524 16160 17564
rect 16669 17561 16681 17595
rect 16715 17561 16727 17595
rect 16669 17555 16727 17561
rect 16684 17524 16712 17555
rect 23198 17552 23204 17604
rect 23256 17592 23262 17604
rect 23385 17595 23443 17601
rect 23385 17592 23397 17595
rect 23256 17564 23397 17592
rect 23256 17552 23262 17564
rect 23385 17561 23397 17564
rect 23431 17561 23443 17595
rect 23385 17555 23443 17561
rect 23477 17595 23535 17601
rect 23477 17561 23489 17595
rect 23523 17592 23535 17595
rect 25314 17592 25320 17604
rect 23523 17564 25320 17592
rect 23523 17561 23535 17564
rect 23477 17555 23535 17561
rect 25314 17552 25320 17564
rect 25372 17552 25378 17604
rect 16132 17496 16712 17524
rect 16025 17487 16083 17493
rect 18046 17484 18052 17536
rect 18104 17524 18110 17536
rect 18325 17527 18383 17533
rect 18325 17524 18337 17527
rect 18104 17496 18337 17524
rect 18104 17484 18110 17496
rect 18325 17493 18337 17496
rect 18371 17493 18383 17527
rect 18325 17487 18383 17493
rect 21177 17527 21235 17533
rect 21177 17493 21189 17527
rect 21223 17524 21235 17527
rect 21450 17524 21456 17536
rect 21223 17496 21456 17524
rect 21223 17493 21235 17496
rect 21177 17487 21235 17493
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 23566 17484 23572 17536
rect 23624 17524 23630 17536
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 23624 17496 24685 17524
rect 23624 17484 23630 17496
rect 24673 17493 24685 17496
rect 24719 17493 24731 17527
rect 24673 17487 24731 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7156 17292 11008 17320
rect 7156 17280 7162 17292
rect 1486 17212 1492 17264
rect 1544 17252 1550 17264
rect 3145 17255 3203 17261
rect 3145 17252 3157 17255
rect 1544 17224 3157 17252
rect 1544 17212 1550 17224
rect 3145 17221 3157 17224
rect 3191 17221 3203 17255
rect 5074 17252 5080 17264
rect 4370 17224 5080 17252
rect 3145 17215 3203 17221
rect 5074 17212 5080 17224
rect 5132 17212 5138 17264
rect 6914 17252 6920 17264
rect 6012 17224 6920 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 1670 17184 1676 17196
rect 1627 17156 1676 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 6012 17193 6040 17224
rect 6914 17212 6920 17224
rect 6972 17212 6978 17264
rect 8294 17252 8300 17264
rect 8050 17224 8300 17252
rect 8294 17212 8300 17224
rect 8352 17212 8358 17264
rect 8846 17252 8852 17264
rect 8807 17224 8852 17252
rect 8846 17212 8852 17224
rect 8904 17212 8910 17264
rect 9677 17255 9735 17261
rect 9677 17221 9689 17255
rect 9723 17252 9735 17255
rect 9766 17252 9772 17264
rect 9723 17224 9772 17252
rect 9723 17221 9735 17224
rect 9677 17215 9735 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 10686 17212 10692 17264
rect 10744 17212 10750 17264
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17153 6055 17187
rect 5997 17147 6055 17153
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 8720 17156 8769 17184
rect 8720 17144 8726 17156
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9401 17187 9459 17193
rect 9180 17182 9352 17184
rect 9401 17182 9413 17187
rect 9180 17156 9413 17182
rect 9180 17144 9186 17156
rect 9324 17154 9413 17156
rect 9401 17153 9413 17154
rect 9447 17153 9459 17187
rect 10980 17184 11008 17292
rect 11054 17280 11060 17332
rect 11112 17320 11118 17332
rect 13446 17320 13452 17332
rect 11112 17292 13452 17320
rect 11112 17280 11118 17292
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 16209 17323 16267 17329
rect 13688 17292 16160 17320
rect 13688 17280 13694 17292
rect 12618 17212 12624 17264
rect 12676 17252 12682 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 12676 17224 14749 17252
rect 12676 17212 12682 17224
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 16132 17252 16160 17292
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 17034 17320 17040 17332
rect 16255 17292 17040 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 18138 17320 18144 17332
rect 18099 17292 18144 17320
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 18782 17320 18788 17332
rect 18743 17292 18788 17320
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 22830 17320 22836 17332
rect 22791 17292 22836 17320
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 38105 17323 38163 17329
rect 38105 17320 38117 17323
rect 35866 17292 38117 17320
rect 22278 17252 22284 17264
rect 16132 17224 22284 17252
rect 14737 17215 14795 17221
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 14093 17187 14151 17193
rect 10980 17182 12480 17184
rect 12544 17182 14044 17184
rect 10980 17156 14044 17182
rect 12452 17154 12572 17156
rect 9401 17147 9459 17153
rect 2869 17119 2927 17125
rect 2869 17116 2881 17119
rect 1596 17088 2881 17116
rect 1596 17060 1624 17088
rect 2869 17085 2881 17088
rect 2915 17116 2927 17119
rect 4890 17116 4896 17128
rect 2915 17088 4752 17116
rect 4851 17088 4896 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 1578 17008 1584 17060
rect 1636 17008 1642 17060
rect 4724 17048 4752 17088
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 10226 17116 10232 17128
rect 6871 17088 9352 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6564 17048 6592 17079
rect 4724 17020 6592 17048
rect 1762 16980 1768 16992
rect 1723 16952 1768 16980
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 5813 16983 5871 16989
rect 5813 16949 5825 16983
rect 5859 16980 5871 16983
rect 8110 16980 8116 16992
rect 5859 16952 8116 16980
rect 5859 16949 5871 16952
rect 5813 16943 5871 16949
rect 8110 16940 8116 16952
rect 8168 16940 8174 16992
rect 8297 16983 8355 16989
rect 8297 16949 8309 16983
rect 8343 16980 8355 16983
rect 8386 16980 8392 16992
rect 8343 16952 8392 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9324 16980 9352 17088
rect 9508 17088 10232 17116
rect 9508 17048 9536 17088
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 10468 17088 12265 17116
rect 10468 17076 10474 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17085 12495 17119
rect 14016 17116 14044 17156
rect 14093 17153 14105 17187
rect 14139 17184 14151 17187
rect 14274 17184 14280 17196
rect 14139 17156 14280 17184
rect 14139 17153 14151 17156
rect 14093 17147 14151 17153
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 16114 17184 16120 17196
rect 16075 17156 16120 17184
rect 16114 17144 16120 17156
rect 16172 17184 16178 17196
rect 16482 17184 16488 17196
rect 16172 17156 16488 17184
rect 16172 17144 16178 17156
rect 16482 17144 16488 17156
rect 16540 17184 16546 17196
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16540 17156 17049 17184
rect 16540 17144 16546 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 17037 17147 17095 17153
rect 17586 17144 17592 17196
rect 17644 17184 17650 17196
rect 18966 17184 18972 17196
rect 17644 17156 18972 17184
rect 17644 17144 17650 17156
rect 18966 17144 18972 17156
rect 19024 17184 19030 17196
rect 19610 17184 19616 17196
rect 19024 17156 19334 17184
rect 19571 17156 19616 17184
rect 19024 17144 19030 17156
rect 14182 17116 14188 17128
rect 14016 17088 14188 17116
rect 12437 17079 12495 17085
rect 12452 17048 12480 17079
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 14645 17119 14703 17125
rect 14645 17085 14657 17119
rect 14691 17116 14703 17119
rect 14826 17116 14832 17128
rect 14691 17088 14832 17116
rect 14691 17085 14703 17088
rect 14645 17079 14703 17085
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 15838 17116 15844 17128
rect 15335 17088 15844 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 16080 17088 17509 17116
rect 16080 17076 16086 17088
rect 17497 17085 17509 17088
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 17681 17119 17739 17125
rect 17681 17085 17693 17119
rect 17727 17085 17739 17119
rect 19306 17116 19334 17156
rect 19610 17144 19616 17156
rect 19668 17144 19674 17196
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20346 17184 20352 17196
rect 20119 17156 20352 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 21450 17184 21456 17196
rect 21411 17156 21456 17184
rect 21450 17144 21456 17156
rect 21508 17144 21514 17196
rect 22370 17184 22376 17196
rect 22331 17156 22376 17184
rect 22370 17144 22376 17156
rect 22428 17144 22434 17196
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17184 23535 17187
rect 23566 17184 23572 17196
rect 23523 17156 23572 17184
rect 23523 17153 23535 17156
rect 23477 17147 23535 17153
rect 23566 17144 23572 17156
rect 23624 17144 23630 17196
rect 23934 17144 23940 17196
rect 23992 17184 23998 17196
rect 24397 17187 24455 17193
rect 24397 17184 24409 17187
rect 23992 17156 24409 17184
rect 23992 17144 23998 17156
rect 24397 17153 24409 17156
rect 24443 17184 24455 17187
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 24443 17156 25881 17184
rect 24443 17153 24455 17156
rect 24397 17147 24455 17153
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17184 33747 17187
rect 35866 17184 35894 17292
rect 38105 17289 38117 17292
rect 38151 17289 38163 17323
rect 38105 17283 38163 17289
rect 38286 17184 38292 17196
rect 33735 17156 35894 17184
rect 38247 17156 38292 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 38286 17144 38292 17156
rect 38344 17144 38350 17196
rect 22186 17116 22192 17128
rect 19306 17088 22094 17116
rect 22147 17088 22192 17116
rect 17681 17079 17739 17085
rect 9416 17020 9536 17048
rect 10704 17020 12480 17048
rect 9416 16980 9444 17020
rect 9324 16952 9444 16980
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 10704 16980 10732 17020
rect 13446 17008 13452 17060
rect 13504 17048 13510 17060
rect 14918 17048 14924 17060
rect 13504 17020 14924 17048
rect 13504 17008 13510 17020
rect 14918 17008 14924 17020
rect 14976 17008 14982 17060
rect 15470 17008 15476 17060
rect 15528 17048 15534 17060
rect 17696 17048 17724 17079
rect 20254 17048 20260 17060
rect 15528 17020 17724 17048
rect 18524 17020 20260 17048
rect 15528 17008 15534 17020
rect 9548 16952 10732 16980
rect 11149 16983 11207 16989
rect 9548 16940 9554 16952
rect 11149 16949 11161 16983
rect 11195 16980 11207 16983
rect 11698 16980 11704 16992
rect 11195 16952 11704 16980
rect 11195 16949 11207 16952
rect 11149 16943 11207 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 12621 16983 12679 16989
rect 12621 16980 12633 16983
rect 11848 16952 12633 16980
rect 11848 16940 11854 16952
rect 12621 16949 12633 16952
rect 12667 16949 12679 16983
rect 12621 16943 12679 16949
rect 13909 16983 13967 16989
rect 13909 16949 13921 16983
rect 13955 16980 13967 16983
rect 16666 16980 16672 16992
rect 13955 16952 16672 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 16853 16983 16911 16989
rect 16853 16949 16865 16983
rect 16899 16980 16911 16983
rect 18524 16980 18552 17020
rect 20254 17008 20260 17020
rect 20312 17008 20318 17060
rect 22066 17048 22094 17088
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 23293 17119 23351 17125
rect 23293 17085 23305 17119
rect 23339 17085 23351 17119
rect 23293 17079 23351 17085
rect 22554 17048 22560 17060
rect 22066 17020 22560 17048
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 23308 17048 23336 17079
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 25041 17119 25099 17125
rect 25041 17116 25053 17119
rect 24636 17088 25053 17116
rect 24636 17076 24642 17088
rect 25041 17085 25053 17088
rect 25087 17085 25099 17119
rect 25041 17079 25099 17085
rect 33781 17051 33839 17057
rect 33781 17048 33793 17051
rect 23308 17020 33793 17048
rect 33781 17017 33793 17020
rect 33827 17017 33839 17051
rect 33781 17011 33839 17017
rect 16899 16952 18552 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 19392 16952 19441 16980
rect 19392 16940 19398 16952
rect 19429 16949 19441 16952
rect 19475 16949 19487 16983
rect 19429 16943 19487 16949
rect 20165 16983 20223 16989
rect 20165 16949 20177 16983
rect 20211 16980 20223 16983
rect 20714 16980 20720 16992
rect 20211 16952 20720 16980
rect 20211 16949 20223 16952
rect 20165 16943 20223 16949
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21358 16980 21364 16992
rect 21315 16952 21364 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 23198 16940 23204 16992
rect 23256 16980 23262 16992
rect 23661 16983 23719 16989
rect 23661 16980 23673 16983
rect 23256 16952 23673 16980
rect 23256 16940 23262 16952
rect 23661 16949 23673 16952
rect 23707 16949 23719 16983
rect 24486 16980 24492 16992
rect 24447 16952 24492 16980
rect 23661 16943 23719 16949
rect 24486 16940 24492 16952
rect 24544 16940 24550 16992
rect 25682 16980 25688 16992
rect 25643 16952 25688 16980
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 11054 16776 11060 16788
rect 4948 16748 11060 16776
rect 4948 16736 4954 16748
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 15194 16736 15200 16788
rect 15252 16776 15258 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 15252 16748 16681 16776
rect 15252 16736 15258 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18196 16748 18337 16776
rect 18196 16736 18202 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 19610 16736 19616 16788
rect 19668 16776 19674 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 19668 16748 20085 16776
rect 19668 16736 19674 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 21542 16776 21548 16788
rect 21503 16748 21548 16776
rect 20073 16739 20131 16745
rect 21542 16736 21548 16748
rect 21600 16736 21606 16788
rect 23198 16776 23204 16788
rect 23159 16748 23204 16776
rect 23198 16736 23204 16748
rect 23256 16736 23262 16788
rect 5810 16668 5816 16720
rect 5868 16708 5874 16720
rect 6730 16708 6736 16720
rect 5868 16680 6736 16708
rect 5868 16668 5874 16680
rect 6730 16668 6736 16680
rect 6788 16668 6794 16720
rect 8386 16708 8392 16720
rect 6840 16680 8392 16708
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16640 2010 16652
rect 2590 16640 2596 16652
rect 2004 16612 2596 16640
rect 2004 16600 2010 16612
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 6840 16640 6868 16680
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 17402 16708 17408 16720
rect 10428 16680 17408 16708
rect 4295 16612 6868 16640
rect 6917 16643 6975 16649
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 7374 16640 7380 16652
rect 6963 16612 7380 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16640 7619 16643
rect 8018 16640 8024 16652
rect 7607 16612 8024 16640
rect 7607 16609 7619 16612
rect 7561 16603 7619 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8404 16640 8432 16668
rect 10428 16640 10456 16680
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 33410 16708 33416 16720
rect 17972 16680 33416 16708
rect 8404 16612 10456 16640
rect 10594 16600 10600 16652
rect 10652 16640 10658 16652
rect 10873 16643 10931 16649
rect 10873 16640 10885 16643
rect 10652 16612 10885 16640
rect 10652 16600 10658 16612
rect 10873 16609 10885 16612
rect 10919 16609 10931 16643
rect 10873 16603 10931 16609
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 13722 16640 13728 16652
rect 12115 16612 13728 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 17972 16649 18000 16680
rect 33410 16668 33416 16680
rect 33468 16668 33474 16720
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 13872 16612 16497 16640
rect 13872 16600 13878 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16609 18015 16643
rect 18138 16640 18144 16652
rect 18099 16612 18144 16640
rect 17957 16603 18015 16609
rect 18138 16600 18144 16612
rect 18196 16600 18202 16652
rect 21174 16640 21180 16652
rect 21135 16612 21180 16640
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 22554 16640 22560 16652
rect 22515 16612 22560 16640
rect 22554 16600 22560 16612
rect 22612 16600 22618 16652
rect 24578 16640 24584 16652
rect 24539 16612 24584 16640
rect 24578 16600 24584 16612
rect 24636 16600 24642 16652
rect 1578 16532 1584 16584
rect 1636 16572 1642 16584
rect 1673 16575 1731 16581
rect 1673 16572 1685 16575
rect 1636 16544 1685 16572
rect 1636 16532 1642 16544
rect 1673 16541 1685 16544
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 9122 16572 9128 16584
rect 9083 16544 9128 16572
rect 3973 16535 4031 16541
rect 2958 16464 2964 16516
rect 3016 16464 3022 16516
rect 3988 16504 4016 16535
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 4154 16504 4160 16516
rect 3988 16476 4160 16504
rect 4154 16464 4160 16476
rect 4212 16464 4218 16516
rect 4890 16464 4896 16516
rect 4948 16464 4954 16516
rect 6270 16504 6276 16516
rect 6231 16476 6276 16504
rect 6270 16464 6276 16476
rect 6328 16464 6334 16516
rect 6365 16507 6423 16513
rect 6365 16473 6377 16507
rect 6411 16473 6423 16507
rect 6365 16467 6423 16473
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 5534 16436 5540 16448
rect 3467 16408 5540 16436
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 5718 16436 5724 16448
rect 5679 16408 5724 16436
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 6086 16396 6092 16448
rect 6144 16436 6150 16448
rect 6380 16436 6408 16467
rect 7650 16464 7656 16516
rect 7708 16504 7714 16516
rect 8205 16507 8263 16513
rect 7708 16476 7753 16504
rect 7708 16464 7714 16476
rect 8205 16473 8217 16507
rect 8251 16473 8263 16507
rect 9398 16504 9404 16516
rect 9359 16476 9404 16504
rect 8205 16467 8263 16473
rect 6144 16408 6408 16436
rect 6144 16396 6150 16408
rect 7190 16396 7196 16448
rect 7248 16436 7254 16448
rect 8018 16436 8024 16448
rect 7248 16408 8024 16436
rect 7248 16396 7254 16408
rect 8018 16396 8024 16408
rect 8076 16436 8082 16448
rect 8220 16436 8248 16467
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 9490 16464 9496 16516
rect 9548 16504 9554 16516
rect 11624 16504 11652 16535
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 12216 16544 12265 16572
rect 12216 16532 12222 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 14274 16532 14280 16584
rect 14332 16572 14338 16584
rect 14461 16575 14519 16581
rect 14461 16572 14473 16575
rect 14332 16544 14473 16572
rect 14332 16532 14338 16544
rect 14461 16541 14473 16544
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 16390 16572 16396 16584
rect 16347 16544 16396 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16572 19671 16575
rect 20162 16572 20168 16584
rect 19659 16544 20168 16572
rect 19659 16541 19671 16544
rect 19613 16535 19671 16541
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16572 20315 16575
rect 20346 16572 20352 16584
rect 20303 16544 20352 16572
rect 20303 16541 20315 16544
rect 20257 16535 20315 16541
rect 20346 16532 20352 16544
rect 20404 16532 20410 16584
rect 22738 16572 22744 16584
rect 22699 16544 22744 16572
rect 22738 16532 22744 16544
rect 22796 16532 22802 16584
rect 23566 16532 23572 16584
rect 23624 16572 23630 16584
rect 23845 16575 23903 16581
rect 23845 16572 23857 16575
rect 23624 16544 23857 16572
rect 23624 16532 23630 16544
rect 23845 16541 23857 16544
rect 23891 16572 23903 16575
rect 24394 16572 24400 16584
rect 23891 16544 24400 16572
rect 23891 16541 23903 16544
rect 23845 16535 23903 16541
rect 24394 16532 24400 16544
rect 24452 16532 24458 16584
rect 24762 16572 24768 16584
rect 24723 16544 24768 16572
rect 24762 16532 24768 16544
rect 24820 16532 24826 16584
rect 14642 16504 14648 16516
rect 9548 16476 9890 16504
rect 11624 16476 14648 16504
rect 9548 16464 9554 16476
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 15194 16504 15200 16516
rect 15155 16476 15200 16504
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15289 16507 15347 16513
rect 15289 16473 15301 16507
rect 15335 16504 15347 16507
rect 15378 16504 15384 16516
rect 15335 16476 15384 16504
rect 15335 16473 15347 16476
rect 15289 16467 15347 16473
rect 15378 16464 15384 16476
rect 15436 16464 15442 16516
rect 15838 16504 15844 16516
rect 15799 16476 15844 16504
rect 15838 16464 15844 16476
rect 15896 16464 15902 16516
rect 8076 16408 8248 16436
rect 8076 16396 8082 16408
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 11146 16436 11152 16448
rect 8444 16408 11152 16436
rect 8444 16396 8450 16408
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 11425 16439 11483 16445
rect 11425 16405 11437 16439
rect 11471 16436 11483 16439
rect 12618 16436 12624 16448
rect 11471 16408 12624 16436
rect 11471 16405 11483 16408
rect 11425 16399 11483 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 13541 16439 13599 16445
rect 12768 16408 12813 16436
rect 12768 16396 12774 16408
rect 13541 16405 13553 16439
rect 13587 16436 13599 16439
rect 14458 16436 14464 16448
rect 13587 16408 14464 16436
rect 13587 16405 13599 16408
rect 13541 16399 13599 16405
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16436 14611 16439
rect 15470 16436 15476 16448
rect 14599 16408 15476 16436
rect 14599 16405 14611 16408
rect 14553 16399 14611 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 19426 16436 19432 16448
rect 19387 16408 19432 16436
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 23658 16436 23664 16448
rect 23619 16408 23664 16436
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 25225 16439 25283 16445
rect 25225 16436 25237 16439
rect 24084 16408 25237 16436
rect 24084 16396 24090 16408
rect 25225 16405 25237 16408
rect 25271 16436 25283 16439
rect 29730 16436 29736 16448
rect 25271 16408 29736 16436
rect 25271 16405 25283 16408
rect 25225 16399 25283 16405
rect 29730 16396 29736 16408
rect 29788 16396 29794 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2096 16204 3648 16232
rect 2096 16192 2102 16204
rect 3620 16176 3648 16204
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 7650 16232 7656 16244
rect 5040 16204 7656 16232
rect 5040 16192 5046 16204
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 11149 16235 11207 16241
rect 7852 16204 11008 16232
rect 3326 16164 3332 16176
rect 3082 16136 3332 16164
rect 3326 16124 3332 16136
rect 3384 16124 3390 16176
rect 3602 16164 3608 16176
rect 3563 16136 3608 16164
rect 3602 16124 3608 16136
rect 3660 16124 3666 16176
rect 5350 16124 5356 16176
rect 5408 16124 5414 16176
rect 5718 16124 5724 16176
rect 5776 16164 5782 16176
rect 7190 16164 7196 16176
rect 5776 16136 7196 16164
rect 5776 16124 5782 16136
rect 7190 16124 7196 16136
rect 7248 16124 7254 16176
rect 7469 16167 7527 16173
rect 7469 16133 7481 16167
rect 7515 16164 7527 16167
rect 7852 16164 7880 16204
rect 7515 16136 7880 16164
rect 7515 16133 7527 16136
rect 7469 16127 7527 16133
rect 10134 16124 10140 16176
rect 10192 16124 10198 16176
rect 10980 16164 11008 16204
rect 11149 16201 11161 16235
rect 11195 16232 11207 16235
rect 11514 16232 11520 16244
rect 11195 16204 11520 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 13265 16235 13323 16241
rect 13265 16201 13277 16235
rect 13311 16232 13323 16235
rect 13814 16232 13820 16244
rect 13311 16204 13820 16232
rect 13311 16201 13323 16204
rect 13265 16195 13323 16201
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 16114 16232 16120 16244
rect 13924 16204 16120 16232
rect 12250 16164 12256 16176
rect 10980 16136 12256 16164
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 13354 16164 13360 16176
rect 12406 16136 13360 16164
rect 1578 16028 1584 16040
rect 1539 16000 1584 16028
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 3234 16028 3240 16040
rect 1903 16000 3240 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 4062 16028 4068 16040
rect 4023 16000 4068 16028
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4341 16031 4399 16037
rect 4341 15997 4353 16031
rect 4387 16028 4399 16031
rect 5736 16028 5764 16124
rect 6546 16096 6552 16108
rect 6507 16068 6552 16096
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 8570 16056 8576 16108
rect 8628 16056 8634 16108
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9180 16068 9413 16096
rect 9180 16056 9186 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 12406 16096 12434 16136
rect 13354 16124 13360 16136
rect 13412 16164 13418 16176
rect 13924 16164 13952 16204
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 18892 16204 20116 16232
rect 14090 16164 14096 16176
rect 13412 16136 13952 16164
rect 14051 16136 14096 16164
rect 13412 16124 13418 16136
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 14458 16124 14464 16176
rect 14516 16164 14522 16176
rect 18322 16164 18328 16176
rect 14516 16136 16896 16164
rect 18283 16136 18328 16164
rect 14516 16124 14522 16136
rect 11204 16068 12434 16096
rect 13449 16099 13507 16105
rect 11204 16056 11210 16068
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 13814 16096 13820 16108
rect 13495 16068 13820 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 16868 16105 16896 16136
rect 18322 16124 18328 16136
rect 18380 16124 18386 16176
rect 18892 16173 18920 16204
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16133 18935 16167
rect 18877 16127 18935 16133
rect 19426 16124 19432 16176
rect 19484 16164 19490 16176
rect 20088 16173 20116 16204
rect 20162 16192 20168 16244
rect 20220 16232 20226 16244
rect 22005 16235 22063 16241
rect 22005 16232 22017 16235
rect 20220 16204 22017 16232
rect 20220 16192 20226 16204
rect 22005 16201 22017 16204
rect 22051 16201 22063 16235
rect 22738 16232 22744 16244
rect 22699 16204 22744 16232
rect 22005 16195 22063 16201
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 24026 16232 24032 16244
rect 23987 16204 24032 16232
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 24489 16235 24547 16241
rect 24489 16201 24501 16235
rect 24535 16232 24547 16235
rect 24762 16232 24768 16244
rect 24535 16204 24768 16232
rect 24535 16201 24547 16204
rect 24489 16195 24547 16201
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 19521 16167 19579 16173
rect 19521 16164 19533 16167
rect 19484 16136 19533 16164
rect 19484 16124 19490 16136
rect 19521 16133 19533 16136
rect 19567 16133 19579 16167
rect 19521 16127 19579 16133
rect 20073 16167 20131 16173
rect 20073 16133 20085 16167
rect 20119 16164 20131 16167
rect 21634 16164 21640 16176
rect 20119 16136 21640 16164
rect 20119 16133 20131 16136
rect 20073 16127 20131 16133
rect 21634 16124 21640 16136
rect 21692 16124 21698 16176
rect 24854 16164 24860 16176
rect 22066 16136 24860 16164
rect 16853 16099 16911 16105
rect 15028 16068 16804 16096
rect 4387 16000 5764 16028
rect 5813 16031 5871 16037
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 6178 16028 6184 16040
rect 5859 16000 6184 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 7182 16031 7240 16037
rect 7182 15997 7194 16031
rect 7228 16028 7240 16031
rect 9140 16028 9168 16056
rect 7228 16000 9168 16028
rect 9677 16031 9735 16037
rect 7228 15997 7240 16000
rect 7182 15991 7240 15997
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 10042 16028 10048 16040
rect 9723 16000 10048 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11514 16028 11520 16040
rect 11020 16000 11520 16028
rect 11020 15988 11026 16000
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 11698 16028 11704 16040
rect 11659 16000 11704 16028
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 11882 16028 11888 16040
rect 11843 16000 11888 16028
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 13998 16028 14004 16040
rect 13959 16000 14004 16028
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 15028 16028 15056 16068
rect 14476 16000 15056 16028
rect 14476 15960 14504 16000
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15289 16031 15347 16037
rect 15160 16000 15205 16028
rect 15160 15988 15166 16000
rect 15289 15997 15301 16031
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 10704 15932 14504 15960
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6641 15895 6699 15901
rect 6641 15892 6653 15895
rect 6052 15864 6653 15892
rect 6052 15852 6058 15864
rect 6641 15861 6653 15864
rect 6687 15861 6699 15895
rect 6641 15855 6699 15861
rect 8941 15895 8999 15901
rect 8941 15861 8953 15895
rect 8987 15892 8999 15895
rect 9398 15892 9404 15904
rect 8987 15864 9404 15892
rect 8987 15861 8999 15864
rect 8941 15855 8999 15861
rect 9398 15852 9404 15864
rect 9456 15892 9462 15904
rect 10704 15892 10732 15932
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 14608 15932 14653 15960
rect 14608 15920 14614 15932
rect 9456 15864 10732 15892
rect 9456 15852 9462 15864
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 10928 15864 12081 15892
rect 10928 15852 10934 15864
rect 12069 15861 12081 15864
rect 12115 15861 12127 15895
rect 12069 15855 12127 15861
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 15304 15892 15332 15991
rect 16776 15960 16804 16068
rect 16853 16065 16865 16099
rect 16899 16065 16911 16099
rect 20714 16096 20720 16108
rect 20675 16068 20720 16096
rect 16853 16059 16911 16065
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 17034 16028 17040 16040
rect 16995 16000 17040 16028
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 18230 16028 18236 16040
rect 18191 16000 18236 16028
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 19426 16028 19432 16040
rect 19387 16000 19432 16028
rect 19426 15988 19432 16000
rect 19484 15988 19490 16040
rect 20070 15988 20076 16040
rect 20128 16028 20134 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20128 16000 20545 16028
rect 20128 15988 20134 16000
rect 20533 15997 20545 16000
rect 20579 16028 20591 16031
rect 22066 16028 22094 16136
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16096 22983 16099
rect 23658 16096 23664 16108
rect 22971 16068 23664 16096
rect 22971 16065 22983 16068
rect 22925 16059 22983 16065
rect 20579 16000 22094 16028
rect 20579 15997 20591 16000
rect 20533 15991 20591 15997
rect 18506 15960 18512 15972
rect 16776 15932 18512 15960
rect 18506 15920 18512 15932
rect 18564 15920 18570 15972
rect 22204 15960 22232 16059
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 24673 16099 24731 16105
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 25682 16096 25688 16108
rect 24719 16068 25688 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 29730 16096 29736 16108
rect 29691 16068 29736 16096
rect 29730 16056 29736 16068
rect 29788 16056 29794 16108
rect 36078 16056 36084 16108
rect 36136 16096 36142 16108
rect 38013 16099 38071 16105
rect 38013 16096 38025 16099
rect 36136 16068 38025 16096
rect 36136 16056 36142 16068
rect 38013 16065 38025 16068
rect 38059 16065 38071 16099
rect 38013 16059 38071 16065
rect 23106 15988 23112 16040
rect 23164 16028 23170 16040
rect 23385 16031 23443 16037
rect 23385 16028 23397 16031
rect 23164 16000 23397 16028
rect 23164 15988 23170 16000
rect 23385 15997 23397 16000
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 23569 16031 23627 16037
rect 23569 15997 23581 16031
rect 23615 16028 23627 16031
rect 24486 16028 24492 16040
rect 23615 16000 24492 16028
rect 23615 15997 23627 16000
rect 23569 15991 23627 15997
rect 24486 15988 24492 16000
rect 24544 15988 24550 16040
rect 20088 15932 22232 15960
rect 15470 15892 15476 15904
rect 13688 15864 15332 15892
rect 15431 15864 15476 15892
rect 13688 15852 13694 15864
rect 15470 15852 15476 15864
rect 15528 15892 15534 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 15528 15864 17233 15892
rect 15528 15852 15534 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 18524 15892 18552 15920
rect 20088 15892 20116 15932
rect 18524 15864 20116 15892
rect 17221 15855 17279 15861
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20312 15864 20913 15892
rect 20312 15852 20318 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 29825 15895 29883 15901
rect 29825 15861 29837 15895
rect 29871 15892 29883 15895
rect 31662 15892 31668 15904
rect 29871 15864 31668 15892
rect 29871 15861 29883 15864
rect 29825 15855 29883 15861
rect 31662 15852 31668 15864
rect 31720 15852 31726 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 3421 15691 3479 15697
rect 3421 15657 3433 15691
rect 3467 15688 3479 15691
rect 6270 15688 6276 15700
rect 3467 15660 6276 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 11146 15688 11152 15700
rect 6604 15660 11152 15688
rect 6604 15648 6610 15660
rect 11146 15648 11152 15660
rect 11204 15688 11210 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11204 15660 11345 15688
rect 11204 15648 11210 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 13633 15691 13691 15697
rect 13633 15657 13645 15691
rect 13679 15688 13691 15691
rect 13906 15688 13912 15700
rect 13679 15660 13912 15688
rect 13679 15657 13691 15660
rect 13633 15651 13691 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14553 15691 14611 15697
rect 14553 15657 14565 15691
rect 14599 15688 14611 15691
rect 17034 15688 17040 15700
rect 14599 15660 17040 15688
rect 14599 15657 14611 15660
rect 14553 15651 14611 15657
rect 17034 15648 17040 15660
rect 17092 15648 17098 15700
rect 20254 15688 20260 15700
rect 20215 15660 20260 15688
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 6641 15623 6699 15629
rect 6641 15589 6653 15623
rect 6687 15620 6699 15623
rect 7926 15620 7932 15632
rect 6687 15592 7932 15620
rect 6687 15589 6699 15592
rect 6641 15583 6699 15589
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 8938 15580 8944 15632
rect 8996 15620 9002 15632
rect 9953 15623 10011 15629
rect 9953 15620 9965 15623
rect 8996 15592 9965 15620
rect 8996 15580 9002 15592
rect 9953 15589 9965 15592
rect 9999 15620 10011 15623
rect 10870 15620 10876 15632
rect 9999 15592 10876 15620
rect 9999 15589 10011 15592
rect 9953 15583 10011 15589
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 15470 15620 15476 15632
rect 10980 15592 15476 15620
rect 2130 15552 2136 15564
rect 2091 15524 2136 15552
rect 2130 15512 2136 15524
rect 2188 15512 2194 15564
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 2866 15552 2872 15564
rect 2823 15524 2872 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 2961 15555 3019 15561
rect 2961 15521 2973 15555
rect 3007 15552 3019 15555
rect 3050 15552 3056 15564
rect 3007 15524 3056 15552
rect 3007 15521 3019 15524
rect 2961 15515 3019 15521
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15552 5227 15555
rect 6730 15552 6736 15564
rect 5215 15524 6736 15552
rect 5215 15521 5227 15524
rect 5169 15515 5227 15521
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 7699 15524 8340 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 1854 15484 1860 15496
rect 1815 15456 1860 15484
rect 1854 15444 1860 15456
rect 1912 15484 1918 15496
rect 3973 15487 4031 15493
rect 1912 15456 2774 15484
rect 1912 15444 1918 15456
rect 2746 15416 2774 15456
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 8312 15484 8340 15524
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 10980 15561 11008 15592
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 16850 15620 16856 15632
rect 16811 15592 16856 15620
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 18046 15620 18052 15632
rect 17696 15592 18052 15620
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 8444 15524 9781 15552
rect 8444 15512 8450 15524
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 10965 15555 11023 15561
rect 10965 15521 10977 15555
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 12802 15552 12808 15564
rect 12115 15524 12808 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 17696 15561 17724 15592
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 17681 15555 17739 15561
rect 14608 15524 15976 15552
rect 14608 15512 14614 15524
rect 9582 15484 9588 15496
rect 8312 15456 8708 15484
rect 9543 15456 9588 15484
rect 4893 15447 4951 15453
rect 3988 15416 4016 15447
rect 2746 15388 4016 15416
rect 4249 15419 4307 15425
rect 4249 15385 4261 15419
rect 4295 15416 4307 15419
rect 4614 15416 4620 15428
rect 4295 15388 4620 15416
rect 4295 15385 4307 15388
rect 4249 15379 4307 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 4908 15416 4936 15447
rect 5442 15416 5448 15428
rect 4908 15388 5448 15416
rect 5442 15376 5448 15388
rect 5500 15376 5506 15428
rect 6454 15416 6460 15428
rect 6394 15388 6460 15416
rect 6454 15376 6460 15388
rect 6512 15376 6518 15428
rect 7742 15376 7748 15428
rect 7800 15416 7806 15428
rect 7800 15388 7845 15416
rect 7800 15376 7806 15388
rect 8018 15376 8024 15428
rect 8076 15416 8082 15428
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 8076 15388 8309 15416
rect 8076 15376 8082 15388
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8680 15416 8708 15456
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15484 11207 15487
rect 11974 15484 11980 15496
rect 11195 15456 11980 15484
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12250 15484 12256 15496
rect 12211 15456 12256 15484
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 13538 15484 13544 15496
rect 12820 15456 13544 15484
rect 12820 15428 12848 15456
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 14826 15484 14832 15496
rect 14783 15456 14832 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 11790 15416 11796 15428
rect 8680 15388 11796 15416
rect 8297 15379 8355 15385
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 12802 15376 12808 15428
rect 12860 15376 12866 15428
rect 15286 15416 15292 15428
rect 15247 15388 15292 15416
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 15381 15419 15439 15425
rect 15381 15385 15393 15419
rect 15427 15416 15439 15419
rect 15746 15416 15752 15428
rect 15427 15388 15752 15416
rect 15427 15385 15439 15388
rect 15381 15379 15439 15385
rect 15746 15376 15752 15388
rect 15804 15376 15810 15428
rect 15948 15425 15976 15524
rect 17681 15521 17693 15555
rect 17727 15521 17739 15555
rect 17681 15515 17739 15521
rect 17862 15512 17868 15564
rect 17920 15552 17926 15564
rect 17957 15555 18015 15561
rect 17957 15552 17969 15555
rect 17920 15524 17969 15552
rect 17920 15512 17926 15524
rect 17957 15521 17969 15524
rect 18003 15521 18015 15555
rect 17957 15515 18015 15521
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19797 15555 19855 15561
rect 19797 15552 19809 15555
rect 19392 15524 19809 15552
rect 19392 15512 19398 15524
rect 19797 15521 19809 15524
rect 19843 15521 19855 15555
rect 19797 15515 19855 15521
rect 20162 15512 20168 15564
rect 20220 15552 20226 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20220 15524 20913 15552
rect 20220 15512 20226 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 22278 15552 22284 15564
rect 22239 15524 22284 15552
rect 20901 15515 20959 15521
rect 22278 15512 22284 15524
rect 22336 15552 22342 15564
rect 25682 15552 25688 15564
rect 22336 15524 25688 15552
rect 22336 15512 22342 15524
rect 25682 15512 25688 15524
rect 25740 15512 25746 15564
rect 16482 15484 16488 15496
rect 16443 15456 16488 15484
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 16669 15487 16727 15493
rect 16669 15453 16681 15487
rect 16715 15484 16727 15487
rect 16942 15484 16948 15496
rect 16715 15456 16948 15484
rect 16715 15453 16727 15456
rect 16669 15447 16727 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 20438 15484 20444 15496
rect 19659 15456 20444 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20806 15484 20812 15496
rect 20763 15456 20812 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 22465 15487 22523 15493
rect 22465 15453 22477 15487
rect 22511 15484 22523 15487
rect 24118 15484 24124 15496
rect 22511 15456 24124 15484
rect 22511 15453 22523 15456
rect 22465 15447 22523 15453
rect 24118 15444 24124 15456
rect 24176 15444 24182 15496
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 25130 15484 25136 15496
rect 24627 15456 25136 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 25130 15444 25136 15456
rect 25188 15444 25194 15496
rect 15933 15419 15991 15425
rect 15933 15385 15945 15419
rect 15979 15416 15991 15419
rect 17218 15416 17224 15428
rect 15979 15388 17224 15416
rect 15979 15385 15991 15388
rect 15933 15379 15991 15385
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 17770 15376 17776 15428
rect 17828 15416 17834 15428
rect 17828 15388 17873 15416
rect 17828 15376 17834 15388
rect 19978 15376 19984 15428
rect 20036 15416 20042 15428
rect 22738 15416 22744 15428
rect 20036 15388 22744 15416
rect 20036 15376 20042 15388
rect 22738 15376 22744 15388
rect 22796 15376 22802 15428
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 9582 15348 9588 15360
rect 3844 15320 9588 15348
rect 3844 15308 3850 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 12710 15348 12716 15360
rect 12671 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 21358 15348 21364 15360
rect 21319 15320 21364 15348
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 22922 15348 22928 15360
rect 22883 15320 22928 15348
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 23382 15348 23388 15360
rect 23343 15320 23388 15348
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 24670 15348 24676 15360
rect 24631 15320 24676 15348
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 5442 15144 5448 15156
rect 4264 15116 5448 15144
rect 2498 15036 2504 15088
rect 2556 15036 2562 15088
rect 3510 15036 3516 15088
rect 3568 15076 3574 15088
rect 3786 15076 3792 15088
rect 3568 15048 3792 15076
rect 3568 15036 3574 15048
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4264 15017 4292 15116
rect 5442 15104 5448 15116
rect 5500 15144 5506 15156
rect 6546 15144 6552 15156
rect 5500 15116 6552 15144
rect 5500 15104 5506 15116
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 9490 15144 9496 15156
rect 6788 15116 9496 15144
rect 6788 15104 6794 15116
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 9824 15116 10609 15144
rect 9824 15104 9830 15116
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 10597 15107 10655 15113
rect 10704 15116 13124 15144
rect 4982 15036 4988 15088
rect 5040 15036 5046 15088
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 6825 15079 6883 15085
rect 6825 15076 6837 15079
rect 6328 15048 6837 15076
rect 6328 15036 6334 15048
rect 6825 15045 6837 15048
rect 6871 15076 6883 15079
rect 7098 15076 7104 15088
rect 6871 15048 7104 15076
rect 6871 15045 6883 15048
rect 6825 15039 6883 15045
rect 7098 15036 7104 15048
rect 7156 15036 7162 15088
rect 7834 15036 7840 15088
rect 7892 15036 7898 15088
rect 9122 15076 9128 15088
rect 8864 15048 9128 15076
rect 8864 15017 8892 15048
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 4249 15011 4307 15017
rect 4249 15008 4261 15011
rect 4120 14980 4261 15008
rect 4120 14968 4126 14980
rect 4249 14977 4261 14980
rect 4295 14977 4307 15011
rect 4249 14971 4307 14977
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 10226 14968 10232 15020
rect 10284 14968 10290 15020
rect 10704 15008 10732 15116
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 13096 15076 13124 15116
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 14461 15147 14519 15153
rect 14461 15144 14473 15147
rect 13872 15116 14473 15144
rect 13872 15104 13878 15116
rect 14461 15113 14473 15116
rect 14507 15113 14519 15147
rect 14461 15107 14519 15113
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16850 15144 16856 15156
rect 15795 15116 16856 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 16960 15116 17540 15144
rect 16960 15076 16988 15116
rect 17402 15076 17408 15088
rect 12400 15048 13032 15076
rect 13096 15048 16988 15076
rect 17363 15048 17408 15076
rect 12400 15036 12406 15048
rect 13004 15017 13032 15048
rect 17402 15036 17408 15048
rect 17460 15036 17466 15088
rect 17512 15076 17540 15116
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 18380 15116 18613 15144
rect 18380 15104 18386 15116
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 22922 15144 22928 15156
rect 18601 15107 18659 15113
rect 18708 15116 22094 15144
rect 22883 15116 22928 15144
rect 18708 15076 18736 15116
rect 19242 15076 19248 15088
rect 17512 15048 18736 15076
rect 19203 15048 19248 15076
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 19337 15079 19395 15085
rect 19337 15045 19349 15079
rect 19383 15076 19395 15079
rect 19978 15076 19984 15088
rect 19383 15048 19984 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 22066 15076 22094 15116
rect 22922 15104 22928 15116
rect 22980 15104 22986 15156
rect 23198 15104 23204 15156
rect 23256 15144 23262 15156
rect 34701 15147 34759 15153
rect 23256 15116 24072 15144
rect 23256 15104 23262 15116
rect 23934 15076 23940 15088
rect 22066 15048 23940 15076
rect 23934 15036 23940 15048
rect 23992 15036 23998 15088
rect 10612 14980 10732 15008
rect 12989 15011 13047 15017
rect 1670 14900 1676 14952
rect 1728 14940 1734 14952
rect 1765 14943 1823 14949
rect 1765 14940 1777 14943
rect 1728 14912 1777 14940
rect 1728 14900 1734 14912
rect 1765 14909 1777 14912
rect 1811 14909 1823 14943
rect 1765 14903 1823 14909
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 3418 14940 3424 14952
rect 2087 14912 3424 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 5810 14940 5816 14952
rect 4571 14912 5816 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 6546 14940 6552 14952
rect 6507 14912 6552 14940
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 9122 14940 9128 14952
rect 7248 14912 8432 14940
rect 9035 14912 9128 14940
rect 7248 14900 7254 14912
rect 6178 14872 6184 14884
rect 5552 14844 6184 14872
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 5552 14804 5580 14844
rect 6178 14832 6184 14844
rect 6236 14832 6242 14884
rect 2740 14776 5580 14804
rect 2740 14764 2746 14776
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5684 14776 6009 14804
rect 5684 14764 5690 14776
rect 5997 14773 6009 14776
rect 6043 14773 6055 14807
rect 5997 14767 6055 14773
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 8168 14776 8309 14804
rect 8168 14764 8174 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8404 14804 8432 14912
rect 9122 14900 9128 14912
rect 9180 14940 9186 14952
rect 10612 14940 10640 14980
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 13596 14980 14657 15008
rect 13596 14968 13602 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 14645 14971 14703 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 15008 19947 15011
rect 22186 15008 22192 15020
rect 19935 14980 22192 15008
rect 19935 14977 19947 14980
rect 19889 14971 19947 14977
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 23382 15008 23388 15020
rect 22327 14980 23388 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 24044 15017 24072 15116
rect 34701 15113 34713 15147
rect 34747 15144 34759 15147
rect 36078 15144 36084 15156
rect 34747 15116 36084 15144
rect 34747 15113 34759 15116
rect 34701 15107 34759 15113
rect 36078 15104 36084 15116
rect 36136 15104 36142 15156
rect 31662 15036 31668 15088
rect 31720 15076 31726 15088
rect 31720 15048 35572 15076
rect 31720 15036 31726 15048
rect 23569 15011 23627 15017
rect 23569 14977 23581 15011
rect 23615 14977 23627 15011
rect 23569 14971 23627 14977
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 15008 24087 15011
rect 24857 15011 24915 15017
rect 24857 15008 24869 15011
rect 24075 14980 24869 15008
rect 24075 14977 24087 14980
rect 24029 14971 24087 14977
rect 24857 14977 24869 14980
rect 24903 14977 24915 15011
rect 24857 14971 24915 14977
rect 33505 15011 33563 15017
rect 33505 14977 33517 15011
rect 33551 14977 33563 15011
rect 33505 14971 33563 14977
rect 9180 14912 10640 14940
rect 9180 14900 9186 14912
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11701 14943 11759 14949
rect 11701 14940 11713 14943
rect 10744 14912 11713 14940
rect 10744 14900 10750 14912
rect 11701 14909 11713 14912
rect 11747 14909 11759 14943
rect 11701 14903 11759 14909
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14940 11943 14943
rect 12526 14940 12532 14952
rect 11931 14928 12204 14940
rect 12360 14928 12532 14940
rect 11931 14912 12532 14928
rect 11931 14909 11943 14912
rect 11885 14903 11943 14909
rect 12176 14900 12388 14912
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 12820 14872 12848 14903
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 15102 14940 15108 14952
rect 13320 14912 15108 14940
rect 13320 14900 13326 14912
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 15286 14940 15292 14952
rect 15247 14912 15292 14940
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 17310 14940 17316 14952
rect 15396 14912 17316 14940
rect 12176 14844 12848 14872
rect 11238 14804 11244 14816
rect 8404 14776 11244 14804
rect 8297 14767 8355 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 11388 14776 12081 14804
rect 11388 14764 11394 14776
rect 12069 14773 12081 14776
rect 12115 14804 12127 14807
rect 12176 14804 12204 14844
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 15396 14872 15424 14912
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 20070 14900 20076 14952
rect 20128 14940 20134 14952
rect 20533 14943 20591 14949
rect 20533 14940 20545 14943
rect 20128 14912 20545 14940
rect 20128 14900 20134 14912
rect 20533 14909 20545 14912
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 20717 14943 20775 14949
rect 20717 14909 20729 14943
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 22465 14943 22523 14949
rect 22465 14909 22477 14943
rect 22511 14940 22523 14943
rect 23584 14940 23612 14971
rect 25314 14940 25320 14952
rect 22511 14912 23428 14940
rect 23584 14912 24716 14940
rect 25275 14912 25320 14940
rect 22511 14909 22523 14912
rect 22465 14903 22523 14909
rect 17862 14872 17868 14884
rect 13872 14844 15424 14872
rect 17823 14844 17868 14872
rect 13872 14832 13878 14844
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 19334 14832 19340 14884
rect 19392 14872 19398 14884
rect 20732 14872 20760 14903
rect 23400 14881 23428 14912
rect 19392 14844 20760 14872
rect 23385 14875 23443 14881
rect 19392 14832 19398 14844
rect 23385 14841 23397 14875
rect 23431 14841 23443 14875
rect 24118 14872 24124 14884
rect 24079 14844 24124 14872
rect 23385 14835 23443 14841
rect 24118 14832 24124 14844
rect 24176 14832 24182 14884
rect 24688 14881 24716 14912
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 25501 14943 25559 14949
rect 25501 14909 25513 14943
rect 25547 14940 25559 14943
rect 26510 14940 26516 14952
rect 25547 14912 26516 14940
rect 25547 14909 25559 14912
rect 25501 14903 25559 14909
rect 26510 14900 26516 14912
rect 26568 14900 26574 14952
rect 33520 14940 33548 14971
rect 33594 14968 33600 15020
rect 33652 15008 33658 15020
rect 35544 15017 35572 15048
rect 34885 15011 34943 15017
rect 34885 15008 34897 15011
rect 33652 14980 34897 15008
rect 33652 14968 33658 14980
rect 34885 14977 34897 14980
rect 34931 14977 34943 15011
rect 34885 14971 34943 14977
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 14977 35587 15011
rect 35529 14971 35587 14977
rect 37182 14940 37188 14952
rect 33520 14912 37188 14940
rect 37182 14900 37188 14912
rect 37240 14900 37246 14952
rect 24673 14875 24731 14881
rect 24673 14841 24685 14875
rect 24719 14841 24731 14875
rect 33597 14875 33655 14881
rect 33597 14872 33609 14875
rect 24673 14835 24731 14841
rect 24780 14844 33609 14872
rect 12115 14776 12204 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13173 14807 13231 14813
rect 13173 14804 13185 14807
rect 13044 14776 13185 14804
rect 13044 14764 13050 14776
rect 13173 14773 13185 14776
rect 13219 14773 13231 14807
rect 13173 14767 13231 14773
rect 17494 14764 17500 14816
rect 17552 14804 17558 14816
rect 20714 14804 20720 14816
rect 17552 14776 20720 14804
rect 17552 14764 17558 14776
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 20901 14807 20959 14813
rect 20901 14804 20913 14807
rect 20864 14776 20913 14804
rect 20864 14764 20870 14776
rect 20901 14773 20913 14776
rect 20947 14773 20959 14807
rect 20901 14767 20959 14773
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 24780 14804 24808 14844
rect 33597 14841 33609 14844
rect 33643 14841 33655 14875
rect 33597 14835 33655 14841
rect 23348 14776 24808 14804
rect 23348 14764 23354 14776
rect 25222 14764 25228 14816
rect 25280 14804 25286 14816
rect 25685 14807 25743 14813
rect 25685 14804 25697 14807
rect 25280 14776 25697 14804
rect 25280 14764 25286 14776
rect 25685 14773 25697 14776
rect 25731 14773 25743 14807
rect 25685 14767 25743 14773
rect 35345 14807 35403 14813
rect 35345 14773 35357 14807
rect 35391 14804 35403 14807
rect 38010 14804 38016 14816
rect 35391 14776 38016 14804
rect 35391 14773 35403 14776
rect 35345 14767 35403 14773
rect 38010 14764 38016 14776
rect 38068 14764 38074 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 6270 14600 6276 14612
rect 3467 14572 6276 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6365 14603 6423 14609
rect 6365 14569 6377 14603
rect 6411 14600 6423 14603
rect 9122 14600 9128 14612
rect 6411 14572 9128 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 12618 14600 12624 14612
rect 10100 14572 12624 14600
rect 10100 14560 10106 14572
rect 12618 14560 12624 14572
rect 12676 14600 12682 14612
rect 13722 14600 13728 14612
rect 12676 14572 13728 14600
rect 12676 14560 12682 14572
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 15562 14560 15568 14612
rect 15620 14600 15626 14612
rect 15620 14572 15665 14600
rect 15620 14560 15626 14572
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 17494 14600 17500 14612
rect 15988 14572 17500 14600
rect 15988 14560 15994 14572
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 18196 14572 18429 14600
rect 18196 14560 18202 14572
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 30009 14603 30067 14609
rect 18417 14563 18475 14569
rect 19076 14572 29960 14600
rect 3789 14535 3847 14541
rect 3789 14501 3801 14535
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2682 14464 2688 14476
rect 1995 14436 2688 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 3804 14464 3832 14495
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 8168 14504 9260 14532
rect 8168 14492 8174 14504
rect 8386 14464 8392 14476
rect 3804 14436 8392 14464
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 9088 14436 9137 14464
rect 9088 14424 9094 14436
rect 9125 14433 9137 14436
rect 9171 14433 9183 14467
rect 9232 14464 9260 14504
rect 10502 14492 10508 14544
rect 10560 14492 10566 14544
rect 10594 14492 10600 14544
rect 10652 14532 10658 14544
rect 13262 14532 13268 14544
rect 10652 14504 13268 14532
rect 10652 14492 10658 14504
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 14645 14535 14703 14541
rect 14645 14532 14657 14535
rect 13372 14504 14657 14532
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 9232 14436 9413 14464
rect 9125 14427 9183 14433
rect 9401 14433 9413 14436
rect 9447 14464 9459 14467
rect 10520 14464 10548 14492
rect 9447 14436 10548 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 10778 14424 10784 14476
rect 10836 14464 10842 14476
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 10836 14436 10885 14464
rect 10836 14424 10842 14436
rect 10873 14433 10885 14436
rect 10919 14433 10931 14467
rect 10873 14427 10931 14433
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14464 11483 14467
rect 12710 14464 12716 14476
rect 11471 14436 12716 14464
rect 11471 14433 11483 14436
rect 11425 14427 11483 14433
rect 12710 14424 12716 14436
rect 12768 14464 12774 14476
rect 13372 14464 13400 14504
rect 14645 14501 14657 14504
rect 14691 14501 14703 14535
rect 19076 14532 19104 14572
rect 25222 14532 25228 14544
rect 14645 14495 14703 14501
rect 16776 14504 19104 14532
rect 19168 14504 24900 14532
rect 25183 14504 25228 14532
rect 12768 14436 13400 14464
rect 13633 14467 13691 14473
rect 12768 14424 12774 14436
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 13814 14464 13820 14476
rect 13679 14436 13820 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14461 14467 14519 14473
rect 14461 14464 14473 14467
rect 13964 14436 14473 14464
rect 13964 14424 13970 14436
rect 14461 14433 14473 14436
rect 14507 14433 14519 14467
rect 15562 14464 15568 14476
rect 14461 14427 14519 14433
rect 15028 14436 15568 14464
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4062 14356 4068 14408
rect 4120 14396 4126 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4120 14368 4629 14396
rect 4120 14356 4126 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6788 14368 6837 14396
rect 6788 14356 6794 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12952 14368 13001 14396
rect 12952 14356 12958 14368
rect 12989 14365 13001 14368
rect 13035 14365 13047 14399
rect 13170 14396 13176 14408
rect 13131 14368 13176 14396
rect 12989 14359 13047 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14396 14335 14399
rect 15028 14396 15056 14436
rect 15562 14424 15568 14436
rect 15620 14464 15626 14476
rect 16022 14464 16028 14476
rect 15620 14436 16028 14464
rect 15620 14424 15626 14436
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 16132 14473 16344 14476
rect 16117 14467 16344 14473
rect 16117 14433 16129 14467
rect 16163 14464 16344 14467
rect 16776 14464 16804 14504
rect 16163 14448 16804 14464
rect 16163 14433 16175 14448
rect 16316 14436 16804 14448
rect 16117 14427 16175 14433
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 17313 14467 17371 14473
rect 17313 14464 17325 14467
rect 16908 14436 17325 14464
rect 16908 14424 16914 14436
rect 17313 14433 17325 14436
rect 17359 14433 17371 14467
rect 17313 14427 17371 14433
rect 17586 14424 17592 14476
rect 17644 14464 17650 14476
rect 17773 14467 17831 14473
rect 17773 14464 17785 14467
rect 17644 14436 17785 14464
rect 17644 14424 17650 14436
rect 17773 14433 17785 14436
rect 17819 14464 17831 14467
rect 19168 14464 19196 14504
rect 17819 14436 19196 14464
rect 17819 14433 17831 14436
rect 17773 14427 17831 14433
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19521 14467 19579 14473
rect 19521 14464 19533 14467
rect 19484 14436 19533 14464
rect 19484 14424 19490 14436
rect 19521 14433 19533 14436
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 20312 14436 20637 14464
rect 20312 14424 20318 14436
rect 20625 14433 20637 14436
rect 20671 14433 20683 14467
rect 20625 14427 20683 14433
rect 21266 14424 21272 14476
rect 21324 14464 21330 14476
rect 21729 14467 21787 14473
rect 21729 14464 21741 14467
rect 21324 14436 21741 14464
rect 21324 14424 21330 14436
rect 21729 14433 21741 14436
rect 21775 14433 21787 14467
rect 21729 14427 21787 14433
rect 22554 14424 22560 14476
rect 22612 14464 22618 14476
rect 23017 14467 23075 14473
rect 23017 14464 23029 14467
rect 22612 14436 23029 14464
rect 22612 14424 22618 14436
rect 23017 14433 23029 14436
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 23201 14467 23259 14473
rect 23201 14433 23213 14467
rect 23247 14464 23259 14467
rect 24670 14464 24676 14476
rect 23247 14436 24676 14464
rect 23247 14433 23259 14436
rect 23201 14427 23259 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 15470 14396 15476 14408
rect 14323 14368 15056 14396
rect 15431 14368 15476 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 16574 14396 16580 14408
rect 16347 14368 16580 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 18601 14399 18659 14405
rect 18601 14365 18613 14399
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14396 21971 14399
rect 22094 14396 22100 14408
rect 21959 14368 22100 14396
rect 21959 14365 21971 14368
rect 21913 14359 21971 14365
rect 2958 14288 2964 14340
rect 3016 14288 3022 14340
rect 4341 14331 4399 14337
rect 4341 14297 4353 14331
rect 4387 14328 4399 14331
rect 4522 14328 4528 14340
rect 4387 14300 4528 14328
rect 4387 14297 4399 14300
rect 4341 14291 4399 14297
rect 4522 14288 4528 14300
rect 4580 14328 4586 14340
rect 4893 14331 4951 14337
rect 4893 14328 4905 14331
rect 4580 14300 4905 14328
rect 4580 14288 4586 14300
rect 4893 14297 4905 14300
rect 4939 14297 4951 14331
rect 4893 14291 4951 14297
rect 5442 14288 5448 14340
rect 5500 14288 5506 14340
rect 7101 14331 7159 14337
rect 7101 14297 7113 14331
rect 7147 14328 7159 14331
rect 7190 14328 7196 14340
rect 7147 14300 7196 14328
rect 7147 14297 7159 14300
rect 7101 14291 7159 14297
rect 7190 14288 7196 14300
rect 7248 14288 7254 14340
rect 9306 14328 9312 14340
rect 7300 14300 7590 14328
rect 8496 14300 9312 14328
rect 7300 14272 7328 14300
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 7006 14260 7012 14272
rect 4856 14232 7012 14260
rect 4856 14220 4862 14232
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7282 14220 7288 14272
rect 7340 14220 7346 14272
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 8496 14260 8524 14300
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 9732 14300 9890 14328
rect 9732 14288 9738 14300
rect 11514 14288 11520 14340
rect 11572 14328 11578 14340
rect 12066 14328 12072 14340
rect 11572 14300 11617 14328
rect 12027 14300 12072 14328
rect 11572 14288 11578 14300
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 13078 14288 13084 14340
rect 13136 14328 13142 14340
rect 16022 14328 16028 14340
rect 13136 14300 16028 14328
rect 13136 14288 13142 14300
rect 16022 14288 16028 14300
rect 16080 14288 16086 14340
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 16724 14300 17356 14328
rect 16724 14288 16730 14300
rect 7432 14232 8524 14260
rect 8573 14263 8631 14269
rect 7432 14220 7438 14232
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 8662 14260 8668 14272
rect 8619 14232 8668 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 15930 14260 15936 14272
rect 9548 14232 15936 14260
rect 9548 14220 9554 14232
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16758 14260 16764 14272
rect 16719 14232 16764 14260
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 17328 14260 17356 14300
rect 17402 14288 17408 14340
rect 17460 14328 17466 14340
rect 17460 14300 17505 14328
rect 17460 14288 17466 14300
rect 18616 14260 18644 14359
rect 22094 14356 22100 14368
rect 22152 14356 22158 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 23860 14368 24593 14396
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 20622 14328 20628 14340
rect 20312 14300 20628 14328
rect 20312 14288 20318 14300
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 20714 14288 20720 14340
rect 20772 14328 20778 14340
rect 21269 14331 21327 14337
rect 20772 14300 20817 14328
rect 20772 14288 20778 14300
rect 21269 14297 21281 14331
rect 21315 14328 21327 14331
rect 21542 14328 21548 14340
rect 21315 14300 21548 14328
rect 21315 14297 21327 14300
rect 21269 14291 21327 14297
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 23860 14272 23888 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24765 14399 24823 14405
rect 24765 14396 24777 14399
rect 24581 14359 24639 14365
rect 24688 14368 24777 14396
rect 17328 14232 18644 14260
rect 22373 14263 22431 14269
rect 22373 14229 22385 14263
rect 22419 14260 22431 14263
rect 23106 14260 23112 14272
rect 22419 14232 23112 14260
rect 22419 14229 22431 14232
rect 22373 14223 22431 14229
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 23661 14263 23719 14269
rect 23661 14229 23673 14263
rect 23707 14260 23719 14263
rect 23842 14260 23848 14272
rect 23707 14232 23848 14260
rect 23707 14229 23719 14232
rect 23661 14223 23719 14229
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 24688 14260 24716 14368
rect 24765 14365 24777 14368
rect 24811 14365 24823 14399
rect 24765 14359 24823 14365
rect 24872 14328 24900 14504
rect 25222 14492 25228 14504
rect 25280 14492 25286 14544
rect 25314 14492 25320 14544
rect 25372 14532 25378 14544
rect 26053 14535 26111 14541
rect 26053 14532 26065 14535
rect 25372 14504 26065 14532
rect 25372 14492 25378 14504
rect 26053 14501 26065 14504
rect 26099 14501 26111 14535
rect 26053 14495 26111 14501
rect 26206 14504 29316 14532
rect 25958 14424 25964 14476
rect 26016 14464 26022 14476
rect 26206 14464 26234 14504
rect 26016 14436 26234 14464
rect 26016 14424 26022 14436
rect 26326 14424 26332 14476
rect 26384 14464 26390 14476
rect 27798 14464 27804 14476
rect 26384 14436 27804 14464
rect 26384 14424 26390 14436
rect 27798 14424 27804 14436
rect 27856 14424 27862 14476
rect 25682 14356 25688 14408
rect 25740 14396 25746 14408
rect 25869 14399 25927 14405
rect 25740 14368 25785 14396
rect 25740 14356 25746 14368
rect 25869 14365 25881 14399
rect 25915 14396 25927 14399
rect 26970 14396 26976 14408
rect 25915 14368 26556 14396
rect 26931 14368 26976 14396
rect 25915 14365 25927 14368
rect 25869 14359 25927 14365
rect 26234 14328 26240 14340
rect 24872 14300 26240 14328
rect 26234 14288 26240 14300
rect 26292 14288 26298 14340
rect 25866 14260 25872 14272
rect 24688 14232 25872 14260
rect 25866 14220 25872 14232
rect 25924 14220 25930 14272
rect 26528 14260 26556 14368
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 29288 14328 29316 14504
rect 29932 14464 29960 14572
rect 30009 14569 30021 14603
rect 30055 14600 30067 14603
rect 33594 14600 33600 14612
rect 30055 14572 33600 14600
rect 30055 14569 30067 14572
rect 30009 14563 30067 14569
rect 33594 14560 33600 14572
rect 33652 14560 33658 14612
rect 33781 14467 33839 14473
rect 33781 14464 33793 14467
rect 29932 14436 33793 14464
rect 33781 14433 33793 14436
rect 33827 14433 33839 14467
rect 33781 14427 33839 14433
rect 29914 14396 29920 14408
rect 29875 14368 29920 14396
rect 29914 14356 29920 14368
rect 29972 14356 29978 14408
rect 33689 14399 33747 14405
rect 33689 14365 33701 14399
rect 33735 14396 33747 14399
rect 38286 14396 38292 14408
rect 33735 14368 35894 14396
rect 38247 14368 38292 14396
rect 33735 14365 33747 14368
rect 33689 14359 33747 14365
rect 32398 14328 32404 14340
rect 29288 14300 32404 14328
rect 32398 14288 32404 14300
rect 32456 14288 32462 14340
rect 26789 14263 26847 14269
rect 26789 14260 26801 14263
rect 26528 14232 26801 14260
rect 26789 14229 26801 14232
rect 26835 14229 26847 14263
rect 35866 14260 35894 14368
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 38105 14263 38163 14269
rect 38105 14260 38117 14263
rect 35866 14232 38117 14260
rect 26789 14223 26847 14229
rect 38105 14229 38117 14232
rect 38151 14229 38163 14263
rect 38105 14223 38163 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1673 14059 1731 14065
rect 1673 14025 1685 14059
rect 1719 14056 1731 14059
rect 5166 14056 5172 14068
rect 1719 14028 5172 14056
rect 1719 14025 1731 14028
rect 1673 14019 1731 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5813 14059 5871 14065
rect 5813 14025 5825 14059
rect 5859 14056 5871 14059
rect 7374 14056 7380 14068
rect 5859 14028 7380 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 7374 14016 7380 14028
rect 7432 14016 7438 14068
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 10042 14056 10048 14068
rect 7607 14028 10048 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 13136 14028 13185 14056
rect 13136 14016 13142 14028
rect 13173 14025 13185 14028
rect 13219 14025 13231 14059
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 13173 14019 13231 14025
rect 13280 14028 15761 14056
rect 5534 13988 5540 14000
rect 4738 13960 5540 13988
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 8110 13988 8116 14000
rect 6012 13960 8116 13988
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1854 13920 1860 13932
rect 1544 13892 1860 13920
rect 1544 13880 1550 13892
rect 1854 13880 1860 13892
rect 1912 13920 1918 13932
rect 6012 13929 6040 13960
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 8754 13988 8760 14000
rect 8220 13960 8760 13988
rect 2317 13923 2375 13929
rect 2317 13920 2329 13923
rect 1912 13892 2329 13920
rect 1912 13880 1918 13892
rect 2317 13889 2329 13892
rect 2363 13889 2375 13923
rect 2317 13883 2375 13889
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 8220 13929 8248 13960
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 8938 13948 8944 14000
rect 8996 13948 9002 14000
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 12345 13991 12403 13997
rect 12345 13988 12357 13991
rect 9824 13960 12357 13988
rect 9824 13948 9830 13960
rect 12345 13957 12357 13960
rect 12391 13988 12403 13991
rect 12986 13988 12992 14000
rect 12391 13960 12992 13988
rect 12391 13957 12403 13960
rect 12345 13951 12403 13957
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 6788 13892 8217 13920
rect 6788 13880 6794 13892
rect 8205 13889 8217 13892
rect 8251 13889 8263 13923
rect 8205 13883 8263 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 13280 13920 13308 14028
rect 15749 14025 15761 14028
rect 15795 14056 15807 14059
rect 16758 14056 16764 14068
rect 15795 14028 16764 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17828 14028 18153 14056
rect 17828 14016 17834 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19429 14059 19487 14065
rect 19429 14056 19441 14059
rect 19392 14028 19441 14056
rect 19392 14016 19398 14028
rect 19429 14025 19441 14028
rect 19475 14025 19487 14059
rect 20070 14056 20076 14068
rect 20031 14028 20076 14056
rect 19429 14019 19487 14025
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 22094 14056 22100 14068
rect 20732 14028 21036 14056
rect 22055 14028 22100 14056
rect 13722 13948 13728 14000
rect 13780 13988 13786 14000
rect 13909 13991 13967 13997
rect 13909 13988 13921 13991
rect 13780 13960 13921 13988
rect 13780 13948 13786 13960
rect 13909 13957 13921 13960
rect 13955 13957 13967 13991
rect 13909 13951 13967 13957
rect 14001 13991 14059 13997
rect 14001 13957 14013 13991
rect 14047 13988 14059 13991
rect 14182 13988 14188 14000
rect 14047 13960 14188 13988
rect 14047 13957 14059 13960
rect 14001 13951 14059 13957
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 14553 13991 14611 13997
rect 14553 13957 14565 13991
rect 14599 13988 14611 13991
rect 16666 13988 16672 14000
rect 14599 13960 16672 13988
rect 14599 13957 14611 13960
rect 14553 13951 14611 13957
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 17034 13988 17040 14000
rect 16995 13960 17040 13988
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 17586 13988 17592 14000
rect 17547 13960 17592 13988
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 20732 13988 20760 14028
rect 20898 13988 20904 14000
rect 19628 13960 20760 13988
rect 20859 13960 20904 13988
rect 10551 13892 13308 13920
rect 13357 13923 13415 13929
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13821 2559 13855
rect 2501 13815 2559 13821
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3510 13852 3516 13864
rect 3283 13824 3372 13852
rect 3471 13824 3516 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 2314 13744 2320 13796
rect 2372 13784 2378 13796
rect 2516 13784 2544 13815
rect 2372 13756 2544 13784
rect 2372 13744 2378 13756
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 2958 13716 2964 13728
rect 1820 13688 2964 13716
rect 1820 13676 1826 13688
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 3344 13716 3372 13824
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 4706 13812 4712 13864
rect 4764 13852 4770 13864
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 4764 13824 5273 13852
rect 4764 13812 4770 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 5261 13815 5319 13821
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6420 13824 6929 13852
rect 6420 13812 6426 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 7064 13824 7113 13852
rect 7064 13812 7070 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8536 13824 8581 13852
rect 8536 13812 8542 13824
rect 9674 13812 9680 13864
rect 9732 13852 9738 13864
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9732 13824 9965 13852
rect 9732 13812 9738 13824
rect 9953 13821 9965 13824
rect 9999 13821 10011 13855
rect 9953 13815 10011 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 11054 13852 11060 13864
rect 10735 13824 11060 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11480 13824 11713 13852
rect 11480 13812 11486 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12802 13852 12808 13864
rect 11931 13824 12808 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13372 13852 13400 13883
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 18322 13920 18328 13932
rect 14792 13892 16252 13920
rect 18283 13892 18328 13920
rect 14792 13880 14798 13892
rect 14918 13852 14924 13864
rect 13372 13824 14924 13852
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15102 13852 15108 13864
rect 15063 13824 15108 13852
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 16114 13852 16120 13864
rect 15335 13824 16120 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 16114 13812 16120 13824
rect 16172 13812 16178 13864
rect 16224 13852 16252 13892
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18782 13920 18788 13932
rect 18743 13892 18788 13920
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 19628 13929 19656 13960
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 21008 13988 21036 14028
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 23842 14056 23848 14068
rect 23803 14028 23848 14056
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 25314 14056 25320 14068
rect 25275 14028 25320 14056
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 26510 14056 26516 14068
rect 26471 14028 26516 14056
rect 26510 14016 26516 14028
rect 26568 14016 26574 14068
rect 22554 13988 22560 14000
rect 21008 13960 22560 13988
rect 22554 13948 22560 13960
rect 22612 13948 22618 14000
rect 25222 13948 25228 14000
rect 25280 13988 25286 14000
rect 29914 13988 29920 14000
rect 25280 13960 29920 13988
rect 25280 13948 25286 13960
rect 29914 13948 29920 13960
rect 29972 13948 29978 14000
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 22278 13920 22284 13932
rect 22239 13892 22284 13920
rect 19613 13883 19671 13889
rect 22278 13880 22284 13892
rect 22336 13880 22342 13932
rect 23201 13923 23259 13929
rect 23201 13889 23213 13923
rect 23247 13920 23259 13923
rect 24578 13920 24584 13932
rect 23247 13892 24584 13920
rect 23247 13889 23259 13892
rect 23201 13883 23259 13889
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 25774 13920 25780 13932
rect 25735 13892 25780 13920
rect 25774 13880 25780 13892
rect 25832 13880 25838 13932
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26421 13923 26479 13929
rect 26421 13920 26433 13923
rect 26292 13892 26433 13920
rect 26292 13880 26298 13892
rect 26421 13889 26433 13892
rect 26467 13889 26479 13923
rect 26421 13883 26479 13889
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 16224 13824 16957 13852
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 16945 13815 17003 13821
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 20162 13852 20168 13864
rect 18923 13824 20168 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20806 13852 20812 13864
rect 20767 13824 20812 13852
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 21453 13855 21511 13861
rect 21453 13821 21465 13855
rect 21499 13852 21511 13855
rect 22186 13852 22192 13864
rect 21499 13824 22192 13852
rect 21499 13821 21511 13824
rect 21453 13815 21511 13821
rect 22186 13812 22192 13824
rect 22244 13852 22250 13864
rect 22830 13852 22836 13864
rect 22244 13824 22836 13852
rect 22244 13812 22250 13824
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 23385 13855 23443 13861
rect 23385 13821 23397 13855
rect 23431 13852 23443 13855
rect 24210 13852 24216 13864
rect 23431 13824 24216 13852
rect 23431 13821 23443 13824
rect 23385 13815 23443 13821
rect 24210 13812 24216 13824
rect 24268 13812 24274 13864
rect 24670 13852 24676 13864
rect 24631 13824 24676 13852
rect 24670 13812 24676 13824
rect 24728 13812 24734 13864
rect 24857 13855 24915 13861
rect 24857 13821 24869 13855
rect 24903 13852 24915 13855
rect 25869 13855 25927 13861
rect 25869 13852 25881 13855
rect 24903 13824 25881 13852
rect 24903 13821 24915 13824
rect 24857 13815 24915 13821
rect 25869 13821 25881 13824
rect 25915 13821 25927 13855
rect 25869 13815 25927 13821
rect 9508 13756 14412 13784
rect 4062 13716 4068 13728
rect 3344 13688 4068 13716
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 9508 13716 9536 13756
rect 4764 13688 9536 13716
rect 4764 13676 4770 13688
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 10318 13716 10324 13728
rect 9732 13688 10324 13716
rect 9732 13676 9738 13688
rect 10318 13676 10324 13688
rect 10376 13716 10382 13728
rect 11146 13716 11152 13728
rect 10376 13688 11152 13716
rect 10376 13676 10382 13688
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 12618 13716 12624 13728
rect 11296 13688 12624 13716
rect 11296 13676 11302 13688
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 14384 13716 14412 13756
rect 14568 13756 17264 13784
rect 14568 13716 14596 13756
rect 14384 13688 14596 13716
rect 14642 13676 14648 13728
rect 14700 13716 14706 13728
rect 16758 13716 16764 13728
rect 14700 13688 16764 13716
rect 14700 13676 14706 13688
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 17236 13716 17264 13756
rect 17604 13756 25452 13784
rect 17604 13716 17632 13756
rect 17236 13688 17632 13716
rect 25424 13716 25452 13756
rect 26234 13716 26240 13728
rect 25424 13688 26240 13716
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 3418 13512 3424 13524
rect 3379 13484 3424 13512
rect 3418 13472 3424 13484
rect 3476 13512 3482 13524
rect 3602 13512 3608 13524
rect 3476 13484 3608 13512
rect 3476 13472 3482 13484
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 4236 13515 4294 13521
rect 4236 13481 4248 13515
rect 4282 13512 4294 13515
rect 4706 13512 4712 13524
rect 4282 13484 4712 13512
rect 4282 13481 4294 13484
rect 4236 13475 4294 13481
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 11238 13512 11244 13524
rect 6656 13484 11244 13512
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 6656 13376 6684 13484
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 13354 13512 13360 13524
rect 11348 13484 13360 13512
rect 8588 13416 9260 13444
rect 1995 13348 6684 13376
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 7009 13379 7067 13385
rect 6788 13348 6833 13376
rect 6788 13336 6794 13348
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 8478 13376 8484 13388
rect 7055 13348 8484 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 3970 13308 3976 13320
rect 3931 13280 3976 13308
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 8588 13308 8616 13416
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9125 13379 9183 13385
rect 9125 13376 9137 13379
rect 9088 13348 9137 13376
rect 9088 13336 9094 13348
rect 9125 13345 9137 13348
rect 9171 13345 9183 13379
rect 9232 13376 9260 13416
rect 11348 13385 11376 13484
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 13630 13512 13636 13524
rect 13591 13484 13636 13512
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14734 13512 14740 13524
rect 14695 13484 14740 13512
rect 14734 13472 14740 13484
rect 14792 13512 14798 13524
rect 14918 13512 14924 13524
rect 14792 13484 14924 13512
rect 14792 13472 14798 13484
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 15657 13515 15715 13521
rect 15657 13481 15669 13515
rect 15703 13512 15715 13515
rect 17034 13512 17040 13524
rect 15703 13484 17040 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 20898 13472 20904 13524
rect 20956 13512 20962 13524
rect 21913 13515 21971 13521
rect 21913 13512 21925 13515
rect 20956 13484 21925 13512
rect 20956 13472 20962 13484
rect 21913 13481 21925 13484
rect 21959 13481 21971 13515
rect 22554 13512 22560 13524
rect 22515 13484 22560 13512
rect 21913 13475 21971 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 25866 13512 25872 13524
rect 25827 13484 25872 13512
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 26513 13515 26571 13521
rect 26513 13481 26525 13515
rect 26559 13512 26571 13515
rect 26970 13512 26976 13524
rect 26559 13484 26976 13512
rect 26559 13481 26571 13484
rect 26513 13475 26571 13481
rect 26970 13472 26976 13484
rect 27028 13472 27034 13524
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 13446 13444 13452 13456
rect 11664 13416 13452 13444
rect 11664 13404 11670 13416
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 13722 13404 13728 13456
rect 13780 13444 13786 13456
rect 14642 13444 14648 13456
rect 13780 13416 14648 13444
rect 13780 13404 13786 13416
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 14826 13404 14832 13456
rect 14884 13444 14890 13456
rect 17405 13447 17463 13453
rect 17405 13444 17417 13447
rect 14884 13416 17417 13444
rect 14884 13404 14890 13416
rect 17405 13413 17417 13416
rect 17451 13413 17463 13447
rect 17405 13407 17463 13413
rect 18877 13447 18935 13453
rect 18877 13413 18889 13447
rect 18923 13444 18935 13447
rect 19797 13447 19855 13453
rect 19797 13444 19809 13447
rect 18923 13416 19809 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 19797 13413 19809 13416
rect 19843 13444 19855 13447
rect 20070 13444 20076 13456
rect 19843 13416 20076 13444
rect 19843 13413 19855 13416
rect 19797 13407 19855 13413
rect 20070 13404 20076 13416
rect 20128 13404 20134 13456
rect 20990 13404 20996 13456
rect 21048 13444 21054 13456
rect 21358 13444 21364 13456
rect 21048 13416 21364 13444
rect 21048 13404 21054 13416
rect 21358 13404 21364 13416
rect 21416 13404 21422 13456
rect 27982 13444 27988 13456
rect 22066 13416 27988 13444
rect 11333 13379 11391 13385
rect 9232 13348 10640 13376
rect 9125 13339 9183 13345
rect 8312 13280 8616 13308
rect 10612 13308 10640 13348
rect 11333 13345 11345 13379
rect 11379 13345 11391 13379
rect 14277 13379 14335 13385
rect 11333 13339 11391 13345
rect 11440 13348 13768 13376
rect 11440 13308 11468 13348
rect 10612 13280 11468 13308
rect 11517 13311 11575 13317
rect 3694 13240 3700 13252
rect 3174 13212 3700 13240
rect 3694 13200 3700 13212
rect 3752 13200 3758 13252
rect 5718 13240 5724 13252
rect 5474 13212 5724 13240
rect 5718 13200 5724 13212
rect 5776 13200 5782 13252
rect 5997 13243 6055 13249
rect 5997 13209 6009 13243
rect 6043 13209 6055 13243
rect 5997 13203 6055 13209
rect 2958 13132 2964 13184
rect 3016 13172 3022 13184
rect 6012 13172 6040 13203
rect 7742 13200 7748 13252
rect 7800 13200 7806 13252
rect 8312 13172 8340 13280
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11698 13308 11704 13320
rect 11563 13280 11704 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11848 13280 11989 13308
rect 11848 13268 11854 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12400 13280 12449 13308
rect 12400 13268 12406 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12618 13308 12624 13320
rect 12579 13280 12624 13308
rect 12437 13271 12495 13277
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8846 13240 8852 13252
rect 8444 13212 8852 13240
rect 8444 13200 8450 13212
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 9398 13240 9404 13252
rect 9359 13212 9404 13240
rect 9398 13200 9404 13212
rect 9456 13200 9462 13252
rect 9950 13200 9956 13252
rect 10008 13200 10014 13252
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 13556 13240 13584 13268
rect 10836 13212 13584 13240
rect 13740 13240 13768 13348
rect 14277 13345 14289 13379
rect 14323 13376 14335 13379
rect 14734 13376 14740 13388
rect 14323 13348 14740 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 14734 13336 14740 13348
rect 14792 13376 14798 13388
rect 15102 13376 15108 13388
rect 14792 13348 15108 13376
rect 14792 13336 14798 13348
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 20162 13376 20168 13388
rect 15212 13348 20168 13376
rect 13998 13268 14004 13320
rect 14056 13308 14062 13320
rect 14182 13308 14188 13320
rect 14056 13280 14188 13308
rect 14056 13268 14062 13280
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14458 13308 14464 13320
rect 14419 13280 14464 13308
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15212 13240 15240 13348
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13376 20867 13379
rect 22066 13376 22094 13416
rect 27982 13404 27988 13416
rect 28040 13404 28046 13456
rect 20855 13348 22094 13376
rect 20855 13345 20867 13348
rect 20809 13339 20867 13345
rect 22922 13336 22928 13388
rect 22980 13376 22986 13388
rect 23293 13379 23351 13385
rect 23293 13376 23305 13379
rect 22980 13348 23305 13376
rect 22980 13336 22986 13348
rect 23293 13345 23305 13348
rect 23339 13345 23351 13379
rect 24578 13376 24584 13388
rect 24539 13348 24584 13376
rect 23293 13339 23351 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13308 15623 13311
rect 15654 13308 15660 13320
rect 15611 13280 15660 13308
rect 15611 13277 15623 13280
rect 15565 13271 15623 13277
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 17586 13308 17592 13320
rect 17547 13280 17592 13308
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 18230 13308 18236 13320
rect 18191 13280 18236 13308
rect 18230 13268 18236 13280
rect 18288 13268 18294 13320
rect 18414 13308 18420 13320
rect 18375 13280 18420 13308
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 19392 13280 19441 13308
rect 19392 13268 19398 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19518 13268 19524 13320
rect 19576 13308 19582 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19576 13280 19625 13308
rect 19576 13268 19582 13280
rect 19613 13277 19625 13280
rect 19659 13277 19671 13311
rect 19613 13271 19671 13277
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13308 21051 13311
rect 21082 13308 21088 13320
rect 21039 13280 21088 13308
rect 21039 13277 21051 13280
rect 20993 13271 21051 13277
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13277 22155 13311
rect 22738 13308 22744 13320
rect 22699 13280 22744 13308
rect 22097 13271 22155 13277
rect 13740 13212 15240 13240
rect 16301 13243 16359 13249
rect 10836 13200 10842 13212
rect 16301 13209 16313 13243
rect 16347 13209 16359 13243
rect 16301 13203 16359 13209
rect 3016 13144 8340 13172
rect 8481 13175 8539 13181
rect 3016 13132 3022 13144
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 9766 13172 9772 13184
rect 8527 13144 9772 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10192 13144 10885 13172
rect 10192 13132 10198 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 13078 13172 13084 13184
rect 13039 13144 13084 13172
rect 10873 13135 10931 13141
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 13446 13132 13452 13184
rect 13504 13172 13510 13184
rect 15470 13172 15476 13184
rect 13504 13144 15476 13172
rect 13504 13132 13510 13144
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 16316 13172 16344 13203
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 16448 13212 16493 13240
rect 16448 13200 16454 13212
rect 16666 13200 16672 13252
rect 16724 13240 16730 13252
rect 16945 13243 17003 13249
rect 16945 13240 16957 13243
rect 16724 13212 16957 13240
rect 16724 13200 16730 13212
rect 16945 13209 16957 13212
rect 16991 13240 17003 13243
rect 17034 13240 17040 13252
rect 16991 13212 17040 13240
rect 16991 13209 17003 13212
rect 16945 13203 17003 13209
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 22112 13240 22140 13271
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 25222 13268 25228 13320
rect 25280 13308 25286 13320
rect 25409 13311 25467 13317
rect 25409 13308 25421 13311
rect 25280 13280 25421 13308
rect 25280 13268 25286 13280
rect 25409 13277 25421 13280
rect 25455 13277 25467 13311
rect 25409 13271 25467 13277
rect 19116 13212 22140 13240
rect 23385 13243 23443 13249
rect 19116 13200 19122 13212
rect 23385 13209 23397 13243
rect 23431 13240 23443 13243
rect 23750 13240 23756 13252
rect 23431 13212 23756 13240
rect 23431 13209 23443 13212
rect 23385 13203 23443 13209
rect 23750 13200 23756 13212
rect 23808 13200 23814 13252
rect 23934 13240 23940 13252
rect 23895 13212 23940 13240
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 25424 13240 25452 13271
rect 25590 13268 25596 13320
rect 25648 13308 25654 13320
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 25648 13280 26065 13308
rect 25648 13268 25654 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26697 13311 26755 13317
rect 26697 13308 26709 13311
rect 26053 13271 26111 13277
rect 26206 13280 26709 13308
rect 25774 13240 25780 13252
rect 25424 13212 25780 13240
rect 25774 13200 25780 13212
rect 25832 13240 25838 13252
rect 26206 13240 26234 13280
rect 26697 13277 26709 13280
rect 26743 13277 26755 13311
rect 26697 13271 26755 13277
rect 25832 13212 26234 13240
rect 25832 13200 25838 13212
rect 16850 13172 16856 13184
rect 16316 13144 16856 13172
rect 16850 13132 16856 13144
rect 16908 13132 16914 13184
rect 24762 13132 24768 13184
rect 24820 13172 24826 13184
rect 25225 13175 25283 13181
rect 25225 13172 25237 13175
rect 24820 13144 25237 13172
rect 24820 13132 24826 13144
rect 25225 13141 25237 13144
rect 25271 13141 25283 13175
rect 25225 13135 25283 13141
rect 25314 13132 25320 13184
rect 25372 13172 25378 13184
rect 27246 13172 27252 13184
rect 25372 13144 27252 13172
rect 25372 13132 25378 13144
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 3694 12928 3700 12980
rect 3752 12968 3758 12980
rect 6086 12968 6092 12980
rect 3752 12940 6092 12968
rect 3752 12928 3758 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 10318 12968 10324 12980
rect 8444 12940 10324 12968
rect 8444 12928 8450 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 11330 12968 11336 12980
rect 10827 12940 11336 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 16206 12968 16212 12980
rect 11624 12940 16212 12968
rect 1854 12900 1860 12912
rect 1815 12872 1860 12900
rect 1854 12860 1860 12872
rect 1912 12860 1918 12912
rect 4338 12900 4344 12912
rect 3082 12872 3832 12900
rect 4299 12872 4344 12900
rect 3804 12776 3832 12872
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 6730 12900 6736 12912
rect 6564 12872 6736 12900
rect 6564 12844 6592 12872
rect 6730 12860 6736 12872
rect 6788 12860 6794 12912
rect 6825 12903 6883 12909
rect 6825 12869 6837 12903
rect 6871 12900 6883 12903
rect 6914 12900 6920 12912
rect 6871 12872 6920 12900
rect 6871 12869 6883 12872
rect 6825 12863 6883 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 7834 12860 7840 12912
rect 7892 12860 7898 12912
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 5442 12792 5448 12844
rect 5500 12792 5506 12844
rect 6546 12832 6552 12844
rect 6459 12804 6552 12832
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 8036 12804 9229 12832
rect 1578 12764 1584 12776
rect 1539 12736 1584 12764
rect 1578 12724 1584 12736
rect 1636 12724 1642 12776
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 2280 12736 3617 12764
rect 2280 12724 2286 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3620 12696 3648 12727
rect 3786 12724 3792 12776
rect 3844 12724 3850 12776
rect 6178 12764 6184 12776
rect 4172 12736 6184 12764
rect 4172 12696 4200 12736
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 7374 12764 7380 12776
rect 6656 12736 7380 12764
rect 5810 12696 5816 12708
rect 3620 12668 4200 12696
rect 5723 12668 5816 12696
rect 5810 12656 5816 12668
rect 5868 12696 5874 12708
rect 6656 12696 6684 12736
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 8036 12764 8064 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 10042 12832 10048 12844
rect 9548 12804 10048 12832
rect 9548 12792 9554 12804
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 11624 12832 11652 12940
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 16482 12928 16488 12980
rect 16540 12968 16546 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 16540 12940 16957 12968
rect 16540 12928 16546 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 18141 12971 18199 12977
rect 18141 12937 18153 12971
rect 18187 12968 18199 12971
rect 18322 12968 18328 12980
rect 18187 12940 18328 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 19058 12968 19064 12980
rect 19019 12940 19064 12968
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19797 12971 19855 12977
rect 19797 12937 19809 12971
rect 19843 12968 19855 12971
rect 19978 12968 19984 12980
rect 19843 12940 19984 12968
rect 19843 12937 19855 12940
rect 19797 12931 19855 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 21269 12971 21327 12977
rect 21269 12968 21281 12971
rect 20864 12940 21281 12968
rect 20864 12928 20870 12940
rect 21269 12937 21281 12940
rect 21315 12937 21327 12971
rect 21269 12931 21327 12937
rect 22278 12928 22284 12980
rect 22336 12968 22342 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 22336 12940 22385 12968
rect 22336 12928 22342 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 23566 12968 23572 12980
rect 22373 12931 22431 12937
rect 22940 12940 23572 12968
rect 12529 12903 12587 12909
rect 12529 12869 12541 12903
rect 12575 12900 12587 12903
rect 13630 12900 13636 12912
rect 12575 12872 13636 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 13725 12903 13783 12909
rect 13725 12869 13737 12903
rect 13771 12900 13783 12903
rect 14921 12903 14979 12909
rect 13771 12872 14872 12900
rect 13771 12869 13783 12872
rect 13725 12863 13783 12869
rect 10183 12804 11652 12832
rect 11701 12835 11759 12841
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 14844 12832 14872 12872
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 15194 12900 15200 12912
rect 14967 12872 15200 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 20162 12860 20168 12912
rect 20220 12900 20226 12912
rect 22940 12900 22968 12940
rect 23566 12928 23572 12940
rect 23624 12928 23630 12980
rect 24210 12968 24216 12980
rect 24171 12940 24216 12968
rect 24210 12928 24216 12940
rect 24268 12928 24274 12980
rect 25590 12968 25596 12980
rect 25551 12940 25596 12968
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 23106 12900 23112 12912
rect 20220 12872 22968 12900
rect 23067 12872 23112 12900
rect 20220 12860 20226 12872
rect 23106 12860 23112 12872
rect 23164 12860 23170 12912
rect 23201 12903 23259 12909
rect 23201 12869 23213 12903
rect 23247 12900 23259 12903
rect 24949 12903 25007 12909
rect 24949 12900 24961 12903
rect 23247 12872 24961 12900
rect 23247 12869 23259 12872
rect 23201 12863 23259 12869
rect 24949 12869 24961 12872
rect 24995 12869 25007 12903
rect 24949 12863 25007 12869
rect 15930 12832 15936 12844
rect 14844 12804 15936 12832
rect 11701 12795 11759 12801
rect 7616 12736 8064 12764
rect 7616 12724 7622 12736
rect 8110 12724 8116 12776
rect 8168 12764 8174 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 8168 12736 8309 12764
rect 8168 12724 8174 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 9030 12764 9036 12776
rect 8991 12736 9036 12764
rect 8297 12727 8355 12733
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 9364 12736 10333 12764
rect 9364 12724 9370 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11716 12764 11744 12795
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 18138 12792 18144 12844
rect 18196 12832 18202 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18196 12804 18337 12832
rect 18196 12792 18202 12804
rect 18325 12801 18337 12804
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 19245 12835 19303 12841
rect 19245 12832 19257 12835
rect 18564 12804 19257 12832
rect 18564 12792 18570 12804
rect 19245 12801 19257 12804
rect 19291 12832 19303 12835
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19291 12804 19717 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12832 20683 12835
rect 21358 12832 21364 12844
rect 20671 12804 21364 12832
rect 20671 12801 20683 12804
rect 20625 12795 20683 12801
rect 21358 12792 21364 12804
rect 21416 12792 21422 12844
rect 22554 12832 22560 12844
rect 22515 12804 22560 12832
rect 22554 12792 22560 12804
rect 22612 12792 22618 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24762 12832 24768 12844
rect 24443 12804 24768 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 25406 12832 25412 12844
rect 24903 12804 25412 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 25406 12792 25412 12804
rect 25464 12792 25470 12844
rect 25777 12835 25835 12841
rect 25777 12801 25789 12835
rect 25823 12832 25835 12835
rect 26234 12832 26240 12844
rect 25823 12804 26240 12832
rect 25823 12801 25835 12804
rect 25777 12795 25835 12801
rect 26234 12792 26240 12804
rect 26292 12792 26298 12844
rect 38010 12832 38016 12844
rect 37971 12804 38016 12832
rect 38010 12792 38016 12804
rect 38068 12792 38074 12844
rect 11204 12736 11744 12764
rect 12437 12767 12495 12773
rect 11204 12724 11210 12736
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 13633 12767 13691 12773
rect 12483 12736 12848 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 5868 12668 6684 12696
rect 7852 12668 10916 12696
rect 5868 12656 5874 12668
rect 6178 12588 6184 12640
rect 6236 12628 6242 12640
rect 7852 12628 7880 12668
rect 6236 12600 7880 12628
rect 6236 12588 6242 12600
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8110 12628 8116 12640
rect 7984 12600 8116 12628
rect 7984 12588 7990 12600
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8628 12600 9413 12628
rect 8628 12588 8634 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10778 12628 10784 12640
rect 9824 12600 10784 12628
rect 9824 12588 9830 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 10888 12628 10916 12668
rect 11606 12628 11612 12640
rect 10888 12600 11612 12628
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 12158 12628 12164 12640
rect 11839 12600 12164 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12820 12628 12848 12736
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 15194 12764 15200 12776
rect 13679 12736 15200 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15562 12764 15568 12776
rect 15475 12736 15568 12764
rect 15562 12724 15568 12736
rect 15620 12724 15626 12776
rect 15749 12767 15807 12773
rect 15749 12733 15761 12767
rect 15795 12764 15807 12767
rect 16758 12764 16764 12776
rect 15795 12736 16764 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 20806 12764 20812 12776
rect 20767 12736 20812 12764
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 23753 12767 23811 12773
rect 23753 12733 23765 12767
rect 23799 12764 23811 12767
rect 23934 12764 23940 12776
rect 23799 12736 23940 12764
rect 23799 12733 23811 12736
rect 23753 12727 23811 12733
rect 23934 12724 23940 12736
rect 23992 12764 23998 12776
rect 28258 12764 28264 12776
rect 23992 12736 28264 12764
rect 23992 12724 23998 12736
rect 28258 12724 28264 12736
rect 28316 12724 28322 12776
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12696 13047 12699
rect 13722 12696 13728 12708
rect 13035 12668 13728 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 14185 12699 14243 12705
rect 14185 12665 14197 12699
rect 14231 12696 14243 12699
rect 15010 12696 15016 12708
rect 14231 12668 15016 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 15580 12696 15608 12724
rect 25314 12696 25320 12708
rect 15580 12668 25320 12696
rect 25314 12656 25320 12668
rect 25372 12656 25378 12708
rect 13078 12628 13084 12640
rect 12820 12600 13084 12628
rect 13078 12588 13084 12600
rect 13136 12628 13142 12640
rect 15933 12631 15991 12637
rect 15933 12628 15945 12631
rect 13136 12600 15945 12628
rect 13136 12588 13142 12600
rect 15933 12597 15945 12600
rect 15979 12597 15991 12631
rect 15933 12591 15991 12597
rect 16206 12588 16212 12640
rect 16264 12628 16270 12640
rect 21174 12628 21180 12640
rect 16264 12600 21180 12628
rect 16264 12588 16270 12600
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 3418 12424 3424 12436
rect 2188 12396 3280 12424
rect 3379 12396 3424 12424
rect 2188 12384 2194 12396
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2038 12288 2044 12300
rect 1995 12260 2044 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3252 12288 3280 12396
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4065 12427 4123 12433
rect 4065 12393 4077 12427
rect 4111 12424 4123 12427
rect 7466 12424 7472 12436
rect 4111 12396 7472 12424
rect 4111 12393 4123 12396
rect 4065 12387 4123 12393
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 10686 12424 10692 12436
rect 7760 12396 10692 12424
rect 3200 12260 3280 12288
rect 3200 12248 3206 12260
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 3252 12220 3280 12260
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 4709 12291 4767 12297
rect 3660 12260 4108 12288
rect 3660 12248 3666 12260
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3252 12192 3985 12220
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 3174 12124 3924 12152
rect 3896 12096 3924 12124
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 4080 12084 4108 12260
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 5534 12288 5540 12300
rect 4755 12260 5540 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 5534 12248 5540 12260
rect 5592 12288 5598 12300
rect 6546 12288 6552 12300
rect 5592 12260 6552 12288
rect 5592 12248 5598 12260
rect 6546 12248 6552 12260
rect 6604 12248 6610 12300
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 6822 12288 6828 12300
rect 6779 12260 6828 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12288 7343 12291
rect 7760 12288 7788 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 16482 12424 16488 12436
rect 10796 12396 16488 12424
rect 8110 12316 8116 12368
rect 8168 12316 8174 12368
rect 8573 12359 8631 12365
rect 8573 12325 8585 12359
rect 8619 12356 8631 12359
rect 9030 12356 9036 12368
rect 8619 12328 9036 12356
rect 8619 12325 8631 12328
rect 8573 12319 8631 12325
rect 9030 12316 9036 12328
rect 9088 12356 9094 12368
rect 10413 12359 10471 12365
rect 10413 12356 10425 12359
rect 9088 12328 10425 12356
rect 9088 12316 9094 12328
rect 10413 12325 10425 12328
rect 10459 12325 10471 12359
rect 10413 12319 10471 12325
rect 10594 12316 10600 12368
rect 10652 12356 10658 12368
rect 10796 12356 10824 12396
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16761 12427 16819 12433
rect 16761 12424 16773 12427
rect 16632 12396 16773 12424
rect 16632 12384 16638 12396
rect 16761 12393 16773 12396
rect 16807 12393 16819 12427
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 16761 12387 16819 12393
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 20165 12427 20223 12433
rect 17972 12396 18184 12424
rect 10652 12328 10824 12356
rect 10652 12316 10658 12328
rect 11422 12316 11428 12368
rect 11480 12356 11486 12368
rect 11517 12359 11575 12365
rect 11517 12356 11529 12359
rect 11480 12328 11529 12356
rect 11480 12316 11486 12328
rect 11517 12325 11529 12328
rect 11563 12325 11575 12359
rect 11517 12319 11575 12325
rect 12526 12316 12532 12368
rect 12584 12356 12590 12368
rect 12710 12356 12716 12368
rect 12584 12328 12716 12356
rect 12584 12316 12590 12328
rect 12710 12316 12716 12328
rect 12768 12316 12774 12368
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16942 12356 16948 12368
rect 16071 12328 16948 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16942 12316 16948 12328
rect 17000 12316 17006 12368
rect 17310 12316 17316 12368
rect 17368 12356 17374 12368
rect 17972 12356 18000 12396
rect 17368 12328 18000 12356
rect 18049 12359 18107 12365
rect 17368 12316 17374 12328
rect 18049 12325 18061 12359
rect 18095 12325 18107 12359
rect 18049 12319 18107 12325
rect 7331 12260 7788 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8128 12288 8156 12316
rect 7975 12260 8156 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 8444 12260 10057 12288
rect 8444 12248 8450 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10502 12288 10508 12300
rect 10045 12251 10103 12257
rect 10152 12260 10508 12288
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7852 12220 7880 12248
rect 8110 12220 8116 12232
rect 7248 12192 7880 12220
rect 8071 12192 8116 12220
rect 7248 12180 7254 12192
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 9490 12220 9496 12232
rect 8220 12192 9496 12220
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4672 12124 4997 12152
rect 4672 12112 4678 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 6270 12152 6276 12164
rect 6210 12124 6276 12152
rect 4985 12115 5043 12121
rect 6270 12112 6276 12124
rect 6328 12112 6334 12164
rect 8220 12152 8248 12192
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 10152 12222 10180 12260
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 14734 12288 14740 12300
rect 11195 12260 14740 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 10060 12220 10180 12222
rect 9631 12194 10180 12220
rect 10229 12223 10287 12229
rect 9631 12192 10088 12194
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 12342 12220 12348 12232
rect 11379 12192 12348 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 6380 12124 8248 12152
rect 6380 12084 6408 12124
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 10042 12152 10048 12164
rect 8720 12124 10048 12152
rect 8720 12112 8726 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10245 12152 10273 12183
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12526 12220 12532 12232
rect 12487 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 13780 12192 13825 12220
rect 13780 12180 13786 12192
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 16080 12192 16221 12220
rect 16080 12180 16086 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16666 12220 16672 12232
rect 16579 12192 16672 12220
rect 16209 12183 16267 12189
rect 16666 12180 16672 12192
rect 16724 12220 16730 12232
rect 17494 12220 17500 12232
rect 16724 12192 17500 12220
rect 16724 12180 16730 12192
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 18064 12220 18092 12319
rect 17635 12192 18092 12220
rect 18156 12220 18184 12396
rect 20165 12393 20177 12427
rect 20211 12424 20223 12427
rect 21082 12424 21088 12436
rect 20211 12396 21088 12424
rect 20211 12393 20223 12396
rect 20165 12387 20223 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 23017 12427 23075 12433
rect 23017 12393 23029 12427
rect 23063 12424 23075 12427
rect 23106 12424 23112 12436
rect 23063 12396 23112 12424
rect 23063 12393 23075 12396
rect 23017 12387 23075 12393
rect 23106 12384 23112 12396
rect 23164 12384 23170 12436
rect 23750 12384 23756 12436
rect 23808 12424 23814 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 23808 12396 24593 12424
rect 23808 12384 23814 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 30653 12427 30711 12433
rect 30653 12424 30665 12427
rect 24912 12396 30665 12424
rect 24912 12384 24918 12396
rect 30653 12393 30665 12396
rect 30699 12393 30711 12427
rect 30653 12387 30711 12393
rect 20346 12356 20352 12368
rect 19996 12328 20352 12356
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 19334 12288 19340 12300
rect 18739 12260 19340 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 19996 12232 20024 12328
rect 20346 12316 20352 12328
rect 20404 12316 20410 12368
rect 33962 12356 33968 12368
rect 22388 12328 33968 12356
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 22388 12297 22416 12328
rect 33962 12316 33968 12328
rect 34020 12316 34026 12368
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20128 12260 20913 12288
rect 20128 12248 20134 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 22373 12291 22431 12297
rect 22373 12257 22385 12291
rect 22419 12257 22431 12291
rect 22373 12251 22431 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 22603 12260 23581 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 23569 12257 23581 12260
rect 23615 12257 23627 12291
rect 23569 12251 23627 12257
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 18156 12192 18245 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 19978 12220 19984 12232
rect 19751 12192 19984 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12220 20407 12223
rect 20622 12220 20628 12232
rect 20395 12192 20628 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 22646 12180 22652 12232
rect 22704 12220 22710 12232
rect 23198 12220 23204 12232
rect 22704 12192 23204 12220
rect 22704 12180 22710 12192
rect 23198 12180 23204 12192
rect 23256 12220 23262 12232
rect 23477 12223 23535 12229
rect 23477 12220 23489 12223
rect 23256 12192 23489 12220
rect 23256 12180 23262 12192
rect 23477 12189 23489 12192
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 25406 12220 25412 12232
rect 24811 12192 25268 12220
rect 25367 12192 25412 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 11146 12152 11152 12164
rect 10245 12124 11152 12152
rect 11146 12112 11152 12124
rect 11204 12112 11210 12164
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13081 12155 13139 12161
rect 13081 12152 13093 12155
rect 12952 12124 13093 12152
rect 12952 12112 12958 12124
rect 13081 12121 13093 12124
rect 13127 12121 13139 12155
rect 13081 12115 13139 12121
rect 13182 12155 13240 12161
rect 13182 12121 13194 12155
rect 13228 12152 13240 12155
rect 14369 12155 14427 12161
rect 13228 12124 13308 12152
rect 13228 12121 13240 12124
rect 13182 12115 13240 12121
rect 4080 12056 6408 12084
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 11606 12084 11612 12096
rect 9447 12056 11612 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12986 12084 12992 12096
rect 12391 12056 12992 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13280 12084 13308 12124
rect 14369 12121 14381 12155
rect 14415 12121 14427 12155
rect 14369 12115 14427 12121
rect 14461 12155 14519 12161
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 14550 12152 14556 12164
rect 14507 12124 14556 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 13814 12084 13820 12096
rect 13280 12056 13820 12084
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 14384 12084 14412 12115
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 15010 12152 15016 12164
rect 14971 12124 15016 12152
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 16482 12112 16488 12164
rect 16540 12152 16546 12164
rect 20898 12152 20904 12164
rect 16540 12124 20904 12152
rect 16540 12112 16546 12124
rect 20898 12112 20904 12124
rect 20956 12112 20962 12164
rect 20990 12112 20996 12164
rect 21048 12152 21054 12164
rect 21542 12152 21548 12164
rect 21048 12124 21093 12152
rect 21503 12124 21548 12152
rect 21048 12112 21054 12124
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 19242 12084 19248 12096
rect 14384 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 25240 12093 25268 12192
rect 25406 12180 25412 12192
rect 25464 12180 25470 12232
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12220 30619 12223
rect 38102 12220 38108 12232
rect 30607 12192 38108 12220
rect 30607 12189 30619 12192
rect 30561 12183 30619 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 19521 12087 19579 12093
rect 19521 12084 19533 12087
rect 19484 12056 19533 12084
rect 19484 12044 19490 12056
rect 19521 12053 19533 12056
rect 19567 12053 19579 12087
rect 19521 12047 19579 12053
rect 25225 12087 25283 12093
rect 25225 12053 25237 12087
rect 25271 12053 25283 12087
rect 25225 12047 25283 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 3510 11880 3516 11892
rect 2884 11852 3516 11880
rect 2884 11821 2912 11852
rect 3510 11840 3516 11852
rect 3568 11880 3574 11892
rect 7006 11880 7012 11892
rect 3568 11852 7012 11880
rect 3568 11840 3574 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7193 11883 7251 11889
rect 7193 11849 7205 11883
rect 7239 11880 7251 11883
rect 9306 11880 9312 11892
rect 7239 11852 9312 11880
rect 7239 11849 7251 11852
rect 7193 11843 7251 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 10318 11880 10324 11892
rect 9548 11852 10324 11880
rect 9548 11840 9554 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 10597 11883 10655 11889
rect 10597 11849 10609 11883
rect 10643 11880 10655 11883
rect 11422 11880 11428 11892
rect 10643 11852 11428 11880
rect 10643 11849 10655 11852
rect 10597 11843 10655 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 12345 11883 12403 11889
rect 12345 11849 12357 11883
rect 12391 11880 12403 11883
rect 13357 11883 13415 11889
rect 12391 11852 13308 11880
rect 12391 11849 12403 11852
rect 12345 11843 12403 11849
rect 2869 11815 2927 11821
rect 2869 11781 2881 11815
rect 2915 11781 2927 11815
rect 4614 11812 4620 11824
rect 4575 11784 4620 11812
rect 2869 11775 2927 11781
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 7926 11812 7932 11824
rect 7760 11784 7932 11812
rect 1486 11704 1492 11756
rect 1544 11744 1550 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1544 11716 1685 11744
rect 1544 11704 1550 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 5997 11731 6055 11737
rect 5997 11697 6009 11731
rect 6043 11697 6055 11731
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 7064 11716 7113 11744
rect 7064 11704 7070 11716
rect 7101 11713 7113 11716
rect 7147 11744 7159 11747
rect 7760 11744 7788 11784
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 9030 11772 9036 11824
rect 9088 11772 9094 11824
rect 9398 11772 9404 11824
rect 9456 11812 9462 11824
rect 12434 11812 12440 11824
rect 9456 11784 12440 11812
rect 9456 11772 9462 11784
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 13280 11812 13308 11852
rect 13357 11849 13369 11883
rect 13403 11880 13415 11883
rect 14090 11880 14096 11892
rect 13403 11852 14096 11880
rect 13403 11849 13415 11852
rect 13357 11843 13415 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14918 11880 14924 11892
rect 14200 11852 14924 11880
rect 14200 11812 14228 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 15286 11880 15292 11892
rect 15247 11852 15292 11880
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 16114 11880 16120 11892
rect 16075 11852 16120 11880
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 16850 11880 16856 11892
rect 16811 11852 16856 11880
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 18414 11840 18420 11892
rect 18472 11880 18478 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 18472 11852 19073 11880
rect 18472 11840 18478 11852
rect 19061 11849 19073 11852
rect 19107 11849 19119 11883
rect 19061 11843 19119 11849
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19613 11883 19671 11889
rect 19613 11880 19625 11883
rect 19392 11852 19625 11880
rect 19392 11840 19398 11852
rect 19613 11849 19625 11852
rect 19659 11849 19671 11883
rect 19613 11843 19671 11849
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20622 11880 20628 11892
rect 20487 11852 20628 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 22005 11883 22063 11889
rect 22005 11880 22017 11883
rect 21048 11852 22017 11880
rect 21048 11840 21054 11852
rect 22005 11849 22017 11852
rect 22051 11849 22063 11883
rect 22005 11843 22063 11849
rect 13280 11784 14228 11812
rect 14645 11815 14703 11821
rect 14645 11781 14657 11815
rect 14691 11812 14703 11815
rect 15378 11812 15384 11824
rect 14691 11784 15384 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 19978 11812 19984 11824
rect 15528 11784 19984 11812
rect 15528 11772 15534 11784
rect 7147 11716 7788 11744
rect 9953 11747 10011 11753
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10686 11744 10692 11756
rect 9999 11716 10692 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 12584 11716 13277 11744
rect 12584 11704 12590 11716
rect 13265 11713 13277 11716
rect 13311 11713 13323 11747
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13265 11707 13323 11713
rect 13740 11716 14105 11744
rect 5997 11691 6055 11697
rect 1854 11676 1860 11688
rect 1815 11648 1860 11676
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11645 2651 11679
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 2593 11639 2651 11645
rect 1670 11568 1676 11620
rect 1728 11608 1734 11620
rect 2608 11608 2636 11639
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 1728 11580 2636 11608
rect 1728 11568 1734 11580
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5626 11540 5632 11552
rect 5224 11512 5632 11540
rect 5224 11500 5230 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 5810 11540 5816 11552
rect 5771 11512 5816 11540
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 6012 11540 6040 11691
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 6788 11648 7757 11676
rect 6788 11636 6794 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8662 11676 8668 11688
rect 8067 11648 8668 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 10042 11676 10048 11688
rect 9508 11648 10048 11676
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 9508 11617 9536 11648
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10410 11676 10416 11688
rect 10183 11648 10416 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11388 11648 11713 11676
rect 11388 11636 11394 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11676 11943 11679
rect 12894 11676 12900 11688
rect 11931 11648 12900 11676
rect 11931 11645 11943 11648
rect 11885 11639 11943 11645
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 9493 11611 9551 11617
rect 9493 11608 9505 11611
rect 9272 11580 9505 11608
rect 9272 11568 9278 11580
rect 9493 11577 9505 11580
rect 9539 11577 9551 11611
rect 10226 11608 10232 11620
rect 9493 11571 9551 11577
rect 9876 11580 10232 11608
rect 9876 11540 9904 11580
rect 10226 11568 10232 11580
rect 10284 11568 10290 11620
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 13740 11608 13768 11716
rect 14093 11713 14105 11716
rect 14139 11744 14151 11747
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 14139 11716 14565 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14553 11713 14565 11716
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 15102 11704 15108 11756
rect 15160 11744 15166 11756
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 15160 11716 15209 11744
rect 15160 11704 15166 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16347 11716 17540 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 10376 11580 13768 11608
rect 13832 11580 15608 11608
rect 10376 11568 10382 11580
rect 6012 11512 9904 11540
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 13832 11540 13860 11580
rect 10100 11512 13860 11540
rect 13909 11543 13967 11549
rect 10100 11500 10106 11512
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14642 11540 14648 11552
rect 13955 11512 14648 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15580 11540 15608 11580
rect 15654 11568 15660 11620
rect 15712 11608 15718 11620
rect 17310 11608 17316 11620
rect 15712 11580 17316 11608
rect 15712 11568 15718 11580
rect 17310 11568 17316 11580
rect 17368 11568 17374 11620
rect 17512 11617 17540 11716
rect 17586 11704 17592 11756
rect 17644 11744 17650 11756
rect 18984 11753 19012 11784
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 20714 11772 20720 11824
rect 20772 11812 20778 11824
rect 21177 11815 21235 11821
rect 21177 11812 21189 11815
rect 20772 11784 21189 11812
rect 20772 11772 20778 11784
rect 21177 11781 21189 11784
rect 21223 11781 21235 11815
rect 21177 11775 21235 11781
rect 22112 11784 22876 11812
rect 17681 11747 17739 11753
rect 17681 11744 17693 11747
rect 17644 11716 17693 11744
rect 17644 11704 17650 11716
rect 17681 11713 17693 11716
rect 17727 11713 17739 11747
rect 17681 11707 17739 11713
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 19426 11704 19432 11756
rect 19484 11744 19490 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19484 11716 19809 11744
rect 19484 11704 19490 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 20622 11744 20628 11756
rect 20583 11716 20628 11744
rect 19797 11707 19855 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20956 11716 21097 11744
rect 20956 11704 20962 11716
rect 21085 11713 21097 11716
rect 21131 11744 21143 11747
rect 22112 11744 22140 11784
rect 22848 11753 22876 11784
rect 21131 11716 22140 11744
rect 22189 11747 22247 11753
rect 21131 11713 21143 11716
rect 21085 11707 21143 11713
rect 22189 11713 22201 11747
rect 22235 11744 22247 11747
rect 22833 11747 22891 11753
rect 22235 11716 22692 11744
rect 22235 11713 22247 11716
rect 22189 11707 22247 11713
rect 18138 11636 18144 11688
rect 18196 11676 18202 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 18196 11648 18245 11676
rect 18196 11636 18202 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 20990 11676 20996 11688
rect 19300 11648 20996 11676
rect 19300 11636 19306 11648
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 22664 11617 22692 11716
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 17497 11611 17555 11617
rect 17497 11577 17509 11611
rect 17543 11577 17555 11611
rect 17497 11571 17555 11577
rect 22649 11611 22707 11617
rect 22649 11577 22661 11611
rect 22695 11577 22707 11611
rect 22649 11571 22707 11577
rect 18782 11540 18788 11552
rect 15580 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11540 18846 11552
rect 20622 11540 20628 11552
rect 18840 11512 20628 11540
rect 18840 11500 18846 11512
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2004 11308 3433 11336
rect 2004 11296 2010 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 7285 11339 7343 11345
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 9398 11336 9404 11348
rect 7331 11308 9404 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 11609 11339 11667 11345
rect 11609 11305 11621 11339
rect 11655 11336 11667 11339
rect 11882 11336 11888 11348
rect 11655 11308 11888 11336
rect 11655 11305 11667 11308
rect 11609 11299 11667 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 12308 11308 12357 11336
rect 12308 11296 12314 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12345 11299 12403 11305
rect 13173 11339 13231 11345
rect 13173 11305 13185 11339
rect 13219 11336 13231 11339
rect 13906 11336 13912 11348
rect 13219 11308 13912 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 16390 11336 16396 11348
rect 15795 11308 16396 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 18506 11336 18512 11348
rect 18467 11308 18512 11336
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 20717 11339 20775 11345
rect 20717 11305 20729 11339
rect 20763 11336 20775 11339
rect 20806 11336 20812 11348
rect 20763 11308 20812 11336
rect 20763 11305 20775 11308
rect 20717 11299 20775 11305
rect 20806 11296 20812 11308
rect 20864 11296 20870 11348
rect 21284 11308 22048 11336
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 7800 11240 8248 11268
rect 7800 11228 7806 11240
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 4672 11172 4905 11200
rect 4672 11160 4678 11172
rect 4893 11169 4905 11172
rect 4939 11200 4951 11203
rect 5534 11200 5540 11212
rect 4939 11172 5540 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 5868 11172 6960 11200
rect 5868 11160 5874 11172
rect 1670 11132 1676 11144
rect 1631 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 3752 11104 4261 11132
rect 3752 11092 3758 11104
rect 4249 11101 4261 11104
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 2038 11064 2044 11076
rect 1995 11036 2044 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 2038 11024 2044 11036
rect 2096 11024 2102 11076
rect 2406 11024 2412 11076
rect 2464 11024 2470 11076
rect 4341 11067 4399 11073
rect 4341 11033 4353 11067
rect 4387 11064 4399 11067
rect 5166 11064 5172 11076
rect 4387 11036 5028 11064
rect 5127 11036 5172 11064
rect 4387 11033 4399 11036
rect 4341 11027 4399 11033
rect 5000 10996 5028 11036
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 6178 11024 6184 11076
rect 6236 11024 6242 11076
rect 6932 11064 6960 11172
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7708 11172 7849 11200
rect 7708 11160 7714 11172
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8220 11200 8248 11240
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 8662 11268 8668 11280
rect 8352 11240 8668 11268
rect 8352 11228 8358 11240
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 9490 11228 9496 11280
rect 9548 11268 9554 11280
rect 10502 11268 10508 11280
rect 9548 11240 10508 11268
rect 9548 11228 9554 11240
rect 10502 11228 10508 11240
rect 10560 11268 10566 11280
rect 12158 11268 12164 11280
rect 10560 11240 12164 11268
rect 10560 11228 10566 11240
rect 12158 11228 12164 11240
rect 12216 11268 12222 11280
rect 12216 11240 12664 11268
rect 12216 11228 12222 11240
rect 9214 11200 9220 11212
rect 8220 11172 9220 11200
rect 8021 11163 8079 11169
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 7156 11104 7205 11132
rect 7156 11092 7162 11104
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 8036 11064 8064 11163
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 12250 11200 12256 11212
rect 9999 11172 12256 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8352 11104 9321 11132
rect 8352 11092 8358 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9490 11132 9496 11144
rect 9451 11104 9496 11132
rect 9309 11095 9367 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9916 11104 10425 11132
rect 9916 11092 9922 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10594 11132 10600 11144
rect 10555 11104 10600 11132
rect 10413 11095 10471 11101
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 10704 11104 11529 11132
rect 8478 11064 8484 11076
rect 6932 11036 8064 11064
rect 8439 11036 8484 11064
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 10704 11064 10732 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 11664 11104 12541 11132
rect 11664 11092 11670 11104
rect 12529 11101 12541 11104
rect 12575 11101 12587 11135
rect 12636 11132 12664 11240
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 15105 11271 15163 11277
rect 13044 11240 14504 11268
rect 13044 11228 13050 11240
rect 14476 11141 14504 11240
rect 15105 11237 15117 11271
rect 15151 11237 15163 11271
rect 21284 11268 21312 11308
rect 15105 11231 15163 11237
rect 16408 11240 21312 11268
rect 15120 11200 15148 11231
rect 16408 11209 16436 11240
rect 21358 11228 21364 11280
rect 21416 11268 21422 11280
rect 22020 11268 22048 11308
rect 22462 11296 22468 11348
rect 22520 11296 22526 11348
rect 37182 11296 37188 11348
rect 37240 11336 37246 11348
rect 38105 11339 38163 11345
rect 38105 11336 38117 11339
rect 37240 11308 38117 11336
rect 37240 11296 37246 11308
rect 38105 11305 38117 11308
rect 38151 11305 38163 11339
rect 38105 11299 38163 11305
rect 22480 11268 22508 11296
rect 21416 11240 21864 11268
rect 22020 11240 22508 11268
rect 21416 11228 21422 11240
rect 16393 11203 16451 11209
rect 15120 11172 15976 11200
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12636 11104 13093 11132
rect 12529 11095 12587 11101
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 15948 11141 15976 11172
rect 16393 11169 16405 11203
rect 16439 11169 16451 11203
rect 18138 11200 18144 11212
rect 18099 11172 18144 11200
rect 16393 11163 16451 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11200 20223 11203
rect 21637 11203 21695 11209
rect 21637 11200 21649 11203
rect 20211 11172 21649 11200
rect 20211 11169 20223 11172
rect 20165 11163 20223 11169
rect 21637 11169 21649 11172
rect 21683 11200 21695 11203
rect 21726 11200 21732 11212
rect 21683 11172 21732 11200
rect 21683 11169 21695 11172
rect 21637 11163 21695 11169
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 21836 11200 21864 11240
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 21836 11172 22477 11200
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 22465 11163 22523 11169
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 14700 11104 15301 11132
rect 14700 11092 14706 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 16574 11132 16580 11144
rect 16535 11104 16580 11132
rect 15933 11095 15991 11101
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 17681 11135 17739 11141
rect 17681 11101 17693 11135
rect 17727 11132 17739 11135
rect 17954 11132 17960 11144
rect 17727 11104 17960 11132
rect 17727 11101 17739 11104
rect 17681 11095 17739 11101
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18322 11132 18328 11144
rect 18283 11104 18328 11132
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11101 20683 11135
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 20625 11095 20683 11101
rect 8628 11036 10732 11064
rect 11057 11067 11115 11073
rect 8628 11024 8634 11036
rect 11057 11033 11069 11067
rect 11103 11064 11115 11067
rect 17037 11067 17095 11073
rect 17037 11064 17049 11067
rect 11103 11036 17049 11064
rect 11103 11033 11115 11036
rect 11057 11027 11115 11033
rect 17037 11033 17049 11036
rect 17083 11064 17095 11067
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 17083 11036 19533 11064
rect 17083 11033 17095 11036
rect 17037 11027 17095 11033
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 19613 11067 19671 11073
rect 19613 11033 19625 11067
rect 19659 11033 19671 11067
rect 19613 11027 19671 11033
rect 5902 10996 5908 11008
rect 5000 10968 5908 10996
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 6546 10956 6552 11008
rect 6604 10996 6610 11008
rect 6641 10999 6699 11005
rect 6641 10996 6653 10999
rect 6604 10968 6653 10996
rect 6604 10956 6610 10968
rect 6641 10965 6653 10968
rect 6687 10965 6699 10999
rect 6641 10959 6699 10965
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 10502 10996 10508 11008
rect 7524 10968 10508 10996
rect 7524 10956 7530 10968
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 14277 10999 14335 11005
rect 14277 10965 14289 10999
rect 14323 10996 14335 10999
rect 15746 10996 15752 11008
rect 14323 10968 15752 10996
rect 14323 10965 14335 10968
rect 14277 10959 14335 10965
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 17494 10996 17500 11008
rect 17455 10968 17500 10996
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 19628 10996 19656 11027
rect 19484 10968 19656 10996
rect 20640 10996 20668 11095
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 21358 11064 21364 11076
rect 21319 11036 21364 11064
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 21450 11024 21456 11076
rect 21508 11064 21514 11076
rect 21508 11036 21553 11064
rect 21508 11024 21514 11036
rect 21726 11024 21732 11076
rect 21784 11064 21790 11076
rect 28350 11064 28356 11076
rect 21784 11036 28356 11064
rect 21784 11024 21790 11036
rect 28350 11024 28356 11036
rect 28408 11024 28414 11076
rect 22738 10996 22744 11008
rect 20640 10968 22744 10996
rect 19484 10956 19490 10968
rect 22738 10956 22744 10968
rect 22796 10956 22802 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 1946 10792 1952 10804
rect 1811 10764 1952 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2774 10792 2780 10804
rect 2455 10764 2780 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 3016 10764 3065 10792
rect 3016 10752 3022 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 4065 10795 4123 10801
rect 3476 10764 3924 10792
rect 3476 10752 3482 10764
rect 3896 10724 3924 10764
rect 4065 10761 4077 10795
rect 4111 10792 4123 10795
rect 4154 10792 4160 10804
rect 4111 10764 4160 10792
rect 4111 10761 4123 10764
rect 4065 10755 4123 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5350 10792 5356 10804
rect 5040 10764 5356 10792
rect 5040 10752 5046 10764
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 7558 10792 7564 10804
rect 7519 10764 7564 10792
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 10410 10792 10416 10804
rect 8496 10764 10416 10792
rect 6917 10727 6975 10733
rect 3896 10696 5212 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2314 10656 2320 10668
rect 1719 10628 2320 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2314 10616 2320 10628
rect 2372 10656 2378 10668
rect 2682 10656 2688 10668
rect 2372 10628 2688 10656
rect 2372 10616 2378 10628
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3142 10656 3148 10668
rect 3007 10628 3148 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 5184 10665 5212 10696
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 8496 10724 8524 10764
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13541 10795 13599 10801
rect 13541 10792 13553 10795
rect 13228 10764 13553 10792
rect 13228 10752 13234 10764
rect 13541 10761 13553 10764
rect 13587 10761 13599 10795
rect 13541 10755 13599 10761
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 14056 10764 14749 10792
rect 14056 10752 14062 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 14737 10755 14795 10761
rect 15194 10752 15200 10804
rect 15252 10792 15258 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 15252 10764 15301 10792
rect 15252 10752 15258 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15930 10792 15936 10804
rect 15891 10764 15936 10792
rect 15289 10755 15347 10761
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 16758 10752 16764 10804
rect 16816 10792 16822 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 16816 10764 16865 10792
rect 16816 10752 16822 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 16853 10755 16911 10761
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19484 10764 19625 10792
rect 19484 10752 19490 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21450 10792 21456 10804
rect 21131 10764 21456 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21542 10752 21548 10804
rect 21600 10792 21606 10804
rect 21600 10764 33824 10792
rect 21600 10752 21606 10764
rect 6963 10696 8524 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 8570 10684 8576 10736
rect 8628 10724 8634 10736
rect 9677 10727 9735 10733
rect 8628 10696 9444 10724
rect 8628 10684 8634 10696
rect 3973 10660 4031 10665
rect 3896 10659 4031 10660
rect 3896 10656 3985 10659
rect 3252 10632 3985 10656
rect 3252 10628 3924 10632
rect 2700 10588 2728 10616
rect 3252 10588 3280 10628
rect 3973 10625 3985 10632
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5994 10656 6000 10668
rect 5955 10628 6000 10656
rect 5169 10619 5227 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 7006 10656 7012 10668
rect 6871 10628 7012 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 7466 10656 7472 10668
rect 7427 10628 7472 10656
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10625 8171 10659
rect 8938 10656 8944 10668
rect 8899 10628 8944 10656
rect 8113 10619 8171 10625
rect 2700 10560 3280 10588
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10588 5319 10591
rect 5307 10560 7052 10588
rect 5307 10557 5319 10560
rect 5261 10551 5319 10557
rect 2314 10480 2320 10532
rect 2372 10520 2378 10532
rect 3418 10520 3424 10532
rect 2372 10492 3424 10520
rect 2372 10480 2378 10492
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 7024 10520 7052 10560
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 8128 10588 8156 10619
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9416 10665 9444 10696
rect 9677 10693 9689 10727
rect 9723 10724 9735 10727
rect 9766 10724 9772 10736
rect 9723 10696 9772 10724
rect 9723 10693 9735 10696
rect 9677 10687 9735 10693
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 9950 10684 9956 10736
rect 10008 10724 10014 10736
rect 12250 10724 12256 10736
rect 10008 10696 10166 10724
rect 12211 10696 12256 10724
rect 10008 10684 10014 10696
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 12345 10727 12403 10733
rect 12345 10693 12357 10727
rect 12391 10724 12403 10727
rect 12986 10724 12992 10736
rect 12391 10696 12992 10724
rect 12391 10693 12403 10696
rect 12345 10687 12403 10693
rect 12986 10684 12992 10696
rect 13044 10684 13050 10736
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 17920 10696 28580 10724
rect 17920 10684 17926 10696
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13320 10628 13461 10656
rect 13320 10616 13326 10628
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 14642 10656 14648 10668
rect 14603 10628 14648 10656
rect 13449 10619 13507 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15620 10628 16129 10656
rect 15620 10616 15626 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17494 10656 17500 10668
rect 17083 10628 17500 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17954 10656 17960 10668
rect 17915 10628 17960 10656
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 19518 10656 19524 10668
rect 18064 10628 19524 10656
rect 7432 10560 8156 10588
rect 8205 10591 8263 10597
rect 7432 10548 7438 10560
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 11698 10588 11704 10600
rect 8251 10560 9260 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 8386 10520 8392 10532
rect 7024 10492 8392 10520
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 9232 10520 9260 10560
rect 9508 10560 11704 10588
rect 9508 10520 9536 10560
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 18064 10588 18092 10628
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 20588 10628 21281 10656
rect 20588 10616 20594 10628
rect 21269 10625 21281 10628
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21634 10616 21640 10668
rect 21692 10656 21698 10668
rect 22741 10659 22799 10665
rect 22741 10656 22753 10659
rect 21692 10628 22753 10656
rect 21692 10616 21698 10628
rect 22741 10625 22753 10628
rect 22787 10625 22799 10659
rect 27154 10656 27160 10668
rect 27115 10628 27160 10656
rect 22741 10619 22799 10625
rect 27154 10616 27160 10628
rect 27212 10616 27218 10668
rect 27246 10616 27252 10668
rect 27304 10656 27310 10668
rect 28552 10665 28580 10696
rect 33796 10665 33824 10764
rect 28537 10659 28595 10665
rect 27304 10628 27349 10656
rect 27304 10616 27310 10628
rect 28537 10625 28549 10659
rect 28583 10625 28595 10659
rect 28537 10619 28595 10625
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10625 33839 10659
rect 33781 10619 33839 10625
rect 18414 10588 18420 10600
rect 12584 10560 18092 10588
rect 18375 10560 18420 10588
rect 12584 10548 12590 10560
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18598 10588 18604 10600
rect 18559 10560 18604 10588
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 9232 10492 9536 10520
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13078 10520 13084 10532
rect 12851 10492 13084 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 18506 10480 18512 10532
rect 18564 10520 18570 10532
rect 18785 10523 18843 10529
rect 18785 10520 18797 10523
rect 18564 10492 18797 10520
rect 18564 10480 18570 10492
rect 18785 10489 18797 10492
rect 18831 10489 18843 10523
rect 18785 10483 18843 10489
rect 28629 10523 28687 10529
rect 28629 10489 28641 10523
rect 28675 10520 28687 10523
rect 34146 10520 34152 10532
rect 28675 10492 34152 10520
rect 28675 10489 28687 10492
rect 28629 10483 28687 10489
rect 34146 10480 34152 10492
rect 34204 10480 34210 10532
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 5813 10455 5871 10461
rect 5813 10452 5825 10455
rect 2648 10424 5825 10452
rect 2648 10412 2654 10424
rect 5813 10421 5825 10424
rect 5859 10421 5871 10455
rect 8754 10452 8760 10464
rect 8715 10424 8760 10452
rect 5813 10415 5871 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 10870 10452 10876 10464
rect 8904 10424 10876 10452
rect 8904 10412 8910 10424
rect 10870 10412 10876 10424
rect 10928 10452 10934 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 10928 10424 11161 10452
rect 10928 10412 10934 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 17773 10455 17831 10461
rect 17773 10421 17785 10455
rect 17819 10452 17831 10455
rect 18690 10452 18696 10464
rect 17819 10424 18696 10452
rect 17819 10421 17831 10424
rect 17773 10415 17831 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 22833 10455 22891 10461
rect 22833 10421 22845 10455
rect 22879 10452 22891 10455
rect 23566 10452 23572 10464
rect 22879 10424 23572 10452
rect 22879 10421 22891 10424
rect 22833 10415 22891 10421
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 33873 10455 33931 10461
rect 33873 10421 33885 10455
rect 33919 10452 33931 10455
rect 36354 10452 36360 10464
rect 33919 10424 36360 10452
rect 33919 10421 33931 10424
rect 33873 10415 33931 10421
rect 36354 10412 36360 10424
rect 36412 10412 36418 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 2041 10251 2099 10257
rect 2041 10248 2053 10251
rect 1360 10220 2053 10248
rect 1360 10208 1366 10220
rect 2041 10217 2053 10220
rect 2087 10217 2099 10251
rect 3326 10248 3332 10260
rect 3287 10220 3332 10248
rect 2041 10211 2099 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3694 10208 3700 10260
rect 3752 10248 3758 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3752 10220 4077 10248
rect 3752 10208 3758 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 4880 10251 4938 10257
rect 4880 10217 4892 10251
rect 4926 10248 4938 10251
rect 6546 10248 6552 10260
rect 4926 10220 6552 10248
rect 4926 10217 4938 10220
rect 4880 10211 4938 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7193 10251 7251 10257
rect 7193 10217 7205 10251
rect 7239 10248 7251 10251
rect 8018 10248 8024 10260
rect 7239 10220 8024 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8389 10251 8447 10257
rect 8389 10248 8401 10251
rect 8168 10220 8401 10248
rect 8168 10208 8174 10220
rect 8389 10217 8401 10220
rect 8435 10217 8447 10251
rect 9950 10248 9956 10260
rect 8389 10211 8447 10217
rect 8496 10220 9956 10248
rect 2685 10183 2743 10189
rect 2685 10149 2697 10183
rect 2731 10180 2743 10183
rect 3786 10180 3792 10192
rect 2731 10152 3792 10180
rect 2731 10149 2743 10152
rect 2685 10143 2743 10149
rect 3786 10140 3792 10152
rect 3844 10140 3850 10192
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 8496 10180 8524 10220
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10778 10208 10784 10260
rect 10836 10248 10842 10260
rect 10836 10220 11652 10248
rect 10836 10208 10842 10220
rect 7524 10152 8524 10180
rect 7524 10140 7530 10152
rect 8570 10140 8576 10192
rect 8628 10140 8634 10192
rect 9122 10140 9128 10192
rect 9180 10180 9186 10192
rect 11517 10183 11575 10189
rect 9180 10152 9352 10180
rect 9180 10140 9186 10152
rect 4614 10112 4620 10124
rect 4575 10084 4620 10112
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6270 10112 6276 10124
rect 5960 10084 6276 10112
rect 5960 10072 5966 10084
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 8588 10112 8616 10140
rect 9217 10115 9275 10121
rect 9217 10112 9229 10115
rect 6972 10084 9229 10112
rect 6972 10072 6978 10084
rect 9217 10081 9229 10084
rect 9263 10081 9275 10115
rect 9324 10112 9352 10152
rect 11517 10149 11529 10183
rect 11563 10149 11575 10183
rect 11624 10180 11652 10220
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 12032 10220 12173 10248
rect 12032 10208 12038 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12768 10220 12817 10248
rect 12768 10208 12774 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 14458 10248 14464 10260
rect 14323 10220 14464 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15562 10248 15568 10260
rect 14752 10220 15056 10248
rect 15523 10220 15568 10248
rect 14642 10180 14648 10192
rect 11624 10152 14648 10180
rect 11517 10143 11575 10149
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9324 10084 9505 10112
rect 9217 10075 9275 10081
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 11532 10112 11560 10143
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 9640 10084 10824 10112
rect 11532 10084 12388 10112
rect 9640 10072 9646 10084
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2593 10047 2651 10053
rect 2593 10044 2605 10047
rect 1995 10016 2605 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2593 10013 2605 10016
rect 2639 10044 2651 10047
rect 2682 10044 2688 10056
rect 2639 10016 2688 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 3142 10004 3148 10056
rect 3200 10044 3206 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 3200 10016 3249 10044
rect 3200 10004 3206 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3973 10047 4031 10053
rect 3973 10044 3985 10047
rect 3660 10016 3985 10044
rect 3660 10004 3666 10016
rect 3973 10013 3985 10016
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7374 10044 7380 10056
rect 7147 10016 7380 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8294 10044 8300 10056
rect 7791 10016 8300 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 4798 9976 4804 9988
rect 4580 9948 4804 9976
rect 4580 9936 4586 9948
rect 4798 9936 4804 9948
rect 4856 9936 4862 9988
rect 5626 9936 5632 9988
rect 5684 9936 5690 9988
rect 6288 9948 9536 9976
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 6288 9908 6316 9948
rect 2096 9880 6316 9908
rect 6365 9911 6423 9917
rect 2096 9868 2102 9880
rect 6365 9877 6377 9911
rect 6411 9908 6423 9911
rect 6730 9908 6736 9920
rect 6411 9880 6736 9908
rect 6411 9877 6423 9880
rect 6365 9871 6423 9877
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 9508 9908 9536 9948
rect 9582 9936 9588 9988
rect 9640 9976 9646 9988
rect 10796 9976 10824 10084
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 12360 10053 12388 10084
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 13541 10115 13599 10121
rect 12768 10084 13492 10112
rect 12768 10072 12774 10084
rect 13464 10053 13492 10084
rect 13541 10081 13553 10115
rect 13587 10112 13599 10115
rect 14752 10112 14780 10220
rect 14921 10183 14979 10189
rect 14921 10149 14933 10183
rect 14967 10149 14979 10183
rect 15028 10180 15056 10220
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 18322 10208 18328 10260
rect 18380 10248 18386 10260
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 18380 10220 18521 10248
rect 18380 10208 18386 10220
rect 18509 10217 18521 10220
rect 18555 10217 18567 10251
rect 18509 10211 18567 10217
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 18656 10220 19533 10248
rect 18656 10208 18662 10220
rect 19521 10217 19533 10220
rect 19567 10217 19579 10251
rect 20530 10248 20536 10260
rect 20491 10220 20536 10248
rect 19521 10211 19579 10217
rect 20530 10208 20536 10220
rect 20588 10208 20594 10260
rect 33962 10248 33968 10260
rect 33923 10220 33968 10248
rect 33962 10208 33968 10220
rect 34020 10208 34026 10260
rect 16206 10180 16212 10192
rect 15028 10152 16212 10180
rect 14921 10143 14979 10149
rect 13587 10084 14780 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 10928 10016 11713 10044
rect 10928 10004 10934 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 14936 10044 14964 10143
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18012 10084 19472 10112
rect 18012 10072 18018 10084
rect 15102 10044 15108 10056
rect 14507 10016 14964 10044
rect 15063 10016 15108 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 9640 9948 9982 9976
rect 10796 9948 11100 9976
rect 9640 9936 9646 9948
rect 10778 9908 10784 9920
rect 9508 9880 10784 9908
rect 10778 9868 10784 9880
rect 10836 9908 10842 9920
rect 10965 9911 11023 9917
rect 10965 9908 10977 9911
rect 10836 9880 10977 9908
rect 10836 9868 10842 9880
rect 10965 9877 10977 9880
rect 11011 9877 11023 9911
rect 11072 9908 11100 9948
rect 11422 9936 11428 9988
rect 11480 9976 11486 9988
rect 12526 9976 12532 9988
rect 11480 9948 12532 9976
rect 11480 9936 11486 9948
rect 12526 9936 12532 9948
rect 12584 9936 12590 9988
rect 13004 9976 13032 10007
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 17218 10044 17224 10056
rect 16807 10016 17224 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 15764 9976 15792 10007
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 18690 10044 18696 10056
rect 18651 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 19444 10053 19472 10084
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 19576 10016 20729 10044
rect 19576 10004 19582 10016
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 28258 10044 28264 10056
rect 28219 10016 28264 10044
rect 20717 10007 20775 10013
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 28350 10004 28356 10056
rect 28408 10044 28414 10056
rect 29733 10047 29791 10053
rect 29733 10044 29745 10047
rect 28408 10016 29745 10044
rect 28408 10004 28414 10016
rect 29733 10013 29745 10016
rect 29779 10013 29791 10047
rect 29733 10007 29791 10013
rect 33873 10047 33931 10053
rect 33873 10013 33885 10047
rect 33919 10044 33931 10047
rect 37182 10044 37188 10056
rect 33919 10016 37188 10044
rect 33919 10013 33931 10016
rect 33873 10007 33931 10013
rect 37182 10004 37188 10016
rect 37240 10004 37246 10056
rect 12728 9948 13032 9976
rect 14476 9948 15792 9976
rect 12728 9908 12756 9948
rect 14476 9920 14504 9948
rect 11072 9880 12756 9908
rect 10965 9871 11023 9877
rect 14458 9868 14464 9920
rect 14516 9868 14522 9920
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 18506 9908 18512 9920
rect 16899 9880 18512 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 28353 9911 28411 9917
rect 28353 9877 28365 9911
rect 28399 9908 28411 9911
rect 29638 9908 29644 9920
rect 28399 9880 29644 9908
rect 28399 9877 28411 9880
rect 28353 9871 28411 9877
rect 29638 9868 29644 9880
rect 29696 9868 29702 9920
rect 29825 9911 29883 9917
rect 29825 9877 29837 9911
rect 29871 9908 29883 9911
rect 31662 9908 31668 9920
rect 29871 9880 31668 9908
rect 29871 9877 29883 9880
rect 29825 9871 29883 9877
rect 31662 9868 31668 9880
rect 31720 9868 31726 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 2648 9676 4660 9704
rect 2648 9664 2654 9676
rect 1210 9596 1216 9648
rect 1268 9636 1274 9648
rect 1857 9639 1915 9645
rect 1857 9636 1869 9639
rect 1268 9608 1869 9636
rect 1268 9596 1274 9608
rect 1857 9605 1869 9608
rect 1903 9605 1915 9639
rect 2498 9636 2504 9648
rect 2459 9608 2504 9636
rect 1857 9599 1915 9605
rect 2498 9596 2504 9608
rect 2556 9596 2562 9648
rect 3602 9636 3608 9648
rect 2700 9608 3608 9636
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 1780 9500 1808 9531
rect 1946 9528 1952 9580
rect 2004 9568 2010 9580
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2004 9540 2421 9568
rect 2004 9528 2010 9540
rect 2409 9537 2421 9540
rect 2455 9568 2467 9571
rect 2590 9568 2596 9580
rect 2455 9540 2596 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 2700 9500 2728 9608
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 4632 9568 4660 9676
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 5442 9704 5448 9716
rect 4856 9676 5448 9704
rect 4856 9664 4862 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5534 9664 5540 9716
rect 5592 9664 5598 9716
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 8110 9704 8116 9716
rect 7064 9676 8116 9704
rect 7064 9664 7070 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 8938 9704 8944 9716
rect 8352 9676 8944 9704
rect 8352 9664 8358 9676
rect 8938 9664 8944 9676
rect 8996 9704 9002 9716
rect 8996 9676 11192 9704
rect 8996 9664 9002 9676
rect 5552 9636 5580 9664
rect 6914 9636 6920 9648
rect 5552 9608 6920 9636
rect 5258 9568 5264 9580
rect 1780 9472 2728 9500
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 3694 9500 3700 9512
rect 3375 9472 3700 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 2590 9364 2596 9376
rect 1636 9336 2596 9364
rect 1636 9324 1642 9336
rect 2590 9324 2596 9336
rect 2648 9364 2654 9376
rect 3068 9364 3096 9463
rect 3694 9460 3700 9472
rect 3752 9460 3758 9512
rect 4448 9432 4476 9554
rect 4632 9540 5264 9568
rect 5258 9528 5264 9540
rect 5316 9568 5322 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5316 9540 5549 9568
rect 5316 9528 5322 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 6086 9568 6092 9580
rect 5675 9540 6092 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 6086 9528 6092 9540
rect 6144 9528 6150 9580
rect 6564 9577 6592 9608
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 8386 9636 8392 9648
rect 8050 9608 8392 9636
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 11054 9636 11060 9648
rect 8812 9608 10548 9636
rect 11015 9608 11060 9636
rect 8812 9596 8818 9608
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9537 6607 9571
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 6549 9531 6607 9537
rect 8312 9540 9229 9568
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5442 9500 5448 9512
rect 5123 9472 5448 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5442 9460 5448 9472
rect 5500 9500 5506 9512
rect 5500 9472 6684 9500
rect 5500 9460 5506 9472
rect 5166 9432 5172 9444
rect 4448 9404 5172 9432
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 2648 9336 3096 9364
rect 2648 9324 2654 9336
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 5810 9364 5816 9376
rect 3844 9336 5816 9364
rect 3844 9324 3850 9336
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6656 9364 6684 9472
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7558 9500 7564 9512
rect 6880 9472 7564 9500
rect 6880 9460 6886 9472
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7926 9392 7932 9444
rect 7984 9432 7990 9444
rect 8312 9441 8340 9540
rect 9217 9537 9229 9540
rect 9263 9568 9275 9571
rect 9398 9568 9404 9580
rect 9263 9540 9404 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10134 9568 10140 9580
rect 9907 9540 10140 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10520 9577 10548 9608
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 10505 9571 10563 9577
rect 10505 9537 10517 9571
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10928 9540 10977 9568
rect 10928 9528 10934 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 11164 9568 11192 9676
rect 12250 9596 12256 9648
rect 12308 9636 12314 9648
rect 12529 9639 12587 9645
rect 12529 9636 12541 9639
rect 12308 9608 12541 9636
rect 12308 9596 12314 9608
rect 12529 9605 12541 9608
rect 12575 9605 12587 9639
rect 12529 9599 12587 9605
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 13081 9639 13139 9645
rect 13081 9636 13093 9639
rect 12860 9608 13093 9636
rect 12860 9596 12866 9608
rect 13081 9605 13093 9608
rect 13127 9605 13139 9639
rect 14550 9636 14556 9648
rect 14511 9608 14556 9636
rect 13081 9599 13139 9605
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 12069 9571 12127 9577
rect 11164 9540 12020 9568
rect 10965 9531 11023 9537
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 10152 9500 10180 9528
rect 10778 9500 10784 9512
rect 8812 9472 9812 9500
rect 10152 9472 10784 9500
rect 8812 9460 8818 9472
rect 8297 9435 8355 9441
rect 8297 9432 8309 9435
rect 7984 9404 8309 9432
rect 7984 9392 7990 9404
rect 8297 9401 8309 9404
rect 8343 9401 8355 9435
rect 8297 9395 8355 9401
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 8628 9404 9689 9432
rect 8628 9392 8634 9404
rect 9677 9401 9689 9404
rect 9723 9401 9735 9435
rect 9677 9395 9735 9401
rect 8754 9364 8760 9376
rect 6656 9336 8760 9364
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9784 9364 9812 9472
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 11882 9500 11888 9512
rect 11843 9472 11888 9500
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 11992 9500 12020 9540
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12434 9568 12440 9580
rect 12115 9540 12440 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 13998 9568 14004 9580
rect 13959 9540 14004 9568
rect 12989 9531 13047 9537
rect 13004 9500 13032 9531
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 14458 9568 14464 9580
rect 14419 9540 14464 9568
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 11992 9472 13032 9500
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 15304 9500 15332 9531
rect 31662 9528 31668 9580
rect 31720 9568 31726 9580
rect 34517 9571 34575 9577
rect 34517 9568 34529 9571
rect 31720 9540 34529 9568
rect 31720 9528 31726 9540
rect 34517 9537 34529 9540
rect 34563 9537 34575 9571
rect 34517 9531 34575 9537
rect 25222 9500 25228 9512
rect 14148 9472 15332 9500
rect 22066 9472 25228 9500
rect 14148 9460 14154 9472
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9432 10379 9435
rect 12066 9432 12072 9444
rect 10367 9404 12072 9432
rect 10367 9401 10379 9404
rect 10321 9395 10379 9401
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 22066 9432 22094 9472
rect 25222 9460 25228 9472
rect 25280 9460 25286 9512
rect 12406 9404 22094 9432
rect 12406 9364 12434 9404
rect 13814 9364 13820 9376
rect 9784 9336 12434 9364
rect 13775 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 15105 9367 15163 9373
rect 15105 9333 15117 9367
rect 15151 9364 15163 9367
rect 16574 9364 16580 9376
rect 15151 9336 16580 9364
rect 15151 9333 15163 9336
rect 15105 9327 15163 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 34333 9367 34391 9373
rect 34333 9333 34345 9367
rect 34379 9364 34391 9367
rect 38010 9364 38016 9376
rect 34379 9336 38016 9364
rect 34379 9333 34391 9336
rect 34333 9327 34391 9333
rect 38010 9324 38016 9336
rect 38068 9324 38074 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 7098 9169 7104 9172
rect 7088 9163 7104 9169
rect 3476 9132 6500 9160
rect 3476 9120 3482 9132
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9092 3387 9095
rect 3510 9092 3516 9104
rect 3375 9064 3516 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2222 9024 2228 9036
rect 1903 8996 2228 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 2648 8996 4353 9024
rect 2648 8984 2654 8996
rect 4341 8993 4353 8996
rect 4387 9024 4399 9027
rect 4614 9024 4620 9036
rect 4387 8996 4620 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2498 8848 2504 8900
rect 2556 8848 2562 8900
rect 4617 8891 4675 8897
rect 4617 8857 4629 8891
rect 4663 8857 4675 8891
rect 4617 8851 4675 8857
rect 4632 8820 4660 8851
rect 5626 8848 5632 8900
rect 5684 8848 5690 8900
rect 6362 8888 6368 8900
rect 6323 8860 6368 8888
rect 6362 8848 6368 8860
rect 6420 8848 6426 8900
rect 6472 8888 6500 9132
rect 7088 9129 7100 9163
rect 7088 9123 7104 9129
rect 7098 9120 7104 9123
rect 7156 9120 7162 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8168 9132 8708 9160
rect 8168 9120 8174 9132
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 8573 9095 8631 9101
rect 8573 9092 8585 9095
rect 8352 9064 8585 9092
rect 8352 9052 8358 9064
rect 8573 9061 8585 9064
rect 8619 9061 8631 9095
rect 8680 9092 8708 9132
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9548 9132 9689 9160
rect 9548 9120 9554 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 9824 9132 12081 9160
rect 9824 9120 9830 9132
rect 12069 9129 12081 9132
rect 12115 9160 12127 9163
rect 12618 9160 12624 9172
rect 12115 9132 12434 9160
rect 12579 9132 12624 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 10134 9092 10140 9104
rect 8680 9064 10140 9092
rect 8573 9055 8631 9061
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 12406 9092 12434 9132
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 13998 9120 14004 9172
rect 14056 9160 14062 9172
rect 14921 9163 14979 9169
rect 14921 9160 14933 9163
rect 14056 9132 14933 9160
rect 14056 9120 14062 9132
rect 14921 9129 14933 9132
rect 14967 9129 14979 9163
rect 14921 9123 14979 9129
rect 20254 9120 20260 9172
rect 20312 9160 20318 9172
rect 25225 9163 25283 9169
rect 25225 9160 25237 9163
rect 20312 9132 25237 9160
rect 20312 9120 20318 9132
rect 25225 9129 25237 9132
rect 25271 9129 25283 9163
rect 25225 9123 25283 9129
rect 13262 9092 13268 9104
rect 12406 9064 13268 9092
rect 13262 9052 13268 9064
rect 13320 9052 13326 9104
rect 14182 9052 14188 9104
rect 14240 9092 14246 9104
rect 14369 9095 14427 9101
rect 14369 9092 14381 9095
rect 14240 9064 14381 9092
rect 14240 9052 14246 9064
rect 14369 9061 14381 9064
rect 14415 9061 14427 9095
rect 14369 9055 14427 9061
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 7616 8996 8432 9024
rect 7616 8984 7622 8996
rect 8404 8888 8432 8996
rect 8938 8984 8944 9036
rect 8996 9024 9002 9036
rect 10597 9027 10655 9033
rect 8996 8996 10180 9024
rect 8996 8984 9002 8996
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9088 8928 9873 8956
rect 9088 8916 9094 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10152 8888 10180 8996
rect 10597 8993 10609 9027
rect 10643 9024 10655 9027
rect 10962 9024 10968 9036
rect 10643 8996 10968 9024
rect 10643 8993 10655 8996
rect 10597 8987 10655 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 17954 9024 17960 9036
rect 11112 8996 17960 9024
rect 11112 8984 11118 8996
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 12406 8956 12434 8996
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12406 8928 12541 8956
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13170 8956 13176 8968
rect 12860 8928 13176 8956
rect 12860 8916 12866 8928
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 13354 8956 13360 8968
rect 13315 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 15105 8959 15163 8965
rect 15105 8956 15117 8959
rect 14323 8928 15117 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 15105 8925 15117 8928
rect 15151 8925 15163 8959
rect 15105 8919 15163 8925
rect 25133 8959 25191 8965
rect 25133 8925 25145 8959
rect 25179 8956 25191 8959
rect 28626 8956 28632 8968
rect 25179 8928 28632 8956
rect 25179 8925 25191 8928
rect 25133 8919 25191 8925
rect 10870 8888 10876 8900
rect 6472 8860 7590 8888
rect 8404 8860 9674 8888
rect 10152 8860 10876 8888
rect 6822 8820 6828 8832
rect 4632 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 7006 8780 7012 8832
rect 7064 8820 7070 8832
rect 8478 8820 8484 8832
rect 7064 8792 8484 8820
rect 7064 8780 7070 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 9646 8820 9674 8860
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 11238 8848 11244 8900
rect 11296 8848 11302 8900
rect 14292 8888 14320 8919
rect 28626 8916 28632 8928
rect 28684 8916 28690 8968
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 12406 8860 14320 8888
rect 12406 8820 12434 8860
rect 9646 8792 12434 8820
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 12584 8792 13185 8820
rect 12584 8780 12590 8792
rect 13173 8789 13185 8792
rect 13219 8789 13231 8823
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 13173 8783 13231 8789
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 4617 8619 4675 8625
rect 2516 8588 4568 8616
rect 2516 8557 2544 8588
rect 2501 8551 2559 8557
rect 2501 8517 2513 8551
rect 2547 8517 2559 8551
rect 4540 8548 4568 8588
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 4890 8616 4896 8628
rect 4663 8588 4896 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 5132 8588 5273 8616
rect 5132 8576 5138 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5776 8588 5917 8616
rect 5776 8576 5782 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 6420 8588 9260 8616
rect 6420 8576 6426 8588
rect 6380 8548 6408 8576
rect 8018 8548 8024 8560
rect 4540 8520 6408 8548
rect 6564 8520 8024 8548
rect 2501 8511 2559 8517
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 1854 8480 1860 8492
rect 1627 8452 1860 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1854 8440 1860 8452
rect 1912 8480 1918 8492
rect 2038 8480 2044 8492
rect 1912 8452 2044 8480
rect 1912 8440 1918 8452
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 3844 8452 4537 8480
rect 3844 8440 3850 8452
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 5132 8452 5181 8480
rect 5132 8440 5138 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5169 8443 5227 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8381 2283 8415
rect 2225 8375 2283 8381
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 2240 8344 2268 8375
rect 3694 8372 3700 8424
rect 3752 8412 3758 8424
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3752 8384 3985 8412
rect 3752 8372 3758 8384
rect 3973 8381 3985 8384
rect 4019 8412 4031 8415
rect 6564 8412 6592 8520
rect 8018 8508 8024 8520
rect 8076 8508 8082 8560
rect 8478 8508 8484 8560
rect 8536 8508 8542 8560
rect 9232 8548 9260 8588
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 9364 8588 9413 8616
rect 9364 8576 9370 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 10284 8588 10333 8616
rect 10284 8576 10290 8588
rect 10321 8585 10333 8588
rect 10367 8585 10379 8619
rect 10321 8579 10379 8585
rect 11057 8619 11115 8625
rect 11057 8585 11069 8619
rect 11103 8616 11115 8619
rect 11146 8616 11152 8628
rect 11103 8588 11152 8616
rect 11103 8585 11115 8588
rect 11057 8579 11115 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11572 8588 11805 8616
rect 11572 8576 11578 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 12342 8616 12348 8628
rect 12303 8588 12348 8616
rect 11793 8579 11851 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12986 8616 12992 8628
rect 12947 8588 12992 8616
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14090 8616 14096 8628
rect 14047 8588 14096 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 14734 8616 14740 8628
rect 14695 8588 14740 8616
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 14826 8576 14832 8628
rect 14884 8616 14890 8628
rect 25406 8616 25412 8628
rect 14884 8588 25412 8616
rect 14884 8576 14890 8588
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 17310 8548 17316 8560
rect 9232 8520 17316 8548
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 17494 8508 17500 8560
rect 17552 8548 17558 8560
rect 22554 8548 22560 8560
rect 17552 8520 22560 8548
rect 17552 8508 17558 8520
rect 22554 8508 22560 8520
rect 22612 8508 22618 8560
rect 7006 8480 7012 8492
rect 6967 8452 7012 8480
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 10502 8480 10508 8492
rect 10463 8452 10508 8480
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 10962 8480 10968 8492
rect 10836 8452 10968 8480
rect 10836 8440 10842 8452
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11698 8480 11704 8492
rect 11659 8452 11704 8480
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 13170 8480 13176 8492
rect 13131 8452 13176 8480
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13320 8452 14197 8480
rect 13320 8440 13326 8452
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14642 8480 14648 8492
rect 14603 8452 14648 8480
rect 14185 8443 14243 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8480 21235 8483
rect 22002 8480 22008 8492
rect 21223 8452 22008 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 4019 8384 5212 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 1636 8316 2268 8344
rect 1636 8304 1642 8316
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 2682 8276 2688 8288
rect 2372 8248 2688 8276
rect 2372 8236 2378 8248
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 5184 8276 5212 8384
rect 5368 8384 6592 8412
rect 5368 8276 5396 8384
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 6972 8384 7665 8412
rect 6972 8372 6978 8384
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7653 8375 7711 8381
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 14826 8412 14832 8424
rect 8076 8384 14832 8412
rect 8076 8372 8082 8384
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 7098 8344 7104 8356
rect 7059 8316 7104 8344
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 11698 8344 11704 8356
rect 9364 8316 11704 8344
rect 9364 8304 9370 8316
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 13354 8344 13360 8356
rect 11808 8316 13360 8344
rect 5184 8248 5396 8276
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 8478 8276 8484 8288
rect 8168 8248 8484 8276
rect 8168 8236 8174 8248
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 11808 8276 11836 8316
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 17034 8304 17040 8356
rect 17092 8344 17098 8356
rect 20180 8344 20208 8443
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 33962 8480 33968 8492
rect 33923 8452 33968 8480
rect 33962 8440 33968 8452
rect 34020 8440 34026 8492
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 22462 8412 22468 8424
rect 21315 8384 22468 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 17092 8316 20208 8344
rect 20257 8347 20315 8353
rect 17092 8304 17098 8316
rect 20257 8313 20269 8347
rect 20303 8344 20315 8347
rect 21174 8344 21180 8356
rect 20303 8316 21180 8344
rect 20303 8313 20315 8316
rect 20257 8307 20315 8313
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 22370 8304 22376 8356
rect 22428 8344 22434 8356
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 22428 8316 34069 8344
rect 22428 8304 22434 8316
rect 34057 8313 34069 8316
rect 34103 8313 34115 8347
rect 34057 8307 34115 8313
rect 10192 8248 11836 8276
rect 10192 8236 10198 8248
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 4798 8072 4804 8084
rect 4755 8044 4804 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 7926 8072 7932 8084
rect 5776 8044 7512 8072
rect 7887 8044 7932 8072
rect 5776 8032 5782 8044
rect 3326 8004 3332 8016
rect 3287 7976 3332 8004
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 4982 8004 4988 8016
rect 4111 7976 4988 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 7484 8004 7512 8044
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 10594 8072 10600 8084
rect 9815 8044 10600 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12894 8072 12900 8084
rect 12759 8044 12900 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13228 8044 13277 8072
rect 13228 8032 13234 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 27982 8072 27988 8084
rect 27943 8044 27988 8072
rect 13265 8035 13323 8041
rect 27982 8032 27988 8044
rect 28040 8032 28046 8084
rect 37182 8032 37188 8084
rect 37240 8072 37246 8084
rect 38105 8075 38163 8081
rect 38105 8072 38117 8075
rect 37240 8044 38117 8072
rect 37240 8032 37246 8044
rect 38105 8041 38117 8044
rect 38151 8041 38163 8075
rect 38105 8035 38163 8041
rect 10042 8004 10048 8016
rect 7484 7976 10048 8004
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 11698 7964 11704 8016
rect 11756 8004 11762 8016
rect 11756 7976 12434 8004
rect 11756 7964 11762 7976
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 6181 7939 6239 7945
rect 3200 7908 4660 7936
rect 3200 7896 3206 7908
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 4632 7877 4660 7908
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 6914 7936 6920 7948
rect 6227 7908 6920 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 11790 7936 11796 7948
rect 10652 7908 11796 7936
rect 10652 7896 10658 7908
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 12406 7936 12434 7976
rect 12406 7908 13492 7936
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3752 7840 3985 7868
rect 3752 7828 3758 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 4617 7831 4675 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 9674 7868 9680 7880
rect 9635 7840 9680 7868
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 13464 7877 13492 7908
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 12406 7840 12633 7868
rect 1857 7803 1915 7809
rect 1857 7769 1869 7803
rect 1903 7769 1915 7803
rect 1857 7763 1915 7769
rect 1872 7732 1900 7763
rect 2866 7760 2872 7812
rect 2924 7760 2930 7812
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 5353 7803 5411 7809
rect 5353 7800 5365 7803
rect 4120 7772 5365 7800
rect 4120 7760 4126 7772
rect 5353 7769 5365 7772
rect 5399 7769 5411 7803
rect 5353 7763 5411 7769
rect 6457 7803 6515 7809
rect 6457 7769 6469 7803
rect 6503 7769 6515 7803
rect 6457 7763 6515 7769
rect 5442 7732 5448 7744
rect 1872 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6472 7732 6500 7763
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 6604 7772 6946 7800
rect 6604 7760 6610 7772
rect 10502 7760 10508 7812
rect 10560 7800 10566 7812
rect 10597 7803 10655 7809
rect 10597 7800 10609 7803
rect 10560 7772 10609 7800
rect 10560 7760 10566 7772
rect 10597 7769 10609 7772
rect 10643 7769 10655 7803
rect 10597 7763 10655 7769
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 10928 7772 11086 7800
rect 10928 7760 10934 7772
rect 8294 7732 8300 7744
rect 6472 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 9950 7692 9956 7744
rect 10008 7732 10014 7744
rect 12069 7735 12127 7741
rect 12069 7732 12081 7735
rect 10008 7704 12081 7732
rect 10008 7692 10014 7704
rect 12069 7701 12081 7704
rect 12115 7732 12127 7735
rect 12406 7732 12434 7840
rect 12621 7837 12633 7840
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7868 27951 7871
rect 33594 7868 33600 7880
rect 27939 7840 33600 7868
rect 27939 7837 27951 7840
rect 27893 7831 27951 7837
rect 12636 7800 12664 7831
rect 33594 7828 33600 7840
rect 33652 7828 33658 7880
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 15102 7800 15108 7812
rect 12636 7772 15108 7800
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 12115 7704 12434 7732
rect 12115 7701 12127 7704
rect 12069 7695 12127 7701
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 3421 7531 3479 7537
rect 3421 7497 3433 7531
rect 3467 7528 3479 7531
rect 4706 7528 4712 7540
rect 3467 7500 4712 7528
rect 3467 7497 3479 7500
rect 3421 7491 3479 7497
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5718 7528 5724 7540
rect 5399 7500 5724 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6512 7500 6653 7528
rect 6512 7488 6518 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 10042 7528 10048 7540
rect 6641 7491 6699 7497
rect 7208 7500 10048 7528
rect 1946 7460 1952 7472
rect 1907 7432 1952 7460
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 2958 7420 2964 7472
rect 3016 7420 3022 7472
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 3936 7432 4077 7460
rect 3936 7420 3942 7432
rect 4065 7429 4077 7432
rect 4111 7429 4123 7463
rect 4065 7423 4123 7429
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 1636 7364 1685 7392
rect 1636 7352 1642 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7392 4675 7395
rect 5074 7392 5080 7404
rect 4663 7364 5080 7392
rect 4663 7361 4675 7364
rect 4617 7355 4675 7361
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3988 7324 4016 7355
rect 5074 7352 5080 7364
rect 5132 7392 5138 7404
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 5132 7364 5273 7392
rect 5132 7352 5138 7364
rect 5261 7361 5273 7364
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6512 7364 6561 7392
rect 6512 7352 6518 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7208 7401 7236 7500
rect 7469 7463 7527 7469
rect 7469 7429 7481 7463
rect 7515 7460 7527 7463
rect 7742 7460 7748 7472
rect 7515 7432 7748 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 8478 7420 8484 7472
rect 8536 7420 8542 7472
rect 9416 7401 9444 7500
rect 10042 7488 10048 7500
rect 10100 7528 10106 7540
rect 10318 7528 10324 7540
rect 10100 7500 10324 7528
rect 10100 7488 10106 7500
rect 10318 7488 10324 7500
rect 10376 7528 10382 7540
rect 10376 7500 11100 7528
rect 10376 7488 10382 7500
rect 9677 7463 9735 7469
rect 9677 7429 9689 7463
rect 9723 7460 9735 7463
rect 9950 7460 9956 7472
rect 9723 7432 9956 7460
rect 9723 7429 9735 7432
rect 9677 7423 9735 7429
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6972 7364 7205 7392
rect 6972 7352 6978 7364
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 11072 7392 11100 7500
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 11848 7500 13461 7528
rect 11848 7488 11854 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 11204 7432 12466 7460
rect 11204 7420 11210 7432
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 9401 7355 9459 7361
rect 3200 7296 4016 7324
rect 3200 7284 3206 7296
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 10796 7324 10824 7378
rect 11072 7364 11713 7392
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 15896 7364 16865 7392
rect 15896 7352 15902 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 36354 7392 36360 7404
rect 36315 7364 36360 7392
rect 16853 7355 16911 7361
rect 36354 7352 36360 7364
rect 36412 7352 36418 7404
rect 7616 7296 10824 7324
rect 7616 7284 7622 7296
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11020 7296 11989 7324
rect 11020 7284 11026 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 4709 7259 4767 7265
rect 4709 7225 4721 7259
rect 4755 7256 4767 7259
rect 4798 7256 4804 7268
rect 4755 7228 4804 7256
rect 4755 7225 4767 7228
rect 4709 7219 4767 7225
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 8938 7188 8944 7200
rect 8899 7160 8944 7188
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10836 7160 11161 7188
rect 10836 7148 10842 7160
rect 11149 7157 11161 7160
rect 11195 7188 11207 7191
rect 15654 7188 15660 7200
rect 11195 7160 15660 7188
rect 11195 7157 11207 7160
rect 11149 7151 11207 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16945 7191 17003 7197
rect 16945 7157 16957 7191
rect 16991 7188 17003 7191
rect 17862 7188 17868 7200
rect 16991 7160 17868 7188
rect 16991 7157 17003 7160
rect 16945 7151 17003 7157
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 36173 7191 36231 7197
rect 36173 7157 36185 7191
rect 36219 7188 36231 7191
rect 38010 7188 38016 7200
rect 36219 7160 38016 7188
rect 36219 7157 36231 7160
rect 36173 7151 36231 7157
rect 38010 7148 38016 7160
rect 38068 7148 38074 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2004 6956 2912 6984
rect 2004 6944 2010 6956
rect 1854 6876 1860 6928
rect 1912 6916 1918 6928
rect 2406 6916 2412 6928
rect 1912 6888 2412 6916
rect 1912 6876 1918 6888
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 2884 6848 2912 6956
rect 3786 6944 3792 6996
rect 3844 6984 3850 6996
rect 5350 6984 5356 6996
rect 3844 6956 5356 6984
rect 3844 6944 3850 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 8938 6944 8944 6996
rect 8996 6984 9002 6996
rect 10394 6987 10452 6993
rect 10394 6984 10406 6987
rect 8996 6956 10406 6984
rect 8996 6944 9002 6956
rect 10394 6953 10406 6956
rect 10440 6984 10452 6987
rect 14458 6984 14464 6996
rect 10440 6956 14464 6984
rect 10440 6953 10452 6956
rect 10394 6947 10452 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 4672 6888 8340 6916
rect 4672 6876 4678 6888
rect 3234 6848 3240 6860
rect 1544 6820 2774 6848
rect 2884 6820 3240 6848
rect 1544 6808 1550 6820
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6780 1823 6783
rect 1946 6780 1952 6792
rect 1811 6752 1952 6780
rect 1811 6749 1823 6752
rect 1765 6743 1823 6749
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 2096 6752 2329 6780
rect 2096 6740 2102 6752
rect 2317 6749 2329 6752
rect 2363 6749 2375 6783
rect 2746 6780 2774 6820
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 5718 6848 5724 6860
rect 4080 6820 5724 6848
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2746 6752 2973 6780
rect 2317 6743 2375 6749
rect 2961 6749 2973 6752
rect 3007 6780 3019 6783
rect 3050 6780 3056 6792
rect 3007 6752 3056 6780
rect 3007 6749 3019 6752
rect 2961 6743 3019 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 4080 6789 4108 6820
rect 5718 6808 5724 6820
rect 5776 6808 5782 6860
rect 5994 6848 6000 6860
rect 5955 6820 6000 6848
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6638 6848 6644 6860
rect 6599 6820 6644 6848
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 8312 6848 8340 6888
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9088 6888 9444 6916
rect 9088 6876 9094 6888
rect 9416 6848 9444 6888
rect 9968 6888 10272 6916
rect 9858 6848 9864 6860
rect 6880 6820 8248 6848
rect 8312 6820 9260 6848
rect 9416 6820 9864 6848
rect 6880 6808 6886 6820
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3568 6752 3985 6780
rect 3568 6740 3574 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4065 6743 4123 6749
rect 4614 6740 4620 6752
rect 4672 6780 4678 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4672 6752 5273 6780
rect 4672 6740 4678 6752
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 6086 6780 6092 6792
rect 5951 6752 6092 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6454 6740 6460 6792
rect 6512 6780 6518 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 6512 6752 6561 6780
rect 6512 6740 6518 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6730 6740 6736 6792
rect 6788 6780 6794 6792
rect 8220 6789 8248 6820
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 6788 6752 7573 6780
rect 6788 6740 6794 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 9122 6780 9128 6792
rect 8343 6752 9128 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9232 6780 9260 6820
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9232 6752 9321 6780
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9968 6780 9996 6888
rect 10042 6808 10048 6860
rect 10100 6848 10106 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 10100 6820 10149 6848
rect 10100 6808 10106 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10244 6848 10272 6888
rect 11882 6848 11888 6860
rect 10244 6820 11888 6848
rect 10137 6811 10195 6817
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12526 6848 12532 6860
rect 12487 6820 12532 6848
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 25406 6848 25412 6860
rect 25367 6820 25412 6848
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 9456 6752 9996 6780
rect 12437 6783 12495 6789
rect 9456 6740 9462 6752
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 25317 6783 25375 6789
rect 25317 6749 25329 6783
rect 25363 6780 25375 6783
rect 27522 6780 27528 6792
rect 25363 6752 27528 6780
rect 25363 6749 25375 6752
rect 25317 6743 25375 6749
rect 1596 6684 9352 6712
rect 1596 6653 1624 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2409 6647 2467 6653
rect 2409 6644 2421 6647
rect 2280 6616 2421 6644
rect 2280 6604 2286 6616
rect 2409 6613 2421 6616
rect 2455 6613 2467 6647
rect 2409 6607 2467 6613
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3234 6644 3240 6656
rect 3099 6616 3240 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 4798 6644 4804 6656
rect 4755 6616 4804 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5442 6644 5448 6656
rect 5399 6616 5448 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 7190 6644 7196 6656
rect 5776 6616 7196 6644
rect 5776 6604 5782 6616
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 9030 6644 9036 6656
rect 7699 6616 9036 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9324 6644 9352 6684
rect 11054 6672 11060 6724
rect 11112 6672 11118 6724
rect 12342 6712 12348 6724
rect 11716 6684 12348 6712
rect 11716 6644 11744 6684
rect 12342 6672 12348 6684
rect 12400 6672 12406 6724
rect 9180 6616 9225 6644
rect 9324 6616 11744 6644
rect 11885 6647 11943 6653
rect 9180 6604 9186 6616
rect 11885 6613 11897 6647
rect 11931 6644 11943 6647
rect 11974 6644 11980 6656
rect 11931 6616 11980 6644
rect 11931 6613 11943 6616
rect 11885 6607 11943 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12158 6604 12164 6656
rect 12216 6644 12222 6656
rect 12452 6644 12480 6743
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 34146 6780 34152 6792
rect 34107 6752 34152 6780
rect 34146 6740 34152 6752
rect 34204 6740 34210 6792
rect 12216 6616 12480 6644
rect 33965 6647 34023 6653
rect 12216 6604 12222 6616
rect 33965 6613 33977 6647
rect 34011 6644 34023 6647
rect 36998 6644 37004 6656
rect 34011 6616 37004 6644
rect 34011 6613 34023 6616
rect 33965 6607 34023 6613
rect 36998 6604 37004 6616
rect 37056 6604 37062 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 2130 6440 2136 6452
rect 1627 6412 2136 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 3142 6440 3148 6452
rect 3103 6412 3148 6440
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3786 6440 3792 6452
rect 3747 6412 3792 6440
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 5902 6440 5908 6452
rect 4080 6412 5908 6440
rect 2222 6332 2228 6384
rect 2280 6372 2286 6384
rect 4080 6372 4108 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6409 6699 6443
rect 6641 6403 6699 6409
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 7926 6440 7932 6452
rect 7791 6412 7932 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 5718 6372 5724 6384
rect 2280 6344 4108 6372
rect 4172 6344 5724 6372
rect 2280 6332 2286 6344
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 3050 6304 3056 6316
rect 2963 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 3142 6264 3148 6316
rect 3200 6304 3206 6316
rect 3694 6304 3700 6316
rect 3200 6276 3700 6304
rect 3200 6264 3206 6276
rect 3694 6264 3700 6276
rect 3752 6304 3758 6316
rect 4172 6304 4200 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 6656 6372 6684 6403
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 10042 6440 10048 6452
rect 8956 6412 10048 6440
rect 8662 6372 8668 6384
rect 6656 6344 8668 6372
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 4614 6304 4620 6316
rect 3752 6276 4200 6304
rect 4527 6276 4620 6304
rect 3752 6264 3758 6276
rect 4614 6264 4620 6276
rect 4672 6304 4678 6316
rect 5258 6304 5264 6316
rect 4672 6276 5264 6304
rect 4672 6264 4678 6276
rect 5258 6264 5264 6276
rect 5316 6304 5322 6316
rect 6454 6304 6460 6316
rect 5316 6276 6460 6304
rect 5316 6264 5322 6276
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 7190 6304 7196 6316
rect 6595 6276 7196 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 3068 6236 3096 6264
rect 4706 6236 4712 6248
rect 3068 6208 4712 6236
rect 4706 6196 4712 6208
rect 4764 6236 4770 6248
rect 5074 6236 5080 6248
rect 4764 6208 5080 6236
rect 4764 6196 4770 6208
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 7668 6236 7696 6267
rect 7926 6264 7932 6316
rect 7984 6304 7990 6316
rect 8956 6313 8984 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 11422 6440 11428 6452
rect 10735 6412 11428 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 9272 6344 9706 6372
rect 9272 6332 9278 6344
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 7984 6276 8309 6304
rect 7984 6264 7990 6276
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8941 6307 8999 6313
rect 8941 6273 8953 6307
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 5500 6208 7696 6236
rect 9217 6239 9275 6245
rect 5500 6196 5506 6208
rect 9217 6205 9229 6239
rect 9263 6236 9275 6239
rect 9674 6236 9680 6248
rect 9263 6208 9680 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 4614 6128 4620 6180
rect 4672 6168 4678 6180
rect 8938 6168 8944 6180
rect 4672 6140 8944 6168
rect 4672 6128 4678 6140
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 4982 6100 4988 6112
rect 4755 6072 4988 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 7926 6100 7932 6112
rect 5776 6072 7932 6100
rect 5776 6060 5782 6072
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 10704 6100 10732 6403
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13504 6412 13921 6440
rect 13504 6400 13510 6412
rect 13909 6409 13921 6412
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 18417 6443 18475 6449
rect 18417 6440 18429 6443
rect 18288 6412 18429 6440
rect 18288 6400 18294 6412
rect 18417 6409 18429 6412
rect 18463 6409 18475 6443
rect 18417 6403 18475 6409
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 22097 6443 22155 6449
rect 22097 6440 22109 6443
rect 21324 6412 22109 6440
rect 21324 6400 21330 6412
rect 22097 6409 22109 6412
rect 22143 6409 22155 6443
rect 38102 6440 38108 6452
rect 38063 6412 38108 6440
rect 22097 6403 22155 6409
rect 38102 6400 38108 6412
rect 38160 6400 38166 6452
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 14918 6304 14924 6316
rect 13863 6276 14924 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 18322 6304 18328 6316
rect 18283 6276 18328 6304
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 22005 6307 22063 6313
rect 22005 6273 22017 6307
rect 22051 6304 22063 6307
rect 22646 6304 22652 6316
rect 22051 6276 22652 6304
rect 22051 6273 22063 6276
rect 22005 6267 22063 6273
rect 22646 6264 22652 6276
rect 22704 6264 22710 6316
rect 31021 6307 31079 6313
rect 31021 6273 31033 6307
rect 31067 6304 31079 6307
rect 32858 6304 32864 6316
rect 31067 6276 32864 6304
rect 31067 6273 31079 6276
rect 31021 6267 31079 6273
rect 32858 6264 32864 6276
rect 32916 6264 32922 6316
rect 32953 6307 33011 6313
rect 32953 6273 32965 6307
rect 32999 6304 33011 6307
rect 35618 6304 35624 6316
rect 32999 6276 35624 6304
rect 32999 6273 33011 6276
rect 32953 6267 33011 6273
rect 35618 6264 35624 6276
rect 35676 6264 35682 6316
rect 38286 6304 38292 6316
rect 38247 6276 38292 6304
rect 38286 6264 38292 6276
rect 38344 6264 38350 6316
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 33045 6239 33103 6245
rect 33045 6236 33057 6239
rect 18472 6208 33057 6236
rect 18472 6196 18478 6208
rect 33045 6205 33057 6208
rect 33091 6205 33103 6239
rect 33045 6199 33103 6205
rect 24670 6128 24676 6180
rect 24728 6168 24734 6180
rect 31113 6171 31171 6177
rect 31113 6168 31125 6171
rect 24728 6140 31125 6168
rect 24728 6128 24734 6140
rect 31113 6137 31125 6140
rect 31159 6137 31171 6171
rect 31113 6131 31171 6137
rect 8352 6072 10732 6100
rect 8352 6060 8358 6072
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2590 5896 2596 5908
rect 2455 5868 2596 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2590 5856 2596 5868
rect 2648 5856 2654 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 4028 5868 4077 5896
rect 4028 5856 4034 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4709 5899 4767 5905
rect 4709 5896 4721 5899
rect 4212 5868 4721 5896
rect 4212 5856 4218 5868
rect 4709 5865 4721 5868
rect 4755 5865 4767 5899
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 4709 5859 4767 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5997 5899 6055 5905
rect 5997 5865 6009 5899
rect 6043 5896 6055 5899
rect 7282 5896 7288 5908
rect 6043 5868 7288 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 9214 5896 9220 5908
rect 7392 5868 9220 5896
rect 1765 5831 1823 5837
rect 1765 5797 1777 5831
rect 1811 5828 1823 5831
rect 2958 5828 2964 5840
rect 1811 5800 2964 5828
rect 1811 5797 1823 5800
rect 1765 5791 1823 5797
rect 2958 5788 2964 5800
rect 3016 5788 3022 5840
rect 6270 5788 6276 5840
rect 6328 5828 6334 5840
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 6328 5800 6653 5828
rect 6328 5788 6334 5800
rect 6641 5797 6653 5800
rect 6687 5797 6699 5831
rect 7392 5828 7420 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 11241 5899 11299 5905
rect 11241 5896 11253 5899
rect 10744 5868 11253 5896
rect 10744 5856 10750 5868
rect 11241 5865 11253 5868
rect 11287 5865 11299 5899
rect 11241 5859 11299 5865
rect 6641 5791 6699 5797
rect 6748 5800 7420 5828
rect 8113 5831 8171 5837
rect 2498 5720 2504 5772
rect 2556 5760 2562 5772
rect 2556 5732 4016 5760
rect 2556 5720 2562 5732
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2038 5692 2044 5704
rect 1719 5664 2044 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2406 5692 2412 5704
rect 2363 5664 2412 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3142 5692 3148 5704
rect 2746 5664 3148 5692
rect 2056 5624 2084 5652
rect 2746 5624 2774 5664
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3988 5701 4016 5732
rect 4632 5732 5948 5760
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4632 5701 4660 5732
rect 4617 5695 4675 5701
rect 4617 5692 4629 5695
rect 4304 5664 4629 5692
rect 4304 5652 4310 5664
rect 4617 5661 4629 5664
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5350 5692 5356 5704
rect 5307 5664 5356 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 5920 5701 5948 5732
rect 5994 5720 6000 5772
rect 6052 5760 6058 5772
rect 6748 5760 6776 5800
rect 8113 5797 8125 5831
rect 8159 5828 8171 5831
rect 11330 5828 11336 5840
rect 8159 5800 11336 5828
rect 8159 5797 8171 5800
rect 8113 5791 8171 5797
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 6052 5732 6776 5760
rect 7285 5763 7343 5769
rect 6052 5720 6058 5732
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 7466 5760 7472 5772
rect 7331 5732 7472 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6086 5692 6092 5704
rect 5951 5664 6092 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6086 5652 6092 5664
rect 6144 5692 6150 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6144 5664 6561 5692
rect 6144 5652 6150 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 6549 5655 6607 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 11146 5692 11152 5704
rect 11107 5664 11152 5692
rect 8021 5655 8079 5661
rect 2056 5596 2774 5624
rect 3237 5627 3295 5633
rect 3237 5593 3249 5627
rect 3283 5624 3295 5627
rect 3283 5596 4844 5624
rect 3283 5593 3295 5596
rect 3237 5587 3295 5593
rect 4816 5556 4844 5596
rect 5718 5584 5724 5636
rect 5776 5624 5782 5636
rect 8036 5624 8064 5655
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 13722 5692 13728 5704
rect 12023 5664 13728 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 17862 5692 17868 5704
rect 17823 5664 17868 5692
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18506 5692 18512 5704
rect 18467 5664 18512 5692
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 21174 5692 21180 5704
rect 21135 5664 21180 5692
rect 21174 5652 21180 5664
rect 21232 5652 21238 5704
rect 23566 5692 23572 5704
rect 23527 5664 23572 5692
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 5776 5596 8064 5624
rect 5776 5584 5782 5596
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 12069 5627 12127 5633
rect 12069 5624 12081 5627
rect 10100 5596 12081 5624
rect 10100 5584 10106 5596
rect 12069 5593 12081 5596
rect 12115 5593 12127 5627
rect 12069 5587 12127 5593
rect 6178 5556 6184 5568
rect 4816 5528 6184 5556
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 7742 5556 7748 5568
rect 6512 5528 7748 5556
rect 6512 5516 6518 5528
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 17681 5559 17739 5565
rect 17681 5525 17693 5559
rect 17727 5556 17739 5559
rect 18138 5556 18144 5568
rect 17727 5528 18144 5556
rect 17727 5525 17739 5528
rect 17681 5519 17739 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18325 5559 18383 5565
rect 18325 5525 18337 5559
rect 18371 5556 18383 5559
rect 19426 5556 19432 5568
rect 18371 5528 19432 5556
rect 18371 5525 18383 5528
rect 18325 5519 18383 5525
rect 19426 5516 19432 5528
rect 19484 5516 19490 5568
rect 20993 5559 21051 5565
rect 20993 5525 21005 5559
rect 21039 5556 21051 5559
rect 23290 5556 23296 5568
rect 21039 5528 23296 5556
rect 21039 5525 21051 5528
rect 20993 5519 21051 5525
rect 23290 5516 23296 5528
rect 23348 5516 23354 5568
rect 23385 5559 23443 5565
rect 23385 5525 23397 5559
rect 23431 5556 23443 5559
rect 24762 5556 24768 5568
rect 23431 5528 24768 5556
rect 23431 5525 23443 5528
rect 23385 5519 23443 5525
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2409 5355 2467 5361
rect 2409 5352 2421 5355
rect 2372 5324 2421 5352
rect 2372 5312 2378 5324
rect 2409 5321 2421 5324
rect 2455 5321 2467 5355
rect 3694 5352 3700 5364
rect 3655 5324 3700 5352
rect 2409 5315 2467 5321
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 4338 5352 4344 5364
rect 4299 5324 4344 5352
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7156 5324 9628 5352
rect 7156 5312 7162 5324
rect 3053 5287 3111 5293
rect 3053 5253 3065 5287
rect 3099 5284 3111 5287
rect 5626 5284 5632 5296
rect 3099 5256 5632 5284
rect 3099 5253 3111 5256
rect 3053 5247 3111 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 8849 5287 8907 5293
rect 8849 5284 8861 5287
rect 6748 5256 8861 5284
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2406 5216 2412 5228
rect 2363 5188 2412 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 1596 5148 1624 5179
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 2958 5216 2964 5228
rect 2871 5188 2964 5216
rect 2958 5176 2964 5188
rect 3016 5216 3022 5228
rect 3510 5216 3516 5228
rect 3016 5188 3516 5216
rect 3016 5176 3022 5188
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3694 5216 3700 5228
rect 3651 5188 3700 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 4246 5176 4252 5228
rect 4304 5225 4310 5228
rect 4304 5216 4315 5225
rect 4304 5188 4349 5216
rect 4304 5179 4315 5188
rect 4304 5176 4310 5179
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 4893 5219 4951 5225
rect 4893 5216 4905 5219
rect 4856 5188 4905 5216
rect 4856 5176 4862 5188
rect 4893 5185 4905 5188
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 6748 5225 6776 5256
rect 8849 5253 8861 5256
rect 8895 5253 8907 5287
rect 8849 5247 8907 5253
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 5132 5188 5549 5216
rect 5132 5176 5138 5188
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7239 5188 7696 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7668 5148 7696 5188
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7800 5188 7849 5216
rect 7800 5176 7806 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 9600 5225 9628 5324
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8260 5188 8769 5216
rect 8260 5176 8266 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 29638 5176 29644 5228
rect 29696 5216 29702 5228
rect 33781 5219 33839 5225
rect 33781 5216 33793 5219
rect 29696 5188 33793 5216
rect 29696 5176 29702 5188
rect 33781 5185 33793 5188
rect 33827 5185 33839 5219
rect 33781 5179 33839 5185
rect 13078 5148 13084 5160
rect 1596 5120 6592 5148
rect 7668 5120 13084 5148
rect 2406 5040 2412 5092
rect 2464 5080 2470 5092
rect 4246 5080 4252 5092
rect 2464 5052 4252 5080
rect 2464 5040 2470 5052
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 6564 5089 6592 5120
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 6549 5083 6607 5089
rect 6549 5049 6561 5083
rect 6595 5049 6607 5083
rect 7929 5083 7987 5089
rect 6549 5043 6607 5049
rect 7116 5052 7420 5080
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4982 5012 4988 5024
rect 3936 4984 4988 5012
rect 3936 4972 3942 4984
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5629 5015 5687 5021
rect 5629 4981 5641 5015
rect 5675 5012 5687 5015
rect 7116 5012 7144 5052
rect 7282 5012 7288 5024
rect 5675 4984 7144 5012
rect 7243 4984 7288 5012
rect 5675 4981 5687 4984
rect 5629 4975 5687 4981
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7392 5012 7420 5052
rect 7929 5049 7941 5083
rect 7975 5080 7987 5083
rect 11238 5080 11244 5092
rect 7975 5052 11244 5080
rect 7975 5049 7987 5052
rect 7929 5043 7987 5049
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 8846 5012 8852 5024
rect 7392 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 9401 5015 9459 5021
rect 9401 5012 9413 5015
rect 9180 4984 9413 5012
rect 9180 4972 9186 4984
rect 9401 4981 9413 4984
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 33597 5015 33655 5021
rect 33597 4981 33609 5015
rect 33643 5012 33655 5015
rect 36906 5012 36912 5024
rect 33643 4984 36912 5012
rect 33643 4981 33655 4984
rect 33597 4975 33655 4981
rect 36906 4972 36912 4984
rect 36964 4972 36970 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2685 4811 2743 4817
rect 2685 4777 2697 4811
rect 2731 4808 2743 4811
rect 2866 4808 2872 4820
rect 2731 4780 2872 4808
rect 2731 4777 2743 4780
rect 2685 4771 2743 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 5629 4811 5687 4817
rect 3375 4780 5580 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 1949 4743 2007 4749
rect 1949 4709 1961 4743
rect 1995 4740 2007 4743
rect 3878 4740 3884 4752
rect 1995 4712 3884 4740
rect 1995 4709 2007 4712
rect 1949 4703 2007 4709
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4706 4740 4712 4752
rect 4080 4712 4712 4740
rect 2958 4672 2964 4684
rect 2746 4644 2964 4672
rect 1854 4604 1860 4616
rect 1815 4576 1860 4604
rect 1854 4564 1860 4576
rect 1912 4564 1918 4616
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 2746 4604 2774 4644
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 2639 4576 2774 4604
rect 3237 4607 3295 4613
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 4080 4604 4108 4712
rect 4706 4700 4712 4712
rect 4764 4740 4770 4752
rect 5258 4740 5264 4752
rect 4764 4712 5264 4740
rect 4764 4700 4770 4712
rect 5258 4700 5264 4712
rect 5316 4700 5322 4752
rect 5552 4740 5580 4780
rect 5629 4777 5641 4811
rect 5675 4808 5687 4811
rect 6546 4808 6552 4820
rect 5675 4780 6552 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7558 4808 7564 4820
rect 6963 4780 7564 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 12802 4808 12808 4820
rect 10091 4780 12808 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 6273 4743 6331 4749
rect 5552 4712 6224 4740
rect 4246 4672 4252 4684
rect 4207 4644 4252 4672
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 6196 4672 6224 4712
rect 6273 4709 6285 4743
rect 6319 4740 6331 4743
rect 10870 4740 10876 4752
rect 6319 4712 10876 4740
rect 6319 4709 6331 4712
rect 6273 4703 6331 4709
rect 10870 4700 10876 4712
rect 10928 4700 10934 4752
rect 10962 4672 10968 4684
rect 4908 4644 5764 4672
rect 6196 4644 10968 4672
rect 3283 4576 4108 4604
rect 4157 4607 4215 4613
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4798 4604 4804 4616
rect 4203 4576 4804 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3694 4536 3700 4548
rect 3016 4508 3700 4536
rect 3016 4496 3022 4508
rect 3694 4496 3700 4508
rect 3752 4536 3758 4548
rect 4172 4536 4200 4567
rect 4798 4564 4804 4576
rect 4856 4604 4862 4616
rect 4908 4613 4936 4644
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4856 4576 4905 4604
rect 4856 4564 4862 4576
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5408 4576 5549 4604
rect 5408 4564 5414 4576
rect 5537 4573 5549 4576
rect 5583 4604 5595 4607
rect 5626 4604 5632 4616
rect 5583 4576 5632 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5736 4604 5764 4644
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5736 4576 6193 4604
rect 6181 4573 6193 4576
rect 6227 4604 6239 4607
rect 6825 4607 6883 4613
rect 6825 4604 6837 4607
rect 6227 4576 6837 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6825 4573 6837 4576
rect 6871 4604 6883 4607
rect 7190 4604 7196 4616
rect 6871 4576 7196 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 3752 4508 4200 4536
rect 3752 4496 3758 4508
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 9968 4536 9996 4567
rect 22830 4564 22836 4616
rect 22888 4604 22894 4616
rect 26237 4607 26295 4613
rect 26237 4604 26249 4607
rect 22888 4576 26249 4604
rect 22888 4564 22894 4576
rect 26237 4573 26249 4576
rect 26283 4573 26295 4607
rect 38010 4604 38016 4616
rect 37971 4576 38016 4604
rect 26237 4567 26295 4573
rect 38010 4564 38016 4576
rect 38068 4564 38074 4616
rect 4764 4508 9996 4536
rect 4764 4496 4770 4508
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 7834 4468 7840 4480
rect 5031 4440 7840 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 26329 4471 26387 4477
rect 26329 4437 26341 4471
rect 26375 4468 26387 4471
rect 28166 4468 28172 4480
rect 26375 4440 28172 4468
rect 26375 4437 26387 4440
rect 26329 4431 26387 4437
rect 28166 4428 28172 4440
rect 28224 4428 28230 4480
rect 38194 4468 38200 4480
rect 38155 4440 38200 4468
rect 38194 4428 38200 4440
rect 38252 4428 38258 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 3326 4264 3332 4276
rect 2363 4236 3332 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 1854 4156 1860 4208
rect 1912 4196 1918 4208
rect 2958 4196 2964 4208
rect 1912 4168 2964 4196
rect 1912 4156 1918 4168
rect 2240 4137 2268 4168
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 3878 4156 3884 4208
rect 3936 4196 3942 4208
rect 5626 4196 5632 4208
rect 3936 4168 5632 4196
rect 3936 4156 3942 4168
rect 5626 4156 5632 4168
rect 5684 4196 5690 4208
rect 5684 4168 5764 4196
rect 5684 4156 5690 4168
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4097 2283 4131
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2225 4091 2283 4097
rect 1780 4060 1808 4091
rect 2866 4088 2872 4100
rect 2924 4128 2930 4140
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 2924 4100 3525 4128
rect 2924 4088 2930 4100
rect 3513 4097 3525 4100
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 4433 4131 4491 4137
rect 3660 4100 3705 4128
rect 3660 4088 3666 4100
rect 4433 4097 4445 4131
rect 4479 4128 4491 4131
rect 4614 4128 4620 4140
rect 4479 4100 4620 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 5074 4128 5080 4140
rect 5035 4100 5080 4128
rect 5074 4088 5080 4100
rect 5132 4088 5138 4140
rect 5736 4137 5764 4168
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 5994 4128 6000 4140
rect 5859 4100 6000 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 2774 4060 2780 4072
rect 1780 4032 2780 4060
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4060 3019 4063
rect 3418 4060 3424 4072
rect 3007 4032 3424 4060
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 3418 4020 3424 4032
rect 3476 4020 3482 4072
rect 4522 4060 4528 4072
rect 4483 4032 4528 4060
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4060 5227 4063
rect 11054 4060 11060 4072
rect 5215 4032 11060 4060
rect 5215 4029 5227 4032
rect 5169 4023 5227 4029
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 2682 3992 2688 4004
rect 1627 3964 2688 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 2682 3952 2688 3964
rect 2740 3952 2746 4004
rect 3234 3952 3240 4004
rect 3292 3992 3298 4004
rect 8110 3992 8116 4004
rect 3292 3964 8116 3992
rect 3292 3952 3298 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1765 3723 1823 3729
rect 1765 3689 1777 3723
rect 1811 3720 1823 3723
rect 3234 3720 3240 3732
rect 1811 3692 3240 3720
rect 1811 3689 1823 3692
rect 1765 3683 1823 3689
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3329 3723 3387 3729
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 5166 3720 5172 3732
rect 3375 3692 5172 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6365 3723 6423 3729
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 6822 3720 6828 3732
rect 6411 3692 6828 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 33962 3680 33968 3732
rect 34020 3720 34026 3732
rect 38105 3723 38163 3729
rect 38105 3720 38117 3723
rect 34020 3692 38117 3720
rect 34020 3680 34026 3692
rect 38105 3689 38117 3692
rect 38151 3689 38163 3723
rect 38105 3683 38163 3689
rect 3142 3652 3148 3664
rect 2240 3624 3148 3652
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 2240 3516 2268 3624
rect 3142 3612 3148 3624
rect 3200 3652 3206 3664
rect 3970 3652 3976 3664
rect 3200 3624 3976 3652
rect 3200 3612 3206 3624
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 4065 3655 4123 3661
rect 4065 3621 4077 3655
rect 4111 3652 4123 3655
rect 5534 3652 5540 3664
rect 4111 3624 5540 3652
rect 4111 3621 4123 3624
rect 4065 3615 4123 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 2590 3544 2596 3596
rect 2648 3584 2654 3596
rect 2648 3556 5948 3584
rect 2648 3544 2654 3556
rect 1719 3488 2268 3516
rect 2317 3519 2375 3525
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 2317 3485 2329 3519
rect 2363 3516 2375 3519
rect 2498 3516 2504 3528
rect 2363 3488 2504 3516
rect 2363 3485 2375 3488
rect 2317 3479 2375 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2924 3488 3249 3516
rect 2924 3476 2930 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3237 3479 3295 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 5074 3516 5080 3528
rect 4080 3488 5080 3516
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 2593 3451 2651 3457
rect 2593 3448 2605 3451
rect 2464 3420 2605 3448
rect 2464 3408 2470 3420
rect 2593 3417 2605 3420
rect 2639 3448 2651 3451
rect 4080 3448 4108 3488
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5920 3525 5948 3556
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3485 6607 3519
rect 38286 3516 38292 3528
rect 38247 3488 38292 3516
rect 6549 3479 6607 3485
rect 2639 3420 4108 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 6564 3448 6592 3479
rect 38286 3476 38292 3488
rect 38344 3476 38350 3528
rect 4212 3420 6592 3448
rect 4212 3408 4218 3420
rect 5169 3383 5227 3389
rect 5169 3349 5181 3383
rect 5215 3380 5227 3383
rect 8478 3380 8484 3392
rect 5215 3352 8484 3380
rect 5215 3349 5227 3352
rect 5169 3343 5227 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5166 3176 5172 3188
rect 2746 3148 5172 3176
rect 2746 3108 2774 3148
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 6549 3179 6607 3185
rect 5316 3148 5361 3176
rect 5316 3136 5322 3148
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6730 3176 6736 3188
rect 6595 3148 6736 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 35618 3136 35624 3188
rect 35676 3176 35682 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 35676 3148 36737 3176
rect 35676 3136 35682 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 2958 3108 2964 3120
rect 2700 3080 2774 3108
rect 2919 3080 2964 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1596 2972 1624 3003
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 2700 3049 2728 3080
rect 2958 3068 2964 3080
rect 3016 3068 3022 3120
rect 3970 3068 3976 3120
rect 4028 3108 4034 3120
rect 4028 3080 6776 3108
rect 4028 3068 4034 3080
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2556 3012 2697 3040
rect 2556 3000 2562 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 3786 3040 3792 3052
rect 3747 3012 3792 3040
rect 2685 3003 2743 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 5166 3040 5172 3052
rect 5079 3012 5172 3040
rect 4249 3003 4307 3009
rect 2774 2972 2780 2984
rect 1596 2944 2780 2972
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 4264 2972 4292 3003
rect 5166 3000 5172 3012
rect 5224 3040 5230 3052
rect 5350 3040 5356 3052
rect 5224 3012 5356 3040
rect 5224 3000 5230 3012
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 6748 3049 6776 3080
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 10042 3040 10048 3052
rect 10003 3012 10048 3040
rect 6733 3003 6791 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 28166 3040 28172 3052
rect 28127 3012 28172 3040
rect 28166 3000 28172 3012
rect 28224 3000 28230 3052
rect 36909 3043 36967 3049
rect 36909 3009 36921 3043
rect 36955 3009 36967 3043
rect 36909 3003 36967 3009
rect 15010 2972 15016 2984
rect 4264 2944 15016 2972
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 36924 2972 36952 3003
rect 36998 3000 37004 3052
rect 37056 3040 37062 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37056 3012 38025 3040
rect 37056 3000 37062 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 39298 2972 39304 2984
rect 36924 2944 39304 2972
rect 39298 2932 39304 2944
rect 39356 2932 39362 2984
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 4706 2904 4712 2916
rect 3651 2876 4712 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 72 2808 1777 2836
rect 72 2796 78 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 1765 2799 1823 2805
rect 4341 2839 4399 2845
rect 4341 2805 4353 2839
rect 4387 2836 4399 2839
rect 4614 2836 4620 2848
rect 4387 2808 4620 2836
rect 4387 2805 4399 2808
rect 4341 2799 4399 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 9861 2839 9919 2845
rect 9861 2836 9873 2839
rect 7064 2808 9873 2836
rect 7064 2796 7070 2808
rect 9861 2805 9873 2808
rect 9907 2805 9919 2839
rect 9861 2799 9919 2805
rect 27985 2839 28043 2845
rect 27985 2805 27997 2839
rect 28031 2836 28043 2839
rect 30190 2836 30196 2848
rect 28031 2808 30196 2836
rect 28031 2805 28043 2808
rect 27985 2799 28043 2805
rect 30190 2796 30196 2808
rect 30248 2796 30254 2848
rect 38194 2836 38200 2848
rect 38155 2808 38200 2836
rect 38194 2796 38200 2808
rect 38252 2796 38258 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 2832 2604 3985 2632
rect 2832 2592 2838 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 5442 2632 5448 2644
rect 4663 2604 5448 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7374 2632 7380 2644
rect 7331 2604 7380 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11204 2604 11713 2632
rect 11204 2592 11210 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 14277 2635 14335 2641
rect 14277 2601 14289 2635
rect 14323 2632 14335 2635
rect 14642 2632 14648 2644
rect 14323 2604 14648 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 16853 2635 16911 2641
rect 16853 2601 16865 2635
rect 16899 2632 16911 2635
rect 18322 2632 18328 2644
rect 16899 2604 18328 2632
rect 16899 2601 16911 2604
rect 16853 2595 16911 2601
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 22002 2632 22008 2644
rect 21963 2604 22008 2632
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22646 2632 22652 2644
rect 22607 2604 22652 2632
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 28626 2592 28632 2644
rect 28684 2632 28690 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 28684 2604 29745 2632
rect 28684 2592 28690 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 33594 2632 33600 2644
rect 33555 2604 33600 2632
rect 29733 2595 29791 2601
rect 33594 2592 33600 2604
rect 33652 2592 33658 2644
rect 36173 2635 36231 2641
rect 36173 2632 36185 2635
rect 35866 2604 36185 2632
rect 5261 2567 5319 2573
rect 5261 2533 5273 2567
rect 5307 2533 5319 2567
rect 5261 2527 5319 2533
rect 5276 2496 5304 2527
rect 5350 2524 5356 2576
rect 5408 2564 5414 2576
rect 5408 2536 16574 2564
rect 5408 2524 5414 2536
rect 7282 2496 7288 2508
rect 1596 2468 5304 2496
rect 5460 2468 7288 2496
rect 1596 2437 1624 2468
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 2498 2428 2504 2440
rect 2459 2400 2504 2428
rect 1581 2391 1639 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 3878 2428 3884 2440
rect 2823 2400 3884 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4614 2428 4620 2440
rect 4203 2400 4620 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5460 2437 5488 2468
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 16546 2496 16574 2536
rect 27522 2524 27528 2576
rect 27580 2564 27586 2576
rect 30377 2567 30435 2573
rect 30377 2564 30389 2567
rect 27580 2536 30389 2564
rect 27580 2524 27586 2536
rect 30377 2533 30389 2536
rect 30423 2533 30435 2567
rect 30377 2527 30435 2533
rect 32858 2524 32864 2576
rect 32916 2564 32922 2576
rect 35866 2564 35894 2604
rect 36173 2601 36185 2604
rect 36219 2601 36231 2635
rect 36173 2595 36231 2601
rect 32916 2536 35894 2564
rect 32916 2524 32922 2536
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 16546 2468 27445 2496
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 30190 2456 30196 2508
rect 30248 2496 30254 2508
rect 30248 2468 32352 2496
rect 30248 2456 30254 2468
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 7006 2428 7012 2440
rect 6595 2400 7012 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4816 2360 4844 2391
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7156 2400 7481 2428
rect 7156 2388 7162 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 7469 2391 7527 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10778 2428 10784 2440
rect 10459 2400 10784 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11664 2400 11897 2428
rect 11664 2388 11670 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13596 2400 14473 2428
rect 13596 2388 13602 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 14884 2400 15117 2428
rect 14884 2388 14890 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16816 2400 17049 2428
rect 16816 2388 16822 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 17037 2391 17095 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22612 2400 22845 2428
rect 22612 2388 22618 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23348 2400 24593 2428
rect 23348 2388 23354 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 24820 2400 25881 2428
rect 24820 2388 24826 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 27154 2388 27160 2440
rect 27212 2428 27218 2440
rect 27212 2400 28948 2428
rect 27212 2388 27218 2400
rect 4580 2332 4844 2360
rect 4580 2320 4586 2332
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27249 2363 27307 2369
rect 27249 2360 27261 2363
rect 27120 2332 27261 2360
rect 27120 2320 27126 2332
rect 27249 2329 27261 2332
rect 27295 2329 27307 2363
rect 28920 2360 28948 2400
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 32324 2437 32352 2468
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30340 2400 30573 2428
rect 30340 2388 30346 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 33560 2400 33793 2428
rect 33560 2388 33566 2400
rect 33781 2397 33793 2400
rect 33827 2397 33839 2431
rect 33781 2391 33839 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34848 2400 35081 2428
rect 34848 2388 34854 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35069 2391 35127 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36136 2400 36369 2428
rect 36136 2388 36142 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 36906 2388 36912 2440
rect 36964 2428 36970 2440
rect 38013 2431 38071 2437
rect 38013 2428 38025 2431
rect 36964 2400 38025 2428
rect 36964 2388 36970 2400
rect 38013 2397 38025 2400
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 28920 2332 34928 2360
rect 27249 2323 27307 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 1360 2264 1777 2292
rect 1360 2252 1366 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 1765 2255 1823 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 5868 2264 6745 2292
rect 5868 2252 5874 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9088 2264 9321 2292
rect 9088 2252 9094 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 23900 2264 24777 2292
rect 23900 2252 23906 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 25774 2252 25780 2304
rect 25832 2292 25838 2304
rect 26053 2295 26111 2301
rect 26053 2292 26065 2295
rect 25832 2264 26065 2292
rect 25832 2252 25838 2264
rect 26053 2261 26065 2264
rect 26099 2261 26111 2295
rect 26053 2255 26111 2261
rect 31570 2252 31576 2304
rect 31628 2292 31634 2304
rect 34900 2301 34928 2332
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 31628 2264 32505 2292
rect 31628 2252 31634 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 34885 2295 34943 2301
rect 34885 2261 34897 2295
rect 34931 2261 34943 2295
rect 34885 2255 34943 2261
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38197 2295 38255 2301
rect 38197 2292 38209 2295
rect 38068 2264 38209 2292
rect 38068 2252 38074 2264
rect 38197 2261 38209 2264
rect 38243 2261 38255 2295
rect 38197 2255 38255 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 2780 37204 2832 37256
rect 3148 37247 3200 37256
rect 3148 37213 3157 37247
rect 3157 37213 3191 37247
rect 3191 37213 3200 37247
rect 3148 37204 3200 37213
rect 3240 37204 3292 37256
rect 4620 37204 4672 37256
rect 6552 37247 6604 37256
rect 6552 37213 6561 37247
rect 6561 37213 6595 37247
rect 6595 37213 6604 37247
rect 6552 37204 6604 37213
rect 7840 37247 7892 37256
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 9036 37204 9088 37256
rect 11612 37204 11664 37256
rect 1308 37068 1360 37120
rect 2320 37111 2372 37120
rect 2320 37077 2329 37111
rect 2329 37077 2363 37111
rect 2363 37077 2372 37111
rect 2320 37068 2372 37077
rect 5632 37136 5684 37188
rect 13544 37204 13596 37256
rect 15568 37247 15620 37256
rect 15568 37213 15577 37247
rect 15577 37213 15611 37247
rect 15611 37213 15620 37247
rect 15568 37204 15620 37213
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 18052 37204 18104 37256
rect 18512 37204 18564 37256
rect 20628 37204 20680 37256
rect 22560 37204 22612 37256
rect 24492 37204 24544 37256
rect 25780 37204 25832 37256
rect 27804 37247 27856 37256
rect 27804 37213 27813 37247
rect 27813 37213 27847 37247
rect 27847 37213 27856 37247
rect 27804 37204 27856 37213
rect 27896 37204 27948 37256
rect 30380 37204 30432 37256
rect 32220 37204 32272 37256
rect 33508 37204 33560 37256
rect 34888 37247 34940 37256
rect 34888 37213 34897 37247
rect 34897 37213 34931 37247
rect 34931 37213 34940 37247
rect 34888 37204 34940 37213
rect 36912 37247 36964 37256
rect 36912 37213 36921 37247
rect 36921 37213 36955 37247
rect 36955 37213 36964 37247
rect 36912 37204 36964 37213
rect 37464 37247 37516 37256
rect 37464 37213 37473 37247
rect 37473 37213 37507 37247
rect 37507 37213 37516 37247
rect 37464 37204 37516 37213
rect 14648 37136 14700 37188
rect 15844 37136 15896 37188
rect 3976 37111 4028 37120
rect 3976 37077 3985 37111
rect 3985 37077 4019 37111
rect 4019 37077 4028 37111
rect 3976 37068 4028 37077
rect 4620 37111 4672 37120
rect 4620 37077 4629 37111
rect 4629 37077 4663 37111
rect 4663 37077 4672 37111
rect 4620 37068 4672 37077
rect 5816 37068 5868 37120
rect 7748 37068 7800 37120
rect 9128 37111 9180 37120
rect 9128 37077 9137 37111
rect 9137 37077 9171 37111
rect 9171 37077 9180 37111
rect 9128 37068 9180 37077
rect 10324 37068 10376 37120
rect 12440 37068 12492 37120
rect 14280 37111 14332 37120
rect 14280 37077 14289 37111
rect 14289 37077 14323 37111
rect 14323 37077 14332 37111
rect 14280 37068 14332 37077
rect 15476 37068 15528 37120
rect 16764 37068 16816 37120
rect 20904 37136 20956 37188
rect 19984 37068 20036 37120
rect 21272 37068 21324 37120
rect 28080 37136 28132 37188
rect 23020 37068 23072 37120
rect 25044 37068 25096 37120
rect 27712 37068 27764 37120
rect 29000 37068 29052 37120
rect 30012 37068 30064 37120
rect 30656 37068 30708 37120
rect 34428 37136 34480 37188
rect 34796 37068 34848 37120
rect 36820 37068 36872 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 20 36864 72 36916
rect 3976 36864 4028 36916
rect 10232 36864 10284 36916
rect 27804 36864 27856 36916
rect 34888 36864 34940 36916
rect 9128 36796 9180 36848
rect 13820 36796 13872 36848
rect 39304 36864 39356 36916
rect 3976 36728 4028 36780
rect 8300 36728 8352 36780
rect 25504 36771 25556 36780
rect 25504 36737 25513 36771
rect 25513 36737 25547 36771
rect 25547 36737 25556 36771
rect 25504 36728 25556 36737
rect 29828 36728 29880 36780
rect 31760 36728 31812 36780
rect 36176 36771 36228 36780
rect 36176 36737 36185 36771
rect 36185 36737 36219 36771
rect 36219 36737 36228 36771
rect 36176 36728 36228 36737
rect 37004 36728 37056 36780
rect 2320 36660 2372 36712
rect 8852 36660 8904 36712
rect 1584 36592 1636 36644
rect 37464 36592 37516 36644
rect 36728 36567 36780 36576
rect 36728 36533 36737 36567
rect 36737 36533 36771 36567
rect 36771 36533 36780 36567
rect 36728 36524 36780 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 11612 36363 11664 36372
rect 11612 36329 11621 36363
rect 11621 36329 11655 36363
rect 11655 36329 11664 36363
rect 11612 36320 11664 36329
rect 29828 36363 29880 36372
rect 29828 36329 29837 36363
rect 29837 36329 29871 36363
rect 29871 36329 29880 36363
rect 29828 36320 29880 36329
rect 36176 36320 36228 36372
rect 4068 36159 4120 36168
rect 4068 36125 4077 36159
rect 4077 36125 4111 36159
rect 4111 36125 4120 36159
rect 4068 36116 4120 36125
rect 11796 36159 11848 36168
rect 11796 36125 11805 36159
rect 11805 36125 11839 36159
rect 11839 36125 11848 36159
rect 11796 36116 11848 36125
rect 29736 36159 29788 36168
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 29736 36116 29788 36125
rect 34796 36116 34848 36168
rect 38016 36116 38068 36168
rect 37280 35980 37332 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 25504 35776 25556 35828
rect 21916 35640 21968 35692
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 8300 35275 8352 35284
rect 8300 35241 8309 35275
rect 8309 35241 8343 35275
rect 8343 35241 8352 35275
rect 8300 35232 8352 35241
rect 16856 35232 16908 35284
rect 8208 35071 8260 35080
rect 8208 35037 8217 35071
rect 8217 35037 8251 35071
rect 8251 35037 8260 35071
rect 8208 35028 8260 35037
rect 14832 35028 14884 35080
rect 35348 35028 35400 35080
rect 38200 34935 38252 34944
rect 38200 34901 38209 34935
rect 38209 34901 38243 34935
rect 38243 34901 38252 34935
rect 38200 34892 38252 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 6552 34688 6604 34740
rect 7840 34688 7892 34740
rect 14648 34731 14700 34740
rect 14648 34697 14657 34731
rect 14657 34697 14691 34731
rect 14691 34697 14700 34731
rect 14648 34688 14700 34697
rect 15568 34688 15620 34740
rect 18512 34688 18564 34740
rect 20628 34688 20680 34740
rect 27896 34688 27948 34740
rect 5816 34552 5868 34604
rect 6552 34552 6604 34604
rect 14740 34552 14792 34604
rect 15016 34552 15068 34604
rect 17868 34595 17920 34604
rect 17868 34561 17877 34595
rect 17877 34561 17911 34595
rect 17911 34561 17920 34595
rect 17868 34552 17920 34561
rect 17500 34484 17552 34536
rect 27252 34552 27304 34604
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 14556 34076 14608 34128
rect 4620 33940 4672 33992
rect 14280 33983 14332 33992
rect 14280 33949 14289 33983
rect 14289 33949 14323 33983
rect 14323 33949 14332 33983
rect 14280 33940 14332 33949
rect 15844 33940 15896 33992
rect 23020 33983 23072 33992
rect 23020 33949 23029 33983
rect 23029 33949 23063 33983
rect 23063 33949 23072 33983
rect 23020 33940 23072 33949
rect 25044 33983 25096 33992
rect 25044 33949 25053 33983
rect 25053 33949 25087 33983
rect 25087 33949 25096 33983
rect 25044 33940 25096 33949
rect 28080 33940 28132 33992
rect 11888 33804 11940 33856
rect 15108 33804 15160 33856
rect 20168 33804 20220 33856
rect 25136 33847 25188 33856
rect 25136 33813 25145 33847
rect 25145 33813 25179 33847
rect 25179 33813 25188 33847
rect 25136 33804 25188 33813
rect 28080 33847 28132 33856
rect 28080 33813 28089 33847
rect 28089 33813 28123 33847
rect 28123 33813 28132 33847
rect 28080 33804 28132 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 1768 33507 1820 33516
rect 1768 33473 1777 33507
rect 1777 33473 1811 33507
rect 1811 33473 1820 33507
rect 1768 33464 1820 33473
rect 38292 33507 38344 33516
rect 38292 33473 38301 33507
rect 38301 33473 38335 33507
rect 38335 33473 38344 33507
rect 38292 33464 38344 33473
rect 3884 33260 3936 33312
rect 38108 33303 38160 33312
rect 38108 33269 38117 33303
rect 38117 33269 38151 33303
rect 38151 33269 38160 33303
rect 38108 33260 38160 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 31760 33056 31812 33108
rect 5632 32895 5684 32904
rect 5632 32861 5641 32895
rect 5641 32861 5675 32895
rect 5675 32861 5684 32895
rect 5632 32852 5684 32861
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 27528 32852 27580 32861
rect 5724 32759 5776 32768
rect 5724 32725 5733 32759
rect 5733 32725 5767 32759
rect 5767 32725 5776 32759
rect 5724 32716 5776 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 1768 32419 1820 32428
rect 1768 32385 1777 32419
rect 1777 32385 1811 32419
rect 1811 32385 1820 32419
rect 1768 32376 1820 32385
rect 35440 32376 35492 32428
rect 3976 32172 4028 32224
rect 38200 32215 38252 32224
rect 38200 32181 38209 32215
rect 38209 32181 38243 32215
rect 38243 32181 38252 32215
rect 38200 32172 38252 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6552 32011 6604 32020
rect 6552 31977 6561 32011
rect 6561 31977 6595 32011
rect 6595 31977 6604 32011
rect 6552 31968 6604 31977
rect 11796 31968 11848 32020
rect 16304 31832 16356 31884
rect 7380 31764 7432 31816
rect 12900 31764 12952 31816
rect 20904 31807 20956 31816
rect 20904 31773 20913 31807
rect 20913 31773 20947 31807
rect 20947 31773 20956 31807
rect 20904 31764 20956 31773
rect 34428 31832 34480 31884
rect 33692 31807 33744 31816
rect 33692 31773 33701 31807
rect 33701 31773 33735 31807
rect 33735 31773 33744 31807
rect 33692 31764 33744 31773
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 13820 31331 13872 31340
rect 13820 31297 13829 31331
rect 13829 31297 13863 31331
rect 13863 31297 13872 31331
rect 13820 31288 13872 31297
rect 30656 31288 30708 31340
rect 11520 31084 11572 31136
rect 16212 31084 16264 31136
rect 24584 31084 24636 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 35348 30880 35400 30932
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 1768 30676 1820 30685
rect 37280 30744 37332 30796
rect 29920 30676 29972 30728
rect 30012 30608 30064 30660
rect 1492 30540 1544 30592
rect 24952 30583 25004 30592
rect 24952 30549 24961 30583
rect 24961 30549 24995 30583
rect 24995 30549 25004 30583
rect 24952 30540 25004 30549
rect 29828 30583 29880 30592
rect 29828 30549 29837 30583
rect 29837 30549 29871 30583
rect 29871 30549 29880 30583
rect 29828 30540 29880 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 8852 30243 8904 30252
rect 8852 30209 8861 30243
rect 8861 30209 8895 30243
rect 8895 30209 8904 30243
rect 8852 30200 8904 30209
rect 36728 30268 36780 30320
rect 33600 30200 33652 30252
rect 12440 29996 12492 30048
rect 30012 30039 30064 30048
rect 30012 30005 30021 30039
rect 30021 30005 30055 30039
rect 30055 30005 30064 30039
rect 30012 29996 30064 30005
rect 38200 30039 38252 30048
rect 38200 30005 38209 30039
rect 38209 30005 38243 30039
rect 38243 30005 38252 30039
rect 38200 29996 38252 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 17868 29792 17920 29844
rect 35440 29792 35492 29844
rect 3884 29588 3936 29640
rect 14740 29631 14792 29640
rect 14740 29597 14749 29631
rect 14749 29597 14783 29631
rect 14783 29597 14792 29631
rect 14740 29588 14792 29597
rect 15844 29588 15896 29640
rect 33784 29588 33836 29640
rect 8116 29452 8168 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 15016 29248 15068 29300
rect 17500 29291 17552 29300
rect 17500 29257 17509 29291
rect 17509 29257 17543 29291
rect 17543 29257 17552 29291
rect 17500 29248 17552 29257
rect 27252 29291 27304 29300
rect 27252 29257 27261 29291
rect 27261 29257 27295 29291
rect 27295 29257 27304 29291
rect 27252 29248 27304 29257
rect 1768 29155 1820 29164
rect 1768 29121 1777 29155
rect 1777 29121 1811 29155
rect 1811 29121 1820 29155
rect 1768 29112 1820 29121
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 15660 29112 15712 29164
rect 24492 29112 24544 29164
rect 38292 29155 38344 29164
rect 38292 29121 38301 29155
rect 38301 29121 38335 29155
rect 38335 29121 38344 29155
rect 38292 29112 38344 29121
rect 6552 28976 6604 29028
rect 33324 28976 33376 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 5816 28704 5868 28756
rect 14832 28704 14884 28756
rect 33784 28704 33836 28756
rect 6184 28500 6236 28552
rect 18328 28500 18380 28552
rect 32772 28543 32824 28552
rect 32772 28509 32781 28543
rect 32781 28509 32815 28543
rect 32815 28509 32824 28543
rect 32772 28500 32824 28509
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3976 28024 4028 28076
rect 38108 28024 38160 28076
rect 4804 27820 4856 27872
rect 30472 27863 30524 27872
rect 30472 27829 30481 27863
rect 30481 27829 30515 27863
rect 30515 27829 30524 27863
rect 30472 27820 30524 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 20628 27412 20680 27464
rect 36728 27412 36780 27464
rect 5724 27276 5776 27328
rect 20904 27276 20956 27328
rect 38200 27319 38252 27328
rect 38200 27285 38209 27319
rect 38209 27285 38243 27319
rect 38243 27285 38252 27319
rect 38200 27276 38252 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 29920 27072 29972 27124
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 20904 26979 20956 26988
rect 20904 26945 20913 26979
rect 20913 26945 20947 26979
rect 20947 26945 20956 26979
rect 20904 26936 20956 26945
rect 24216 26936 24268 26988
rect 8852 26732 8904 26784
rect 20536 26732 20588 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 14464 26460 14516 26512
rect 17224 26460 17276 26512
rect 11796 26324 11848 26376
rect 12532 26324 12584 26376
rect 15292 26324 15344 26376
rect 16856 26256 16908 26308
rect 20628 26324 20680 26376
rect 20444 26256 20496 26308
rect 11980 26188 12032 26240
rect 17684 26188 17736 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 33600 26027 33652 26036
rect 33600 25993 33609 26027
rect 33609 25993 33643 26027
rect 33643 25993 33652 26027
rect 33600 25984 33652 25993
rect 36728 26027 36780 26036
rect 36728 25993 36737 26027
rect 36737 25993 36771 26027
rect 36771 25993 36780 26027
rect 36728 25984 36780 25993
rect 12532 25916 12584 25968
rect 5448 25848 5500 25900
rect 11796 25848 11848 25900
rect 11980 25891 12032 25900
rect 11980 25857 11989 25891
rect 11989 25857 12023 25891
rect 12023 25857 12032 25891
rect 11980 25848 12032 25857
rect 12624 25891 12676 25900
rect 12624 25857 12633 25891
rect 12633 25857 12667 25891
rect 12667 25857 12676 25891
rect 12624 25848 12676 25857
rect 15292 25891 15344 25900
rect 15292 25857 15301 25891
rect 15301 25857 15335 25891
rect 15335 25857 15344 25891
rect 15292 25848 15344 25857
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 17684 25891 17736 25900
rect 17684 25857 17693 25891
rect 17693 25857 17727 25891
rect 17727 25857 17736 25891
rect 17684 25848 17736 25857
rect 23480 25848 23532 25900
rect 31760 25848 31812 25900
rect 36912 25891 36964 25900
rect 36912 25857 36921 25891
rect 36921 25857 36955 25891
rect 36955 25857 36964 25891
rect 36912 25848 36964 25857
rect 13544 25823 13596 25832
rect 13544 25789 13553 25823
rect 13553 25789 13587 25823
rect 13587 25789 13596 25823
rect 13544 25780 13596 25789
rect 15936 25823 15988 25832
rect 15936 25789 15945 25823
rect 15945 25789 15979 25823
rect 15979 25789 15988 25823
rect 15936 25780 15988 25789
rect 10600 25644 10652 25696
rect 11796 25687 11848 25696
rect 11796 25653 11805 25687
rect 11805 25653 11839 25687
rect 11839 25653 11848 25687
rect 11796 25644 11848 25653
rect 14004 25644 14056 25696
rect 14280 25687 14332 25696
rect 14280 25653 14289 25687
rect 14289 25653 14323 25687
rect 14323 25653 14332 25687
rect 14280 25644 14332 25653
rect 15200 25644 15252 25696
rect 16948 25687 17000 25696
rect 16948 25653 16957 25687
rect 16957 25653 16991 25687
rect 16991 25653 17000 25687
rect 16948 25644 17000 25653
rect 17500 25687 17552 25696
rect 17500 25653 17509 25687
rect 17509 25653 17543 25687
rect 17543 25653 17552 25687
rect 17500 25644 17552 25653
rect 23572 25644 23624 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 12624 25440 12676 25492
rect 14740 25483 14792 25492
rect 14740 25449 14749 25483
rect 14749 25449 14783 25483
rect 14783 25449 14792 25483
rect 14740 25440 14792 25449
rect 5816 25372 5868 25424
rect 13360 25372 13412 25424
rect 8116 25304 8168 25356
rect 10600 25347 10652 25356
rect 10600 25313 10609 25347
rect 10609 25313 10643 25347
rect 10643 25313 10652 25347
rect 10600 25304 10652 25313
rect 11796 25304 11848 25356
rect 13544 25304 13596 25356
rect 14464 25347 14516 25356
rect 14464 25313 14473 25347
rect 14473 25313 14507 25347
rect 14507 25313 14516 25347
rect 14464 25304 14516 25313
rect 15936 25347 15988 25356
rect 15936 25313 15945 25347
rect 15945 25313 15979 25347
rect 15979 25313 15988 25347
rect 15936 25304 15988 25313
rect 17500 25304 17552 25356
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 7196 25236 7248 25288
rect 9864 25236 9916 25288
rect 11520 25236 11572 25288
rect 14188 25236 14240 25288
rect 17224 25279 17276 25288
rect 17224 25245 17233 25279
rect 17233 25245 17267 25279
rect 17267 25245 17276 25279
rect 17224 25236 17276 25245
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 38292 25279 38344 25288
rect 38292 25245 38301 25279
rect 38301 25245 38335 25279
rect 38335 25245 38344 25279
rect 38292 25236 38344 25245
rect 5172 25100 5224 25152
rect 13360 25100 13412 25152
rect 16580 25143 16632 25152
rect 16580 25109 16589 25143
rect 16589 25109 16623 25143
rect 16623 25109 16632 25143
rect 16580 25100 16632 25109
rect 17040 25143 17092 25152
rect 17040 25109 17049 25143
rect 17049 25109 17083 25143
rect 17083 25109 17092 25143
rect 17040 25100 17092 25109
rect 20352 25143 20404 25152
rect 20352 25109 20361 25143
rect 20361 25109 20395 25143
rect 20395 25109 20404 25143
rect 20352 25100 20404 25109
rect 23388 25143 23440 25152
rect 23388 25109 23397 25143
rect 23397 25109 23431 25143
rect 23431 25109 23440 25143
rect 23388 25100 23440 25109
rect 33968 25100 34020 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14740 24896 14792 24948
rect 15200 24871 15252 24880
rect 15200 24837 15209 24871
rect 15209 24837 15243 24871
rect 15243 24837 15252 24871
rect 15200 24828 15252 24837
rect 17040 24871 17092 24880
rect 17040 24837 17049 24871
rect 17049 24837 17083 24871
rect 17083 24837 17092 24871
rect 17040 24828 17092 24837
rect 5172 24803 5224 24812
rect 5172 24769 5181 24803
rect 5181 24769 5215 24803
rect 5215 24769 5224 24803
rect 5172 24760 5224 24769
rect 7288 24803 7340 24812
rect 7288 24769 7297 24803
rect 7297 24769 7331 24803
rect 7331 24769 7340 24803
rect 7288 24760 7340 24769
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 9864 24760 9916 24812
rect 11244 24760 11296 24812
rect 12348 24760 12400 24812
rect 13360 24760 13412 24812
rect 13728 24735 13780 24744
rect 13728 24701 13737 24735
rect 13737 24701 13771 24735
rect 13771 24701 13780 24735
rect 13728 24692 13780 24701
rect 14280 24760 14332 24812
rect 20352 24803 20404 24812
rect 20352 24769 20361 24803
rect 20361 24769 20395 24803
rect 20395 24769 20404 24803
rect 20352 24760 20404 24769
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 22008 24760 22060 24812
rect 22560 24760 22612 24812
rect 23480 24760 23532 24812
rect 33324 24803 33376 24812
rect 33324 24769 33333 24803
rect 33333 24769 33367 24803
rect 33367 24769 33376 24803
rect 33324 24760 33376 24769
rect 35532 24803 35584 24812
rect 35532 24769 35541 24803
rect 35541 24769 35575 24803
rect 35575 24769 35584 24803
rect 35532 24760 35584 24769
rect 36912 24760 36964 24812
rect 16580 24692 16632 24744
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 4988 24599 5040 24608
rect 4988 24565 4997 24599
rect 4997 24565 5031 24599
rect 5031 24565 5040 24599
rect 4988 24556 5040 24565
rect 7564 24556 7616 24608
rect 11796 24599 11848 24608
rect 11796 24565 11805 24599
rect 11805 24565 11839 24599
rect 11839 24565 11848 24599
rect 11796 24556 11848 24565
rect 32772 24624 32824 24676
rect 13176 24556 13228 24608
rect 20812 24599 20864 24608
rect 20812 24565 20821 24599
rect 20821 24565 20855 24599
rect 20855 24565 20864 24599
rect 20812 24556 20864 24565
rect 21456 24556 21508 24608
rect 22744 24556 22796 24608
rect 33416 24599 33468 24608
rect 33416 24565 33425 24599
rect 33425 24565 33459 24599
rect 33459 24565 33468 24599
rect 33416 24556 33468 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 13728 24352 13780 24404
rect 16580 24395 16632 24404
rect 16580 24361 16589 24395
rect 16589 24361 16623 24395
rect 16623 24361 16632 24395
rect 16580 24352 16632 24361
rect 20812 24395 20864 24404
rect 20812 24361 20821 24395
rect 20821 24361 20855 24395
rect 20855 24361 20864 24395
rect 20812 24352 20864 24361
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 2320 24191 2372 24200
rect 2320 24157 2329 24191
rect 2329 24157 2363 24191
rect 2363 24157 2372 24191
rect 2320 24148 2372 24157
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 7564 24191 7616 24200
rect 7564 24157 7573 24191
rect 7573 24157 7607 24191
rect 7607 24157 7616 24191
rect 7564 24148 7616 24157
rect 12624 24216 12676 24268
rect 14004 24216 14056 24268
rect 16212 24259 16264 24268
rect 16212 24225 16221 24259
rect 16221 24225 16255 24259
rect 16255 24225 16264 24259
rect 16212 24216 16264 24225
rect 16948 24216 17000 24268
rect 20168 24259 20220 24268
rect 20168 24225 20177 24259
rect 20177 24225 20211 24259
rect 20211 24225 20220 24259
rect 20168 24216 20220 24225
rect 20444 24216 20496 24268
rect 21640 24284 21692 24336
rect 21916 24327 21968 24336
rect 21916 24293 21925 24327
rect 21925 24293 21959 24327
rect 21959 24293 21968 24327
rect 21916 24284 21968 24293
rect 22744 24259 22796 24268
rect 22744 24225 22753 24259
rect 22753 24225 22787 24259
rect 22787 24225 22796 24259
rect 22744 24216 22796 24225
rect 11796 24148 11848 24200
rect 11520 24080 11572 24132
rect 12348 24080 12400 24132
rect 13084 24148 13136 24200
rect 17960 24148 18012 24200
rect 24768 24191 24820 24200
rect 17868 24080 17920 24132
rect 21456 24123 21508 24132
rect 21456 24089 21465 24123
rect 21465 24089 21499 24123
rect 21499 24089 21508 24123
rect 24768 24157 24777 24191
rect 24777 24157 24811 24191
rect 24811 24157 24820 24191
rect 24768 24148 24820 24157
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 21456 24080 21508 24089
rect 33692 24080 33744 24132
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 1952 24012 2004 24064
rect 5080 24012 5132 24064
rect 6736 24055 6788 24064
rect 6736 24021 6745 24055
rect 6745 24021 6779 24055
rect 6779 24021 6788 24055
rect 6736 24012 6788 24021
rect 6920 24012 6972 24064
rect 12072 24012 12124 24064
rect 12808 24012 12860 24064
rect 12992 24055 13044 24064
rect 12992 24021 13001 24055
rect 13001 24021 13035 24055
rect 13035 24021 13044 24055
rect 12992 24012 13044 24021
rect 14464 24012 14516 24064
rect 23204 24055 23256 24064
rect 23204 24021 23213 24055
rect 23213 24021 23247 24055
rect 23247 24021 23256 24055
rect 23204 24012 23256 24021
rect 25228 24012 25280 24064
rect 37004 24012 37056 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23808 1636 23860
rect 10876 23808 10928 23860
rect 13084 23808 13136 23860
rect 1952 23715 2004 23724
rect 1952 23681 1961 23715
rect 1961 23681 1995 23715
rect 1995 23681 2004 23715
rect 1952 23672 2004 23681
rect 2136 23672 2188 23724
rect 2688 23672 2740 23724
rect 3884 23715 3936 23724
rect 3884 23681 3893 23715
rect 3893 23681 3927 23715
rect 3927 23681 3936 23715
rect 3884 23672 3936 23681
rect 5356 23715 5408 23724
rect 2596 23604 2648 23656
rect 4160 23604 4212 23656
rect 5356 23681 5365 23715
rect 5365 23681 5399 23715
rect 5399 23681 5408 23715
rect 5356 23672 5408 23681
rect 5724 23672 5776 23724
rect 7196 23672 7248 23724
rect 9404 23715 9456 23724
rect 9404 23681 9413 23715
rect 9413 23681 9447 23715
rect 9447 23681 9456 23715
rect 9404 23672 9456 23681
rect 10968 23672 11020 23724
rect 12624 23672 12676 23724
rect 22008 23851 22060 23860
rect 15844 23783 15896 23792
rect 15844 23749 15853 23783
rect 15853 23749 15887 23783
rect 15887 23749 15896 23783
rect 15844 23740 15896 23749
rect 22008 23817 22017 23851
rect 22017 23817 22051 23851
rect 22051 23817 22060 23851
rect 22008 23808 22060 23817
rect 23204 23808 23256 23860
rect 18420 23715 18472 23724
rect 6828 23604 6880 23656
rect 4896 23536 4948 23588
rect 9588 23536 9640 23588
rect 13084 23604 13136 23656
rect 18420 23681 18429 23715
rect 18429 23681 18463 23715
rect 18463 23681 18472 23715
rect 18420 23672 18472 23681
rect 20076 23672 20128 23724
rect 24768 23740 24820 23792
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22652 23715 22704 23724
rect 22652 23681 22661 23715
rect 22661 23681 22695 23715
rect 22695 23681 22704 23715
rect 22652 23672 22704 23681
rect 23388 23672 23440 23724
rect 25228 23715 25280 23724
rect 24400 23647 24452 23656
rect 24400 23613 24409 23647
rect 24409 23613 24443 23647
rect 24443 23613 24452 23647
rect 24400 23604 24452 23613
rect 25228 23681 25237 23715
rect 25237 23681 25271 23715
rect 25271 23681 25280 23715
rect 25228 23672 25280 23681
rect 25504 23604 25556 23656
rect 2872 23468 2924 23520
rect 3148 23468 3200 23520
rect 4620 23511 4672 23520
rect 4620 23477 4629 23511
rect 4629 23477 4663 23511
rect 4663 23477 4672 23511
rect 4620 23468 4672 23477
rect 6644 23468 6696 23520
rect 8024 23468 8076 23520
rect 9680 23468 9732 23520
rect 12256 23468 12308 23520
rect 14832 23468 14884 23520
rect 17684 23511 17736 23520
rect 17684 23477 17693 23511
rect 17693 23477 17727 23511
rect 17727 23477 17736 23511
rect 17684 23468 17736 23477
rect 18512 23511 18564 23520
rect 18512 23477 18521 23511
rect 18521 23477 18555 23511
rect 18555 23477 18564 23511
rect 18512 23468 18564 23477
rect 18696 23468 18748 23520
rect 20996 23511 21048 23520
rect 20996 23477 21005 23511
rect 21005 23477 21039 23511
rect 21039 23477 21048 23511
rect 20996 23468 21048 23477
rect 23756 23511 23808 23520
rect 23756 23477 23765 23511
rect 23765 23477 23799 23511
rect 23799 23477 23808 23511
rect 23756 23468 23808 23477
rect 25044 23511 25096 23520
rect 25044 23477 25053 23511
rect 25053 23477 25087 23511
rect 25087 23477 25096 23511
rect 25044 23468 25096 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3884 23196 3936 23248
rect 5540 23196 5592 23248
rect 4896 23171 4948 23180
rect 4896 23137 4905 23171
rect 4905 23137 4939 23171
rect 4939 23137 4948 23171
rect 4896 23128 4948 23137
rect 4988 23128 5040 23180
rect 1676 22924 1728 22976
rect 2688 23060 2740 23112
rect 4160 23060 4212 23112
rect 5172 23060 5224 23112
rect 7288 23196 7340 23248
rect 9404 23264 9456 23316
rect 12440 23264 12492 23316
rect 20076 23307 20128 23316
rect 9312 23196 9364 23248
rect 15016 23196 15068 23248
rect 6736 23171 6788 23180
rect 6736 23137 6745 23171
rect 6745 23137 6779 23171
rect 6779 23137 6788 23171
rect 6736 23128 6788 23137
rect 7380 23171 7432 23180
rect 7380 23137 7389 23171
rect 7389 23137 7423 23171
rect 7423 23137 7432 23171
rect 7380 23128 7432 23137
rect 9680 23171 9732 23180
rect 9680 23137 9689 23171
rect 9689 23137 9723 23171
rect 9723 23137 9732 23171
rect 9680 23128 9732 23137
rect 11888 23171 11940 23180
rect 11888 23137 11897 23171
rect 11897 23137 11931 23171
rect 11931 23137 11940 23171
rect 11888 23128 11940 23137
rect 12072 23171 12124 23180
rect 12072 23137 12081 23171
rect 12081 23137 12115 23171
rect 12115 23137 12124 23171
rect 12072 23128 12124 23137
rect 13084 23171 13136 23180
rect 13084 23137 13093 23171
rect 13093 23137 13127 23171
rect 13127 23137 13136 23171
rect 13084 23128 13136 23137
rect 14096 23128 14148 23180
rect 14464 23171 14516 23180
rect 14464 23137 14473 23171
rect 14473 23137 14507 23171
rect 14507 23137 14516 23171
rect 14464 23128 14516 23137
rect 20076 23273 20085 23307
rect 20085 23273 20119 23307
rect 20119 23273 20128 23307
rect 20076 23264 20128 23273
rect 20536 23196 20588 23248
rect 17684 23128 17736 23180
rect 18512 23128 18564 23180
rect 21364 23264 21416 23316
rect 29828 23264 29880 23316
rect 28080 23196 28132 23248
rect 20996 23171 21048 23180
rect 6552 22992 6604 23044
rect 6920 22992 6972 23044
rect 7564 22992 7616 23044
rect 9404 23060 9456 23112
rect 11244 23103 11296 23112
rect 11244 23069 11253 23103
rect 11253 23069 11287 23103
rect 11287 23069 11296 23103
rect 11244 23060 11296 23069
rect 14280 23103 14332 23112
rect 14280 23069 14289 23103
rect 14289 23069 14323 23103
rect 14323 23069 14332 23103
rect 14280 23060 14332 23069
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 23204 23128 23256 23180
rect 24400 23128 24452 23180
rect 25044 23128 25096 23180
rect 20168 23060 20220 23112
rect 20812 23103 20864 23112
rect 2780 22924 2832 22976
rect 3240 22967 3292 22976
rect 3240 22933 3249 22967
rect 3249 22933 3283 22967
rect 3283 22933 3292 22967
rect 3240 22924 3292 22933
rect 6092 22967 6144 22976
rect 6092 22933 6101 22967
rect 6101 22933 6135 22967
rect 6135 22933 6144 22967
rect 6092 22924 6144 22933
rect 9680 22924 9732 22976
rect 10600 22967 10652 22976
rect 10600 22933 10609 22967
rect 10609 22933 10643 22967
rect 10643 22933 10652 22967
rect 10600 22924 10652 22933
rect 12348 22924 12400 22976
rect 13176 23035 13228 23044
rect 13176 23001 13185 23035
rect 13185 23001 13219 23035
rect 13219 23001 13228 23035
rect 13176 22992 13228 23001
rect 16120 22992 16172 23044
rect 18420 22992 18472 23044
rect 20812 23069 20821 23103
rect 20821 23069 20855 23103
rect 20855 23069 20864 23103
rect 20812 23060 20864 23069
rect 23572 23060 23624 23112
rect 33968 23103 34020 23112
rect 33968 23069 33977 23103
rect 33977 23069 34011 23103
rect 34011 23069 34020 23103
rect 33968 23060 34020 23069
rect 20536 22992 20588 23044
rect 22100 22992 22152 23044
rect 22468 23035 22520 23044
rect 22468 23001 22477 23035
rect 22477 23001 22511 23035
rect 22511 23001 22520 23035
rect 22468 22992 22520 23001
rect 22652 22992 22704 23044
rect 34796 22992 34848 23044
rect 15108 22924 15160 22976
rect 16028 22967 16080 22976
rect 16028 22933 16037 22967
rect 16037 22933 16071 22967
rect 16071 22933 16080 22967
rect 16028 22924 16080 22933
rect 18604 22924 18656 22976
rect 19248 22924 19300 22976
rect 20812 22924 20864 22976
rect 21364 22924 21416 22976
rect 23480 22924 23532 22976
rect 25044 22924 25096 22976
rect 34060 22967 34112 22976
rect 34060 22933 34069 22967
rect 34069 22933 34103 22967
rect 34103 22933 34112 22967
rect 34060 22924 34112 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9404 22763 9456 22772
rect 3884 22652 3936 22704
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 4160 22584 4212 22636
rect 5356 22584 5408 22636
rect 6276 22584 6328 22636
rect 9404 22729 9413 22763
rect 9413 22729 9447 22763
rect 9447 22729 9456 22763
rect 9404 22720 9456 22729
rect 8576 22652 8628 22704
rect 15384 22720 15436 22772
rect 18236 22720 18288 22772
rect 18604 22763 18656 22772
rect 18604 22729 18613 22763
rect 18613 22729 18647 22763
rect 18647 22729 18656 22763
rect 18604 22720 18656 22729
rect 20168 22763 20220 22772
rect 20168 22729 20177 22763
rect 20177 22729 20211 22763
rect 20211 22729 20220 22763
rect 20168 22720 20220 22729
rect 25044 22763 25096 22772
rect 10600 22652 10652 22704
rect 12256 22695 12308 22704
rect 12256 22661 12265 22695
rect 12265 22661 12299 22695
rect 12299 22661 12308 22695
rect 12256 22652 12308 22661
rect 12900 22652 12952 22704
rect 13452 22652 13504 22704
rect 15108 22695 15160 22704
rect 15108 22661 15117 22695
rect 15117 22661 15151 22695
rect 15151 22661 15160 22695
rect 15108 22652 15160 22661
rect 15660 22695 15712 22704
rect 15660 22661 15669 22695
rect 15669 22661 15703 22695
rect 15703 22661 15712 22695
rect 15660 22652 15712 22661
rect 25044 22729 25053 22763
rect 25053 22729 25087 22763
rect 25087 22729 25096 22763
rect 25044 22720 25096 22729
rect 25504 22763 25556 22772
rect 25504 22729 25513 22763
rect 25513 22729 25547 22763
rect 25547 22729 25556 22763
rect 25504 22720 25556 22729
rect 23480 22652 23532 22704
rect 7196 22584 7248 22636
rect 7564 22584 7616 22636
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 9588 22584 9640 22636
rect 14556 22584 14608 22636
rect 15936 22584 15988 22636
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 16488 22584 16540 22636
rect 17960 22627 18012 22636
rect 17960 22593 17969 22627
rect 17969 22593 18003 22627
rect 18003 22593 18012 22627
rect 17960 22584 18012 22593
rect 18696 22584 18748 22636
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 20168 22584 20220 22636
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 25228 22584 25280 22636
rect 37004 22584 37056 22636
rect 1584 22516 1636 22568
rect 3516 22516 3568 22568
rect 10232 22559 10284 22568
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 12808 22516 12860 22568
rect 15016 22559 15068 22568
rect 15016 22525 15025 22559
rect 15025 22525 15059 22559
rect 15059 22525 15068 22559
rect 15016 22516 15068 22525
rect 19064 22559 19116 22568
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 22100 22559 22152 22568
rect 22100 22525 22109 22559
rect 22109 22525 22143 22559
rect 22143 22525 22152 22559
rect 22100 22516 22152 22525
rect 24400 22559 24452 22568
rect 24400 22525 24409 22559
rect 24409 22525 24443 22559
rect 24443 22525 24452 22559
rect 24400 22516 24452 22525
rect 25412 22516 25464 22568
rect 9220 22448 9272 22500
rect 29736 22448 29788 22500
rect 4712 22380 4764 22432
rect 4988 22423 5040 22432
rect 4988 22389 4997 22423
rect 4997 22389 5031 22423
rect 5031 22389 5040 22423
rect 4988 22380 5040 22389
rect 6000 22380 6052 22432
rect 6368 22380 6420 22432
rect 6920 22380 6972 22432
rect 13912 22380 13964 22432
rect 14004 22380 14056 22432
rect 16212 22423 16264 22432
rect 16212 22389 16221 22423
rect 16221 22389 16255 22423
rect 16255 22389 16264 22423
rect 16212 22380 16264 22389
rect 16856 22423 16908 22432
rect 16856 22389 16865 22423
rect 16865 22389 16899 22423
rect 16899 22389 16908 22423
rect 16856 22380 16908 22389
rect 19432 22423 19484 22432
rect 19432 22389 19441 22423
rect 19441 22389 19475 22423
rect 19475 22389 19484 22423
rect 19432 22380 19484 22389
rect 19524 22380 19576 22432
rect 24952 22380 25004 22432
rect 32404 22423 32456 22432
rect 32404 22389 32413 22423
rect 32413 22389 32447 22423
rect 32447 22389 32456 22423
rect 32404 22380 32456 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6644 22176 6696 22228
rect 10232 22176 10284 22228
rect 11152 22176 11204 22228
rect 6828 22108 6880 22160
rect 1584 21972 1636 22024
rect 5632 22040 5684 22092
rect 5908 22083 5960 22092
rect 5908 22049 5917 22083
rect 5917 22049 5951 22083
rect 5951 22049 5960 22083
rect 5908 22040 5960 22049
rect 6736 21972 6788 22024
rect 7012 21972 7064 22024
rect 7656 21972 7708 22024
rect 7840 22015 7892 22024
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 2964 21904 3016 21956
rect 4436 21947 4488 21956
rect 4436 21913 4445 21947
rect 4445 21913 4479 21947
rect 4479 21913 4488 21947
rect 4436 21904 4488 21913
rect 8024 22083 8076 22092
rect 8024 22049 8033 22083
rect 8033 22049 8067 22083
rect 8067 22049 8076 22083
rect 8024 22040 8076 22049
rect 8116 21972 8168 22024
rect 8484 22040 8536 22092
rect 10968 22040 11020 22092
rect 8392 21972 8444 22024
rect 9956 21972 10008 22024
rect 2688 21836 2740 21888
rect 6184 21879 6236 21888
rect 6184 21845 6193 21879
rect 6193 21845 6227 21879
rect 6227 21845 6236 21879
rect 6184 21836 6236 21845
rect 7104 21836 7156 21888
rect 10508 21904 10560 21956
rect 11336 21904 11388 21956
rect 12348 22108 12400 22160
rect 14280 22176 14332 22228
rect 23296 22176 23348 22228
rect 24400 22176 24452 22228
rect 33784 22176 33836 22228
rect 12440 21836 12492 21888
rect 12900 21972 12952 22024
rect 14556 21972 14608 22024
rect 15752 21972 15804 22024
rect 16856 22040 16908 22092
rect 16488 22015 16540 22024
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 19340 22108 19392 22160
rect 19064 22040 19116 22092
rect 19524 22040 19576 22092
rect 21272 22040 21324 22092
rect 23112 22040 23164 22092
rect 23756 22040 23808 22092
rect 25412 22040 25464 22092
rect 13912 21904 13964 21956
rect 14832 21947 14884 21956
rect 14832 21913 14841 21947
rect 14841 21913 14875 21947
rect 14875 21913 14884 21947
rect 14832 21904 14884 21913
rect 12808 21836 12860 21888
rect 14004 21836 14056 21888
rect 15844 21879 15896 21888
rect 15844 21845 15853 21879
rect 15853 21845 15887 21879
rect 15887 21845 15896 21879
rect 15844 21836 15896 21845
rect 16672 21836 16724 21888
rect 17684 21947 17736 21956
rect 17684 21913 17693 21947
rect 17693 21913 17727 21947
rect 17727 21913 17736 21947
rect 17684 21904 17736 21913
rect 18328 21904 18380 21956
rect 20720 22015 20772 22024
rect 20720 21981 20729 22015
rect 20729 21981 20763 22015
rect 20763 21981 20772 22015
rect 20720 21972 20772 21981
rect 20628 21904 20680 21956
rect 22008 21972 22060 22024
rect 22192 21904 22244 21956
rect 24492 21972 24544 22024
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 24860 21972 24912 22024
rect 38292 22015 38344 22024
rect 19432 21836 19484 21888
rect 20536 21879 20588 21888
rect 20536 21845 20545 21879
rect 20545 21845 20579 21879
rect 20579 21845 20588 21879
rect 20536 21836 20588 21845
rect 20904 21836 20956 21888
rect 22468 21836 22520 21888
rect 23112 21836 23164 21888
rect 23664 21904 23716 21956
rect 31852 21947 31904 21956
rect 31852 21913 31861 21947
rect 31861 21913 31895 21947
rect 31895 21913 31904 21947
rect 31852 21904 31904 21913
rect 25136 21836 25188 21888
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1308 21632 1360 21684
rect 2688 21607 2740 21616
rect 2688 21573 2697 21607
rect 2697 21573 2731 21607
rect 2731 21573 2740 21607
rect 2688 21564 2740 21573
rect 3700 21632 3752 21684
rect 5356 21632 5408 21684
rect 6184 21632 6236 21684
rect 7748 21632 7800 21684
rect 7840 21632 7892 21684
rect 8760 21607 8812 21616
rect 8760 21573 8769 21607
rect 8769 21573 8803 21607
rect 8803 21573 8812 21607
rect 8760 21564 8812 21573
rect 10416 21564 10468 21616
rect 12440 21564 12492 21616
rect 12992 21564 13044 21616
rect 14096 21607 14148 21616
rect 14096 21573 14105 21607
rect 14105 21573 14139 21607
rect 14139 21573 14148 21607
rect 14096 21564 14148 21573
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 5080 21539 5132 21548
rect 5080 21505 5089 21539
rect 5089 21505 5123 21539
rect 5123 21505 5132 21539
rect 5080 21496 5132 21505
rect 5724 21496 5776 21548
rect 6920 21496 6972 21548
rect 8116 21496 8168 21548
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 12624 21496 12676 21548
rect 14648 21632 14700 21684
rect 15016 21564 15068 21616
rect 17224 21607 17276 21616
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 15844 21496 15896 21505
rect 1584 21428 1636 21480
rect 4436 21471 4488 21480
rect 4436 21437 4445 21471
rect 4445 21437 4479 21471
rect 4479 21437 4488 21471
rect 4436 21428 4488 21437
rect 4896 21428 4948 21480
rect 4620 21360 4672 21412
rect 1952 21292 2004 21344
rect 3056 21292 3108 21344
rect 6368 21292 6420 21344
rect 6736 21360 6788 21412
rect 7840 21292 7892 21344
rect 8760 21428 8812 21480
rect 9772 21428 9824 21480
rect 10508 21428 10560 21480
rect 12900 21360 12952 21412
rect 14188 21428 14240 21480
rect 14740 21471 14792 21480
rect 14740 21437 14749 21471
rect 14749 21437 14783 21471
rect 14783 21437 14792 21471
rect 14740 21428 14792 21437
rect 15752 21428 15804 21480
rect 17224 21573 17233 21607
rect 17233 21573 17267 21607
rect 17267 21573 17276 21607
rect 17224 21564 17276 21573
rect 17684 21632 17736 21684
rect 22008 21675 22060 21684
rect 20536 21564 20588 21616
rect 20904 21607 20956 21616
rect 20904 21573 20913 21607
rect 20913 21573 20947 21607
rect 20947 21573 20956 21607
rect 20904 21564 20956 21573
rect 21640 21564 21692 21616
rect 22008 21641 22017 21675
rect 22017 21641 22051 21675
rect 22051 21641 22060 21675
rect 22008 21632 22060 21641
rect 23480 21632 23532 21684
rect 33784 21675 33836 21684
rect 33784 21641 33793 21675
rect 33793 21641 33827 21675
rect 33827 21641 33836 21675
rect 33784 21632 33836 21641
rect 24216 21607 24268 21616
rect 24216 21573 24225 21607
rect 24225 21573 24259 21607
rect 24259 21573 24268 21607
rect 24216 21564 24268 21573
rect 24492 21564 24544 21616
rect 19340 21496 19392 21548
rect 19984 21496 20036 21548
rect 20444 21496 20496 21548
rect 22100 21496 22152 21548
rect 20628 21428 20680 21480
rect 20904 21428 20956 21480
rect 21272 21428 21324 21480
rect 24584 21496 24636 21548
rect 25228 21496 25280 21548
rect 25504 21539 25556 21548
rect 25504 21505 25513 21539
rect 25513 21505 25547 21539
rect 25547 21505 25556 21539
rect 25504 21496 25556 21505
rect 23664 21428 23716 21480
rect 24860 21428 24912 21480
rect 38108 21496 38160 21548
rect 18144 21360 18196 21412
rect 19432 21360 19484 21412
rect 9772 21292 9824 21344
rect 9956 21292 10008 21344
rect 10508 21292 10560 21344
rect 14556 21292 14608 21344
rect 14832 21292 14884 21344
rect 15200 21292 15252 21344
rect 16396 21292 16448 21344
rect 20444 21292 20496 21344
rect 20536 21292 20588 21344
rect 25596 21292 25648 21344
rect 25964 21335 26016 21344
rect 25964 21301 25973 21335
rect 25973 21301 26007 21335
rect 26007 21301 26016 21335
rect 25964 21292 26016 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5908 21088 5960 21140
rect 4252 20952 4304 21004
rect 9864 21088 9916 21140
rect 10324 21088 10376 21140
rect 16396 21088 16448 21140
rect 16764 21088 16816 21140
rect 20536 21088 20588 21140
rect 25504 21088 25556 21140
rect 25596 21088 25648 21140
rect 8484 21020 8536 21072
rect 9312 21020 9364 21072
rect 14832 21063 14884 21072
rect 14832 21029 14841 21063
rect 14841 21029 14875 21063
rect 14875 21029 14884 21063
rect 14832 21020 14884 21029
rect 15108 21020 15160 21072
rect 19984 21020 20036 21072
rect 7196 20952 7248 21004
rect 8116 20952 8168 21004
rect 9956 20952 10008 21004
rect 10232 20995 10284 21004
rect 10232 20961 10241 20995
rect 10241 20961 10275 20995
rect 10275 20961 10284 20995
rect 10508 20995 10560 21004
rect 10232 20952 10284 20961
rect 10508 20961 10517 20995
rect 10517 20961 10551 20995
rect 10551 20961 10560 20995
rect 10508 20952 10560 20961
rect 10600 20952 10652 21004
rect 1584 20927 1636 20936
rect 1584 20893 1593 20927
rect 1593 20893 1627 20927
rect 1627 20893 1636 20927
rect 1584 20884 1636 20893
rect 6736 20884 6788 20936
rect 8484 20884 8536 20936
rect 2872 20816 2924 20868
rect 3608 20816 3660 20868
rect 5264 20816 5316 20868
rect 7564 20816 7616 20868
rect 10048 20884 10100 20936
rect 4160 20748 4212 20800
rect 4896 20748 4948 20800
rect 10600 20816 10652 20868
rect 11060 20816 11112 20868
rect 11796 20748 11848 20800
rect 13268 20952 13320 21004
rect 13452 20995 13504 21004
rect 13452 20961 13461 20995
rect 13461 20961 13495 20995
rect 13495 20961 13504 20995
rect 13452 20952 13504 20961
rect 14924 20952 14976 21004
rect 16672 20952 16724 21004
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 15936 20884 15988 20936
rect 16304 20927 16356 20936
rect 16304 20893 16313 20927
rect 16313 20893 16347 20927
rect 16347 20893 16356 20927
rect 16304 20884 16356 20893
rect 12900 20859 12952 20868
rect 12900 20825 12909 20859
rect 12909 20825 12943 20859
rect 12943 20825 12952 20859
rect 19340 20952 19392 21004
rect 20076 20952 20128 21004
rect 20444 20995 20496 21004
rect 20444 20961 20453 20995
rect 20453 20961 20487 20995
rect 20487 20961 20496 20995
rect 20444 20952 20496 20961
rect 25964 21020 26016 21072
rect 31760 21088 31812 21140
rect 38108 21131 38160 21140
rect 38108 21097 38117 21131
rect 38117 21097 38151 21131
rect 38151 21097 38160 21131
rect 38108 21088 38160 21097
rect 30472 21020 30524 21072
rect 18512 20884 18564 20936
rect 20812 20884 20864 20936
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 22284 20927 22336 20936
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 22744 20884 22796 20936
rect 24676 20884 24728 20936
rect 25780 20884 25832 20936
rect 25872 20927 25924 20936
rect 25872 20893 25881 20927
rect 25881 20893 25915 20927
rect 25915 20893 25924 20927
rect 25872 20884 25924 20893
rect 27804 20927 27856 20936
rect 27804 20893 27813 20927
rect 27813 20893 27847 20927
rect 27847 20893 27856 20927
rect 27804 20884 27856 20893
rect 38292 20927 38344 20936
rect 38292 20893 38301 20927
rect 38301 20893 38335 20927
rect 38335 20893 38344 20927
rect 38292 20884 38344 20893
rect 17684 20859 17736 20868
rect 12900 20816 12952 20825
rect 17684 20825 17693 20859
rect 17693 20825 17727 20859
rect 17727 20825 17736 20859
rect 17684 20816 17736 20825
rect 18052 20816 18104 20868
rect 18144 20816 18196 20868
rect 15292 20748 15344 20800
rect 15752 20748 15804 20800
rect 16764 20748 16816 20800
rect 35532 20816 35584 20868
rect 19432 20791 19484 20800
rect 19432 20757 19441 20791
rect 19441 20757 19475 20791
rect 19475 20757 19484 20791
rect 19432 20748 19484 20757
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 21364 20791 21416 20800
rect 21364 20757 21373 20791
rect 21373 20757 21407 20791
rect 21407 20757 21416 20791
rect 21364 20748 21416 20757
rect 22468 20748 22520 20800
rect 24032 20791 24084 20800
rect 24032 20757 24041 20791
rect 24041 20757 24075 20791
rect 24075 20757 24084 20791
rect 24032 20748 24084 20757
rect 25412 20791 25464 20800
rect 25412 20757 25421 20791
rect 25421 20757 25455 20791
rect 25455 20757 25464 20791
rect 25412 20748 25464 20757
rect 25964 20791 26016 20800
rect 25964 20757 25973 20791
rect 25973 20757 26007 20791
rect 26007 20757 26016 20791
rect 25964 20748 26016 20757
rect 26516 20791 26568 20800
rect 26516 20757 26525 20791
rect 26525 20757 26559 20791
rect 26559 20757 26568 20791
rect 26516 20748 26568 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 11152 20587 11204 20596
rect 3240 20476 3292 20528
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 4528 20519 4580 20528
rect 4528 20485 4537 20519
rect 4537 20485 4571 20519
rect 4571 20485 4580 20519
rect 4528 20476 4580 20485
rect 5540 20476 5592 20528
rect 7564 20476 7616 20528
rect 4252 20451 4304 20460
rect 3608 20408 3660 20417
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 9772 20476 9824 20528
rect 11152 20553 11161 20587
rect 11161 20553 11195 20587
rect 11195 20553 11204 20587
rect 11152 20544 11204 20553
rect 11336 20544 11388 20596
rect 11704 20544 11756 20596
rect 12532 20544 12584 20596
rect 10784 20408 10836 20460
rect 5908 20340 5960 20392
rect 6736 20383 6788 20392
rect 6736 20349 6745 20383
rect 6745 20349 6779 20383
rect 6779 20349 6788 20383
rect 6736 20340 6788 20349
rect 7564 20340 7616 20392
rect 8576 20340 8628 20392
rect 9128 20340 9180 20392
rect 10048 20340 10100 20392
rect 12624 20476 12676 20528
rect 14648 20476 14700 20528
rect 13544 20408 13596 20460
rect 15292 20476 15344 20528
rect 17684 20544 17736 20596
rect 18052 20544 18104 20596
rect 22284 20544 22336 20596
rect 24860 20544 24912 20596
rect 25412 20587 25464 20596
rect 25412 20553 25421 20587
rect 25421 20553 25455 20587
rect 25455 20553 25464 20587
rect 25412 20544 25464 20553
rect 25780 20544 25832 20596
rect 18144 20476 18196 20528
rect 18328 20519 18380 20528
rect 18328 20485 18337 20519
rect 18337 20485 18371 20519
rect 18371 20485 18380 20519
rect 18328 20476 18380 20485
rect 20076 20476 20128 20528
rect 14372 20340 14424 20392
rect 4252 20204 4304 20256
rect 5080 20204 5132 20256
rect 5908 20204 5960 20256
rect 12256 20272 12308 20324
rect 12440 20272 12492 20324
rect 13728 20272 13780 20324
rect 19432 20408 19484 20460
rect 19984 20408 20036 20460
rect 21364 20408 21416 20460
rect 22376 20408 22428 20460
rect 22744 20451 22796 20460
rect 22744 20417 22753 20451
rect 22753 20417 22787 20451
rect 22787 20417 22796 20451
rect 22744 20408 22796 20417
rect 24124 20408 24176 20460
rect 24676 20408 24728 20460
rect 25964 20408 26016 20460
rect 26516 20408 26568 20460
rect 15476 20340 15528 20392
rect 15568 20383 15620 20392
rect 15568 20349 15577 20383
rect 15577 20349 15611 20383
rect 15611 20349 15620 20383
rect 15568 20340 15620 20349
rect 16028 20272 16080 20324
rect 17960 20340 18012 20392
rect 24032 20272 24084 20324
rect 14464 20204 14516 20256
rect 15384 20204 15436 20256
rect 20536 20204 20588 20256
rect 22192 20204 22244 20256
rect 22284 20204 22336 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4528 20000 4580 20052
rect 4896 20000 4948 20052
rect 7196 20000 7248 20052
rect 11980 20000 12032 20052
rect 8300 19975 8352 19984
rect 8300 19941 8309 19975
rect 8309 19941 8343 19975
rect 8343 19941 8352 19975
rect 8300 19932 8352 19941
rect 9772 19932 9824 19984
rect 3792 19864 3844 19916
rect 5080 19907 5132 19916
rect 5080 19873 5089 19907
rect 5089 19873 5123 19907
rect 5123 19873 5132 19907
rect 5080 19864 5132 19873
rect 5448 19864 5500 19916
rect 8392 19864 8444 19916
rect 14740 20000 14792 20052
rect 17224 20000 17276 20052
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 21548 20000 21600 20052
rect 23296 20000 23348 20052
rect 31852 20000 31904 20052
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 10140 19796 10192 19848
rect 3148 19728 3200 19780
rect 3240 19660 3292 19712
rect 5080 19728 5132 19780
rect 5632 19728 5684 19780
rect 5908 19728 5960 19780
rect 6736 19660 6788 19712
rect 7840 19771 7892 19780
rect 7840 19737 7849 19771
rect 7849 19737 7883 19771
rect 7883 19737 7892 19771
rect 7840 19728 7892 19737
rect 8024 19728 8076 19780
rect 10600 19728 10652 19780
rect 10968 19728 11020 19780
rect 11428 19728 11480 19780
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 15200 19932 15252 19984
rect 15568 19975 15620 19984
rect 15568 19941 15577 19975
rect 15577 19941 15611 19975
rect 15611 19941 15620 19975
rect 15568 19932 15620 19941
rect 15384 19907 15436 19916
rect 15384 19873 15393 19907
rect 15393 19873 15427 19907
rect 15427 19873 15436 19907
rect 15384 19864 15436 19873
rect 16212 19864 16264 19916
rect 14556 19796 14608 19848
rect 15752 19796 15804 19848
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 18512 19932 18564 19984
rect 19248 19864 19300 19916
rect 20720 19864 20772 19916
rect 17408 19796 17460 19805
rect 18144 19796 18196 19848
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 19984 19796 20036 19848
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 22376 19932 22428 19984
rect 22928 19932 22980 19984
rect 24400 19932 24452 19984
rect 24216 19864 24268 19916
rect 25412 19864 25464 19916
rect 23296 19839 23348 19848
rect 12440 19728 12492 19780
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 24676 19796 24728 19848
rect 26332 19839 26384 19848
rect 26332 19805 26341 19839
rect 26341 19805 26375 19839
rect 26375 19805 26384 19839
rect 26332 19796 26384 19805
rect 21548 19728 21600 19780
rect 22284 19771 22336 19780
rect 22284 19737 22293 19771
rect 22293 19737 22327 19771
rect 22327 19737 22336 19771
rect 25136 19771 25188 19780
rect 22284 19728 22336 19737
rect 25136 19737 25145 19771
rect 25145 19737 25179 19771
rect 25179 19737 25188 19771
rect 25136 19728 25188 19737
rect 12256 19660 12308 19712
rect 13820 19660 13872 19712
rect 15016 19660 15068 19712
rect 15108 19660 15160 19712
rect 18420 19660 18472 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 19340 19660 19392 19712
rect 20352 19703 20404 19712
rect 20352 19669 20361 19703
rect 20361 19669 20395 19703
rect 20395 19669 20404 19703
rect 20352 19660 20404 19669
rect 26056 19660 26108 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 5448 19456 5500 19508
rect 6000 19456 6052 19508
rect 3792 19431 3844 19440
rect 3792 19397 3801 19431
rect 3801 19397 3835 19431
rect 3835 19397 3844 19431
rect 3792 19388 3844 19397
rect 11888 19456 11940 19508
rect 13820 19456 13872 19508
rect 6920 19388 6972 19440
rect 3148 19320 3200 19372
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 4896 19320 4948 19329
rect 6276 19320 6328 19372
rect 9312 19388 9364 19440
rect 9772 19388 9824 19440
rect 12624 19388 12676 19440
rect 16396 19456 16448 19508
rect 17960 19456 18012 19508
rect 20904 19456 20956 19508
rect 22928 19499 22980 19508
rect 22928 19465 22937 19499
rect 22937 19465 22971 19499
rect 22971 19465 22980 19499
rect 22928 19456 22980 19465
rect 24676 19499 24728 19508
rect 14188 19388 14240 19440
rect 16304 19388 16356 19440
rect 10784 19320 10836 19372
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 12256 19320 12308 19372
rect 1584 19252 1636 19304
rect 3332 19252 3384 19304
rect 4712 19252 4764 19304
rect 5448 19252 5500 19304
rect 6644 19295 6696 19304
rect 6644 19261 6653 19295
rect 6653 19261 6687 19295
rect 6687 19261 6696 19295
rect 6644 19252 6696 19261
rect 7564 19252 7616 19304
rect 6552 19184 6604 19236
rect 7932 19184 7984 19236
rect 9036 19184 9088 19236
rect 10876 19252 10928 19304
rect 11980 19295 12032 19304
rect 11980 19261 11989 19295
rect 11989 19261 12023 19295
rect 12023 19261 12032 19295
rect 11980 19252 12032 19261
rect 4160 19116 4212 19168
rect 4896 19116 4948 19168
rect 9128 19116 9180 19168
rect 12348 19184 12400 19236
rect 12716 19320 12768 19372
rect 15200 19320 15252 19372
rect 17868 19320 17920 19372
rect 21548 19388 21600 19440
rect 23572 19431 23624 19440
rect 13360 19252 13412 19304
rect 13636 19252 13688 19304
rect 13820 19252 13872 19304
rect 14464 19252 14516 19304
rect 14924 19184 14976 19236
rect 15108 19295 15160 19304
rect 15108 19261 15117 19295
rect 15117 19261 15151 19295
rect 15151 19261 15160 19295
rect 15108 19252 15160 19261
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 17316 19252 17368 19304
rect 19340 19252 19392 19304
rect 20352 19320 20404 19372
rect 23572 19397 23581 19431
rect 23581 19397 23615 19431
rect 23615 19397 23624 19431
rect 23572 19388 23624 19397
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 25136 19456 25188 19508
rect 34060 19388 34112 19440
rect 22192 19320 22244 19372
rect 22836 19320 22888 19372
rect 20260 19252 20312 19304
rect 21272 19252 21324 19304
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 22468 19295 22520 19304
rect 22468 19261 22477 19295
rect 22477 19261 22511 19295
rect 22511 19261 22520 19295
rect 22468 19252 22520 19261
rect 25412 19363 25464 19372
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 26056 19363 26108 19372
rect 26056 19329 26065 19363
rect 26065 19329 26099 19363
rect 26099 19329 26108 19363
rect 26056 19320 26108 19329
rect 15476 19227 15528 19236
rect 15476 19193 15485 19227
rect 15485 19193 15519 19227
rect 15519 19193 15528 19227
rect 15476 19184 15528 19193
rect 11060 19116 11112 19168
rect 12072 19116 12124 19168
rect 12164 19116 12216 19168
rect 22744 19184 22796 19236
rect 16304 19116 16356 19168
rect 19064 19116 19116 19168
rect 19248 19116 19300 19168
rect 22376 19116 22428 19168
rect 23940 19184 23992 19236
rect 27528 19184 27580 19236
rect 25228 19159 25280 19168
rect 25228 19125 25237 19159
rect 25237 19125 25271 19159
rect 25271 19125 25280 19159
rect 25228 19116 25280 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3332 18955 3384 18964
rect 3332 18921 3341 18955
rect 3341 18921 3375 18955
rect 3375 18921 3384 18955
rect 3332 18912 3384 18921
rect 7564 18844 7616 18896
rect 8300 18844 8352 18896
rect 10048 18912 10100 18964
rect 13912 18912 13964 18964
rect 14372 18912 14424 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 15660 18912 15712 18964
rect 18052 18912 18104 18964
rect 30012 18912 30064 18964
rect 12072 18887 12124 18896
rect 4896 18776 4948 18828
rect 8944 18776 8996 18828
rect 9772 18776 9824 18828
rect 12072 18853 12081 18887
rect 12081 18853 12115 18887
rect 12115 18853 12124 18887
rect 12072 18844 12124 18853
rect 23940 18887 23992 18896
rect 1584 18751 1636 18760
rect 1584 18717 1593 18751
rect 1593 18717 1627 18751
rect 1627 18717 1636 18751
rect 1584 18708 1636 18717
rect 5816 18708 5868 18760
rect 6920 18708 6972 18760
rect 7196 18708 7248 18760
rect 8300 18708 8352 18760
rect 10140 18708 10192 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 1216 18572 1268 18624
rect 4988 18640 5040 18692
rect 6644 18640 6696 18692
rect 6736 18640 6788 18692
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 8576 18640 8628 18692
rect 10324 18640 10376 18692
rect 10600 18683 10652 18692
rect 10600 18649 10609 18683
rect 10609 18649 10643 18683
rect 10643 18649 10652 18683
rect 10600 18640 10652 18649
rect 11612 18640 11664 18692
rect 8852 18572 8904 18624
rect 13360 18708 13412 18760
rect 15016 18708 15068 18760
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 19064 18776 19116 18828
rect 20076 18776 20128 18828
rect 22284 18776 22336 18828
rect 22928 18776 22980 18828
rect 23940 18853 23949 18887
rect 23949 18853 23983 18887
rect 23983 18853 23992 18887
rect 23940 18844 23992 18853
rect 16304 18708 16356 18760
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 17592 18751 17644 18760
rect 14280 18640 14332 18692
rect 16856 18640 16908 18692
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 17960 18708 18012 18760
rect 19524 18708 19576 18760
rect 22100 18708 22152 18760
rect 24124 18708 24176 18760
rect 26332 18708 26384 18760
rect 18696 18640 18748 18692
rect 23480 18683 23532 18692
rect 23480 18649 23489 18683
rect 23489 18649 23523 18683
rect 23523 18649 23532 18683
rect 23480 18640 23532 18649
rect 13360 18572 13412 18624
rect 15660 18572 15712 18624
rect 16304 18615 16356 18624
rect 16304 18581 16313 18615
rect 16313 18581 16347 18615
rect 16347 18581 16356 18615
rect 16304 18572 16356 18581
rect 18144 18572 18196 18624
rect 19156 18572 19208 18624
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 22928 18572 22980 18624
rect 25320 18615 25372 18624
rect 25320 18581 25329 18615
rect 25329 18581 25363 18615
rect 25363 18581 25372 18615
rect 25320 18572 25372 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 2872 18368 2924 18420
rect 4804 18368 4856 18420
rect 9128 18368 9180 18420
rect 9404 18368 9456 18420
rect 12164 18368 12216 18420
rect 6644 18300 6696 18352
rect 2504 18232 2556 18284
rect 3608 18232 3660 18284
rect 3792 18164 3844 18216
rect 4896 18232 4948 18284
rect 5632 18232 5684 18284
rect 4988 18096 5040 18148
rect 5080 18096 5132 18148
rect 5816 18139 5868 18148
rect 5816 18105 5825 18139
rect 5825 18105 5859 18139
rect 5859 18105 5868 18139
rect 5816 18096 5868 18105
rect 6736 18232 6788 18284
rect 7196 18232 7248 18284
rect 7104 18164 7156 18216
rect 7840 18300 7892 18352
rect 9128 18232 9180 18284
rect 9772 18232 9824 18284
rect 10140 18300 10192 18352
rect 10876 18300 10928 18352
rect 11888 18343 11940 18352
rect 10508 18232 10560 18284
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 11888 18309 11897 18343
rect 11897 18309 11931 18343
rect 11931 18309 11940 18343
rect 11888 18300 11940 18309
rect 17040 18368 17092 18420
rect 17132 18368 17184 18420
rect 21272 18411 21324 18420
rect 17684 18300 17736 18352
rect 10048 18164 10100 18216
rect 13912 18232 13964 18284
rect 15200 18232 15252 18284
rect 16304 18275 16356 18284
rect 16304 18241 16313 18275
rect 16313 18241 16347 18275
rect 16347 18241 16356 18275
rect 16304 18232 16356 18241
rect 18052 18300 18104 18352
rect 19156 18343 19208 18352
rect 19156 18309 19165 18343
rect 19165 18309 19199 18343
rect 19199 18309 19208 18343
rect 19156 18300 19208 18309
rect 20628 18300 20680 18352
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 23572 18368 23624 18420
rect 7656 18028 7708 18080
rect 8208 18096 8260 18148
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 13728 18164 13780 18216
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 20904 18232 20956 18284
rect 22376 18232 22428 18284
rect 22928 18275 22980 18284
rect 22928 18241 22937 18275
rect 22937 18241 22971 18275
rect 22971 18241 22980 18275
rect 22928 18232 22980 18241
rect 23480 18300 23532 18352
rect 25412 18300 25464 18352
rect 25228 18232 25280 18284
rect 10508 18028 10560 18080
rect 11336 18028 11388 18080
rect 12164 18096 12216 18148
rect 12348 18139 12400 18148
rect 12348 18105 12357 18139
rect 12357 18105 12391 18139
rect 12391 18105 12400 18139
rect 12348 18096 12400 18105
rect 17132 18096 17184 18148
rect 22652 18164 22704 18216
rect 23296 18164 23348 18216
rect 24032 18164 24084 18216
rect 20260 18096 20312 18148
rect 20628 18096 20680 18148
rect 12624 18028 12676 18080
rect 13084 18028 13136 18080
rect 18052 18028 18104 18080
rect 19248 18028 19300 18080
rect 22376 18028 22428 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4436 17756 4488 17808
rect 3700 17688 3752 17740
rect 1952 17663 2004 17672
rect 1952 17629 1961 17663
rect 1961 17629 1995 17663
rect 1995 17629 2004 17663
rect 1952 17620 2004 17629
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 7104 17824 7156 17876
rect 9680 17867 9732 17876
rect 5172 17756 5224 17808
rect 5448 17756 5500 17808
rect 6552 17756 6604 17808
rect 6460 17731 6512 17740
rect 3976 17552 4028 17604
rect 4068 17552 4120 17604
rect 6460 17697 6469 17731
rect 6469 17697 6503 17731
rect 6503 17697 6512 17731
rect 6460 17688 6512 17697
rect 6644 17731 6696 17740
rect 6644 17697 6653 17731
rect 6653 17697 6687 17731
rect 6687 17697 6696 17731
rect 6644 17688 6696 17697
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 8208 17799 8260 17808
rect 8208 17765 8217 17799
rect 8217 17765 8251 17799
rect 8251 17765 8260 17799
rect 8208 17756 8260 17765
rect 8668 17756 8720 17808
rect 10600 17756 10652 17808
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 9220 17688 9272 17740
rect 9404 17688 9456 17740
rect 11796 17824 11848 17876
rect 11244 17688 11296 17740
rect 12624 17731 12676 17740
rect 7196 17620 7248 17672
rect 10508 17663 10560 17672
rect 10508 17629 10517 17663
rect 10517 17629 10551 17663
rect 10551 17629 10560 17663
rect 10508 17620 10560 17629
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 12624 17697 12633 17731
rect 12633 17697 12667 17731
rect 12667 17697 12676 17731
rect 12624 17688 12676 17697
rect 13084 17731 13136 17740
rect 13084 17697 13093 17731
rect 13093 17697 13127 17731
rect 13127 17697 13136 17731
rect 13084 17688 13136 17697
rect 12532 17620 12584 17672
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14924 17688 14976 17740
rect 15108 17620 15160 17672
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 18880 17824 18932 17876
rect 19432 17867 19484 17876
rect 19432 17833 19441 17867
rect 19441 17833 19475 17867
rect 19475 17833 19484 17867
rect 19432 17824 19484 17833
rect 17132 17799 17184 17808
rect 17132 17765 17141 17799
rect 17141 17765 17175 17799
rect 17175 17765 17184 17799
rect 17132 17756 17184 17765
rect 17684 17731 17736 17740
rect 17684 17697 17693 17731
rect 17693 17697 17727 17731
rect 17727 17697 17736 17731
rect 17684 17688 17736 17697
rect 24400 17756 24452 17808
rect 18144 17620 18196 17672
rect 18788 17620 18840 17672
rect 20260 17663 20312 17672
rect 20260 17629 20269 17663
rect 20269 17629 20303 17663
rect 20303 17629 20312 17663
rect 20260 17620 20312 17629
rect 20904 17620 20956 17672
rect 24400 17620 24452 17672
rect 25872 17620 25924 17672
rect 4804 17484 4856 17536
rect 5172 17484 5224 17536
rect 5356 17595 5408 17604
rect 5356 17561 5365 17595
rect 5365 17561 5399 17595
rect 5399 17561 5408 17595
rect 5356 17552 5408 17561
rect 5448 17484 5500 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 7748 17595 7800 17604
rect 7748 17561 7757 17595
rect 7757 17561 7791 17595
rect 7791 17561 7800 17595
rect 7748 17552 7800 17561
rect 8024 17552 8076 17604
rect 9404 17484 9456 17536
rect 13084 17484 13136 17536
rect 13452 17484 13504 17536
rect 23204 17552 23256 17604
rect 25320 17552 25372 17604
rect 18052 17484 18104 17536
rect 21456 17484 21508 17536
rect 23572 17484 23624 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7104 17280 7156 17332
rect 1492 17212 1544 17264
rect 5080 17212 5132 17264
rect 1676 17144 1728 17196
rect 6920 17212 6972 17264
rect 8300 17212 8352 17264
rect 8852 17255 8904 17264
rect 8852 17221 8861 17255
rect 8861 17221 8895 17255
rect 8895 17221 8904 17255
rect 8852 17212 8904 17221
rect 9772 17212 9824 17264
rect 10692 17212 10744 17264
rect 8668 17144 8720 17196
rect 9128 17144 9180 17196
rect 11060 17280 11112 17332
rect 13452 17280 13504 17332
rect 13636 17280 13688 17332
rect 12624 17212 12676 17264
rect 17040 17280 17092 17332
rect 18144 17323 18196 17332
rect 18144 17289 18153 17323
rect 18153 17289 18187 17323
rect 18187 17289 18196 17323
rect 18144 17280 18196 17289
rect 18788 17323 18840 17332
rect 18788 17289 18797 17323
rect 18797 17289 18831 17323
rect 18831 17289 18840 17323
rect 18788 17280 18840 17289
rect 22836 17323 22888 17332
rect 22836 17289 22845 17323
rect 22845 17289 22879 17323
rect 22879 17289 22888 17323
rect 22836 17280 22888 17289
rect 22284 17212 22336 17264
rect 4896 17119 4948 17128
rect 1584 17008 1636 17060
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 8116 16940 8168 16992
rect 8392 16940 8444 16992
rect 10232 17076 10284 17128
rect 10416 17076 10468 17128
rect 14280 17144 14332 17196
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 16488 17144 16540 17196
rect 17592 17144 17644 17196
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 19616 17187 19668 17196
rect 18972 17144 19024 17153
rect 14188 17076 14240 17128
rect 14832 17076 14884 17128
rect 15844 17076 15896 17128
rect 16028 17076 16080 17128
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 20352 17144 20404 17196
rect 21456 17187 21508 17196
rect 21456 17153 21465 17187
rect 21465 17153 21499 17187
rect 21499 17153 21508 17187
rect 21456 17144 21508 17153
rect 22376 17187 22428 17196
rect 22376 17153 22385 17187
rect 22385 17153 22419 17187
rect 22419 17153 22428 17187
rect 22376 17144 22428 17153
rect 23572 17144 23624 17196
rect 23940 17144 23992 17196
rect 38292 17187 38344 17196
rect 38292 17153 38301 17187
rect 38301 17153 38335 17187
rect 38335 17153 38344 17187
rect 38292 17144 38344 17153
rect 22192 17119 22244 17128
rect 9496 16940 9548 16992
rect 13452 17008 13504 17060
rect 14924 17008 14976 17060
rect 15476 17008 15528 17060
rect 11704 16940 11756 16992
rect 11796 16940 11848 16992
rect 16672 16940 16724 16992
rect 20260 17008 20312 17060
rect 22192 17085 22201 17119
rect 22201 17085 22235 17119
rect 22235 17085 22244 17119
rect 22192 17076 22244 17085
rect 22560 17008 22612 17060
rect 24584 17076 24636 17128
rect 19340 16940 19392 16992
rect 20720 16940 20772 16992
rect 21364 16940 21416 16992
rect 23204 16940 23256 16992
rect 24492 16983 24544 16992
rect 24492 16949 24501 16983
rect 24501 16949 24535 16983
rect 24535 16949 24544 16983
rect 24492 16940 24544 16949
rect 25688 16983 25740 16992
rect 25688 16949 25697 16983
rect 25697 16949 25731 16983
rect 25731 16949 25740 16983
rect 25688 16940 25740 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4896 16736 4948 16788
rect 11060 16736 11112 16788
rect 15200 16736 15252 16788
rect 18144 16736 18196 16788
rect 19616 16736 19668 16788
rect 21548 16779 21600 16788
rect 21548 16745 21557 16779
rect 21557 16745 21591 16779
rect 21591 16745 21600 16779
rect 21548 16736 21600 16745
rect 23204 16779 23256 16788
rect 23204 16745 23213 16779
rect 23213 16745 23247 16779
rect 23247 16745 23256 16779
rect 23204 16736 23256 16745
rect 5816 16668 5868 16720
rect 6736 16668 6788 16720
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2596 16600 2648 16652
rect 8392 16668 8444 16720
rect 7380 16600 7432 16652
rect 8024 16600 8076 16652
rect 17408 16668 17460 16720
rect 10600 16600 10652 16652
rect 13728 16600 13780 16652
rect 13820 16600 13872 16652
rect 33416 16668 33468 16720
rect 18144 16643 18196 16652
rect 18144 16609 18153 16643
rect 18153 16609 18187 16643
rect 18187 16609 18196 16643
rect 18144 16600 18196 16609
rect 21180 16643 21232 16652
rect 21180 16609 21189 16643
rect 21189 16609 21223 16643
rect 21223 16609 21232 16643
rect 21180 16600 21232 16609
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 22560 16643 22612 16652
rect 22560 16609 22569 16643
rect 22569 16609 22603 16643
rect 22603 16609 22612 16643
rect 22560 16600 22612 16609
rect 24584 16643 24636 16652
rect 24584 16609 24593 16643
rect 24593 16609 24627 16643
rect 24627 16609 24636 16643
rect 24584 16600 24636 16609
rect 1584 16532 1636 16584
rect 9128 16575 9180 16584
rect 2964 16464 3016 16516
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 4160 16464 4212 16516
rect 4896 16464 4948 16516
rect 6276 16507 6328 16516
rect 6276 16473 6285 16507
rect 6285 16473 6319 16507
rect 6319 16473 6328 16507
rect 6276 16464 6328 16473
rect 5540 16396 5592 16448
rect 5724 16439 5776 16448
rect 5724 16405 5733 16439
rect 5733 16405 5767 16439
rect 5767 16405 5776 16439
rect 5724 16396 5776 16405
rect 6092 16396 6144 16448
rect 7656 16507 7708 16516
rect 7656 16473 7665 16507
rect 7665 16473 7699 16507
rect 7699 16473 7708 16507
rect 7656 16464 7708 16473
rect 9404 16507 9456 16516
rect 7196 16396 7248 16448
rect 8024 16396 8076 16448
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 9496 16464 9548 16516
rect 12164 16532 12216 16584
rect 14280 16532 14332 16584
rect 16396 16532 16448 16584
rect 20168 16532 20220 16584
rect 20352 16532 20404 16584
rect 22744 16575 22796 16584
rect 22744 16541 22753 16575
rect 22753 16541 22787 16575
rect 22787 16541 22796 16575
rect 22744 16532 22796 16541
rect 23572 16532 23624 16584
rect 24400 16532 24452 16584
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 14648 16464 14700 16516
rect 15200 16507 15252 16516
rect 15200 16473 15209 16507
rect 15209 16473 15243 16507
rect 15243 16473 15252 16507
rect 15200 16464 15252 16473
rect 15384 16464 15436 16516
rect 15844 16507 15896 16516
rect 15844 16473 15853 16507
rect 15853 16473 15887 16507
rect 15887 16473 15896 16507
rect 15844 16464 15896 16473
rect 8392 16396 8444 16448
rect 11152 16396 11204 16448
rect 12624 16396 12676 16448
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 12716 16396 12768 16405
rect 14464 16396 14516 16448
rect 15476 16396 15528 16448
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 23664 16439 23716 16448
rect 23664 16405 23673 16439
rect 23673 16405 23707 16439
rect 23707 16405 23716 16439
rect 23664 16396 23716 16405
rect 24032 16396 24084 16448
rect 29736 16396 29788 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2044 16192 2096 16244
rect 4988 16192 5040 16244
rect 7656 16192 7708 16244
rect 3332 16124 3384 16176
rect 3608 16167 3660 16176
rect 3608 16133 3617 16167
rect 3617 16133 3651 16167
rect 3651 16133 3660 16167
rect 3608 16124 3660 16133
rect 5356 16124 5408 16176
rect 5724 16124 5776 16176
rect 7196 16124 7248 16176
rect 10140 16124 10192 16176
rect 11520 16192 11572 16244
rect 13820 16192 13872 16244
rect 12256 16124 12308 16176
rect 1584 16031 1636 16040
rect 1584 15997 1593 16031
rect 1593 15997 1627 16031
rect 1627 15997 1636 16031
rect 1584 15988 1636 15997
rect 3240 15988 3292 16040
rect 4068 16031 4120 16040
rect 4068 15997 4077 16031
rect 4077 15997 4111 16031
rect 4111 15997 4120 16031
rect 4068 15988 4120 15997
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 8576 16056 8628 16108
rect 9128 16056 9180 16108
rect 11152 16056 11204 16108
rect 13360 16124 13412 16176
rect 16120 16192 16172 16244
rect 14096 16167 14148 16176
rect 14096 16133 14105 16167
rect 14105 16133 14139 16167
rect 14139 16133 14148 16167
rect 14096 16124 14148 16133
rect 14464 16124 14516 16176
rect 18328 16167 18380 16176
rect 13820 16056 13872 16108
rect 18328 16133 18337 16167
rect 18337 16133 18371 16167
rect 18371 16133 18380 16167
rect 18328 16124 18380 16133
rect 19432 16124 19484 16176
rect 20168 16192 20220 16244
rect 22744 16235 22796 16244
rect 22744 16201 22753 16235
rect 22753 16201 22787 16235
rect 22787 16201 22796 16235
rect 22744 16192 22796 16201
rect 24032 16235 24084 16244
rect 24032 16201 24041 16235
rect 24041 16201 24075 16235
rect 24075 16201 24084 16235
rect 24032 16192 24084 16201
rect 24768 16192 24820 16244
rect 21640 16124 21692 16176
rect 6184 15988 6236 16040
rect 10048 15988 10100 16040
rect 10968 15988 11020 16040
rect 11520 15988 11572 16040
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 11888 16031 11940 16040
rect 11888 15997 11897 16031
rect 11897 15997 11931 16031
rect 11931 15997 11940 16031
rect 11888 15988 11940 15997
rect 14004 16031 14056 16040
rect 14004 15997 14013 16031
rect 14013 15997 14047 16031
rect 14047 15997 14056 16031
rect 14004 15988 14056 15997
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 6000 15852 6052 15904
rect 9404 15852 9456 15904
rect 14556 15963 14608 15972
rect 14556 15929 14565 15963
rect 14565 15929 14599 15963
rect 14599 15929 14608 15963
rect 14556 15920 14608 15929
rect 10876 15852 10928 15904
rect 13636 15852 13688 15904
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 17040 16031 17092 16040
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 19432 16031 19484 16040
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 20076 15988 20128 16040
rect 24860 16124 24912 16176
rect 18512 15920 18564 15972
rect 23664 16056 23716 16108
rect 25688 16056 25740 16108
rect 29736 16099 29788 16108
rect 29736 16065 29745 16099
rect 29745 16065 29779 16099
rect 29779 16065 29788 16099
rect 29736 16056 29788 16065
rect 36084 16056 36136 16108
rect 23112 15988 23164 16040
rect 24492 15988 24544 16040
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 20260 15852 20312 15904
rect 31668 15852 31720 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6276 15648 6328 15700
rect 6552 15648 6604 15700
rect 11152 15648 11204 15700
rect 13912 15648 13964 15700
rect 17040 15648 17092 15700
rect 20260 15691 20312 15700
rect 20260 15657 20269 15691
rect 20269 15657 20303 15691
rect 20303 15657 20312 15691
rect 20260 15648 20312 15657
rect 7932 15580 7984 15632
rect 8944 15580 8996 15632
rect 10876 15580 10928 15632
rect 2136 15555 2188 15564
rect 2136 15521 2145 15555
rect 2145 15521 2179 15555
rect 2179 15521 2188 15555
rect 2136 15512 2188 15521
rect 2872 15512 2924 15564
rect 3056 15512 3108 15564
rect 6736 15512 6788 15564
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 8392 15512 8444 15564
rect 15476 15580 15528 15632
rect 16856 15623 16908 15632
rect 16856 15589 16865 15623
rect 16865 15589 16899 15623
rect 16899 15589 16908 15623
rect 16856 15580 16908 15589
rect 12808 15512 12860 15564
rect 14556 15512 14608 15564
rect 18052 15580 18104 15632
rect 9588 15487 9640 15496
rect 4620 15376 4672 15428
rect 5448 15376 5500 15428
rect 6460 15376 6512 15428
rect 7748 15419 7800 15428
rect 7748 15385 7757 15419
rect 7757 15385 7791 15419
rect 7791 15385 7800 15419
rect 7748 15376 7800 15385
rect 8024 15376 8076 15428
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 11980 15444 12032 15496
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 14832 15444 14884 15496
rect 11796 15376 11848 15428
rect 12808 15376 12860 15428
rect 15292 15419 15344 15428
rect 15292 15385 15301 15419
rect 15301 15385 15335 15419
rect 15335 15385 15344 15419
rect 15292 15376 15344 15385
rect 15752 15376 15804 15428
rect 17868 15512 17920 15564
rect 19340 15512 19392 15564
rect 20168 15512 20220 15564
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 25688 15512 25740 15564
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 16488 15444 16540 15453
rect 16948 15444 17000 15496
rect 20444 15444 20496 15496
rect 20812 15444 20864 15496
rect 24124 15444 24176 15496
rect 25136 15444 25188 15496
rect 17224 15376 17276 15428
rect 17776 15419 17828 15428
rect 17776 15385 17785 15419
rect 17785 15385 17819 15419
rect 17819 15385 17828 15419
rect 17776 15376 17828 15385
rect 19984 15376 20036 15428
rect 22744 15376 22796 15428
rect 3792 15308 3844 15360
rect 9588 15308 9640 15360
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 12716 15308 12768 15317
rect 21364 15351 21416 15360
rect 21364 15317 21373 15351
rect 21373 15317 21407 15351
rect 21407 15317 21416 15351
rect 21364 15308 21416 15317
rect 22928 15351 22980 15360
rect 22928 15317 22937 15351
rect 22937 15317 22971 15351
rect 22971 15317 22980 15351
rect 22928 15308 22980 15317
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 23388 15308 23440 15317
rect 24676 15351 24728 15360
rect 24676 15317 24685 15351
rect 24685 15317 24719 15351
rect 24719 15317 24728 15351
rect 24676 15308 24728 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2504 15036 2556 15088
rect 3516 15036 3568 15088
rect 3792 15079 3844 15088
rect 3792 15045 3801 15079
rect 3801 15045 3835 15079
rect 3835 15045 3844 15079
rect 3792 15036 3844 15045
rect 4068 14968 4120 15020
rect 5448 15104 5500 15156
rect 6552 15104 6604 15156
rect 6736 15104 6788 15156
rect 9496 15104 9548 15156
rect 9772 15104 9824 15156
rect 4988 15036 5040 15088
rect 6276 15036 6328 15088
rect 7104 15036 7156 15088
rect 7840 15036 7892 15088
rect 9128 15036 9180 15088
rect 10232 14968 10284 15020
rect 12348 15036 12400 15088
rect 13820 15104 13872 15156
rect 16856 15104 16908 15156
rect 17408 15079 17460 15088
rect 17408 15045 17417 15079
rect 17417 15045 17451 15079
rect 17451 15045 17460 15079
rect 17408 15036 17460 15045
rect 18328 15104 18380 15156
rect 22928 15147 22980 15156
rect 19248 15079 19300 15088
rect 19248 15045 19257 15079
rect 19257 15045 19291 15079
rect 19291 15045 19300 15079
rect 19248 15036 19300 15045
rect 19984 15036 20036 15088
rect 22928 15113 22937 15147
rect 22937 15113 22971 15147
rect 22971 15113 22980 15147
rect 22928 15104 22980 15113
rect 23204 15104 23256 15156
rect 23940 15036 23992 15088
rect 1676 14900 1728 14952
rect 3424 14900 3476 14952
rect 5816 14900 5868 14952
rect 6552 14943 6604 14952
rect 6552 14909 6561 14943
rect 6561 14909 6595 14943
rect 6595 14909 6604 14943
rect 6552 14900 6604 14909
rect 7196 14900 7248 14952
rect 9128 14943 9180 14952
rect 2688 14764 2740 14816
rect 6184 14832 6236 14884
rect 5632 14764 5684 14816
rect 8116 14764 8168 14816
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 13544 14968 13596 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 22192 14968 22244 15020
rect 23388 14968 23440 15020
rect 36084 15104 36136 15156
rect 31668 15036 31720 15088
rect 9128 14900 9180 14909
rect 10692 14900 10744 14952
rect 12532 14900 12584 14952
rect 13268 14900 13320 14952
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 17316 14943 17368 14952
rect 11244 14764 11296 14816
rect 11336 14764 11388 14816
rect 13820 14832 13872 14884
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 20076 14900 20128 14952
rect 25320 14943 25372 14952
rect 17868 14875 17920 14884
rect 17868 14841 17877 14875
rect 17877 14841 17911 14875
rect 17911 14841 17920 14875
rect 17868 14832 17920 14841
rect 19340 14832 19392 14884
rect 24124 14875 24176 14884
rect 24124 14841 24133 14875
rect 24133 14841 24167 14875
rect 24167 14841 24176 14875
rect 24124 14832 24176 14841
rect 25320 14909 25329 14943
rect 25329 14909 25363 14943
rect 25363 14909 25372 14943
rect 25320 14900 25372 14909
rect 26516 14900 26568 14952
rect 33600 14968 33652 15020
rect 37188 14900 37240 14952
rect 12992 14764 13044 14816
rect 17500 14764 17552 14816
rect 20720 14764 20772 14816
rect 20812 14764 20864 14816
rect 23296 14764 23348 14816
rect 25228 14764 25280 14816
rect 38016 14764 38068 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 6276 14560 6328 14612
rect 9128 14560 9180 14612
rect 10048 14560 10100 14612
rect 12624 14560 12676 14612
rect 13728 14560 13780 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 15936 14560 15988 14612
rect 17500 14560 17552 14612
rect 18144 14560 18196 14612
rect 2688 14424 2740 14476
rect 8116 14492 8168 14544
rect 8392 14424 8444 14476
rect 9036 14424 9088 14476
rect 10508 14492 10560 14544
rect 10600 14492 10652 14544
rect 13268 14492 13320 14544
rect 10784 14424 10836 14476
rect 12716 14424 12768 14476
rect 25228 14535 25280 14544
rect 13820 14424 13872 14476
rect 13912 14424 13964 14476
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4068 14356 4120 14408
rect 6736 14356 6788 14408
rect 12900 14356 12952 14408
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 15568 14424 15620 14476
rect 16028 14424 16080 14476
rect 16856 14424 16908 14476
rect 17592 14424 17644 14476
rect 19432 14424 19484 14476
rect 20260 14424 20312 14476
rect 21272 14424 21324 14476
rect 22560 14424 22612 14476
rect 24676 14424 24728 14476
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 16580 14356 16632 14408
rect 2964 14288 3016 14340
rect 4528 14288 4580 14340
rect 5448 14288 5500 14340
rect 7196 14288 7248 14340
rect 4804 14220 4856 14272
rect 7012 14220 7064 14272
rect 7288 14220 7340 14272
rect 7380 14220 7432 14272
rect 9312 14288 9364 14340
rect 9680 14288 9732 14340
rect 11520 14331 11572 14340
rect 11520 14297 11529 14331
rect 11529 14297 11563 14331
rect 11563 14297 11572 14331
rect 12072 14331 12124 14340
rect 11520 14288 11572 14297
rect 12072 14297 12081 14331
rect 12081 14297 12115 14331
rect 12115 14297 12124 14331
rect 12072 14288 12124 14297
rect 13084 14288 13136 14340
rect 16028 14288 16080 14340
rect 16672 14288 16724 14340
rect 8668 14220 8720 14272
rect 9496 14220 9548 14272
rect 15936 14220 15988 14272
rect 16764 14263 16816 14272
rect 16764 14229 16773 14263
rect 16773 14229 16807 14263
rect 16807 14229 16816 14263
rect 16764 14220 16816 14229
rect 17408 14331 17460 14340
rect 17408 14297 17417 14331
rect 17417 14297 17451 14331
rect 17451 14297 17460 14331
rect 17408 14288 17460 14297
rect 22100 14356 22152 14408
rect 20260 14288 20312 14340
rect 20628 14288 20680 14340
rect 20720 14331 20772 14340
rect 20720 14297 20729 14331
rect 20729 14297 20763 14331
rect 20763 14297 20772 14331
rect 20720 14288 20772 14297
rect 21548 14288 21600 14340
rect 23112 14220 23164 14272
rect 23848 14220 23900 14272
rect 25228 14501 25237 14535
rect 25237 14501 25271 14535
rect 25271 14501 25280 14535
rect 25228 14492 25280 14501
rect 25320 14492 25372 14544
rect 25964 14424 26016 14476
rect 26332 14424 26384 14476
rect 27804 14424 27856 14476
rect 25688 14399 25740 14408
rect 25688 14365 25697 14399
rect 25697 14365 25731 14399
rect 25731 14365 25740 14399
rect 25688 14356 25740 14365
rect 26976 14399 27028 14408
rect 26240 14288 26292 14340
rect 25872 14220 25924 14272
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 33600 14560 33652 14612
rect 29920 14399 29972 14408
rect 29920 14365 29929 14399
rect 29929 14365 29963 14399
rect 29963 14365 29972 14399
rect 29920 14356 29972 14365
rect 38292 14399 38344 14408
rect 32404 14288 32456 14340
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 5172 14016 5224 14068
rect 7380 14016 7432 14068
rect 10048 14016 10100 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 13084 14016 13136 14068
rect 5540 13948 5592 14000
rect 1492 13880 1544 13932
rect 1860 13880 1912 13932
rect 8116 13948 8168 14000
rect 6736 13880 6788 13932
rect 8760 13948 8812 14000
rect 8944 13948 8996 14000
rect 9772 13948 9824 14000
rect 12992 13948 13044 14000
rect 16764 14016 16816 14068
rect 17776 14016 17828 14068
rect 19340 14016 19392 14068
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 22100 14059 22152 14068
rect 13728 13948 13780 14000
rect 14188 13948 14240 14000
rect 16672 13948 16724 14000
rect 17040 13991 17092 14000
rect 17040 13957 17049 13991
rect 17049 13957 17083 13991
rect 17083 13957 17092 13991
rect 17040 13948 17092 13957
rect 17592 13991 17644 14000
rect 17592 13957 17601 13991
rect 17601 13957 17635 13991
rect 17635 13957 17644 13991
rect 17592 13948 17644 13957
rect 20904 13991 20956 14000
rect 3516 13855 3568 13864
rect 2320 13744 2372 13796
rect 1768 13676 1820 13728
rect 2964 13676 3016 13728
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 4712 13812 4764 13864
rect 6368 13812 6420 13864
rect 7012 13812 7064 13864
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 9680 13812 9732 13864
rect 11060 13812 11112 13864
rect 11428 13812 11480 13864
rect 12808 13812 12860 13864
rect 14740 13880 14792 13932
rect 18328 13923 18380 13932
rect 14924 13812 14976 13864
rect 15108 13855 15160 13864
rect 15108 13821 15117 13855
rect 15117 13821 15151 13855
rect 15151 13821 15160 13855
rect 15108 13812 15160 13821
rect 16120 13812 16172 13864
rect 18328 13889 18337 13923
rect 18337 13889 18371 13923
rect 18371 13889 18380 13923
rect 18328 13880 18380 13889
rect 18788 13923 18840 13932
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 20904 13957 20913 13991
rect 20913 13957 20947 13991
rect 20947 13957 20956 13991
rect 20904 13948 20956 13957
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 22100 14016 22152 14025
rect 23848 14059 23900 14068
rect 23848 14025 23857 14059
rect 23857 14025 23891 14059
rect 23891 14025 23900 14059
rect 23848 14016 23900 14025
rect 25320 14059 25372 14068
rect 25320 14025 25329 14059
rect 25329 14025 25363 14059
rect 25363 14025 25372 14059
rect 25320 14016 25372 14025
rect 26516 14059 26568 14068
rect 26516 14025 26525 14059
rect 26525 14025 26559 14059
rect 26559 14025 26568 14059
rect 26516 14016 26568 14025
rect 22560 13948 22612 14000
rect 25228 13948 25280 14000
rect 29920 13948 29972 14000
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 24584 13880 24636 13932
rect 25780 13923 25832 13932
rect 25780 13889 25789 13923
rect 25789 13889 25823 13923
rect 25823 13889 25832 13923
rect 25780 13880 25832 13889
rect 26240 13880 26292 13932
rect 20168 13812 20220 13864
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 22192 13812 22244 13864
rect 22836 13812 22888 13864
rect 24216 13812 24268 13864
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 4068 13676 4120 13728
rect 4712 13676 4764 13728
rect 9680 13676 9732 13728
rect 10324 13676 10376 13728
rect 11152 13676 11204 13728
rect 11244 13676 11296 13728
rect 12624 13676 12676 13728
rect 14648 13676 14700 13728
rect 16764 13676 16816 13728
rect 26240 13676 26292 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 3608 13472 3660 13524
rect 4712 13472 4764 13524
rect 11244 13472 11296 13524
rect 6736 13379 6788 13388
rect 6736 13345 6745 13379
rect 6745 13345 6779 13379
rect 6779 13345 6788 13379
rect 6736 13336 6788 13345
rect 8484 13336 8536 13388
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 9036 13336 9088 13388
rect 13360 13472 13412 13524
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 14740 13515 14792 13524
rect 14740 13481 14749 13515
rect 14749 13481 14783 13515
rect 14783 13481 14792 13515
rect 14740 13472 14792 13481
rect 14924 13472 14976 13524
rect 17040 13472 17092 13524
rect 20904 13472 20956 13524
rect 22560 13515 22612 13524
rect 22560 13481 22569 13515
rect 22569 13481 22603 13515
rect 22603 13481 22612 13515
rect 22560 13472 22612 13481
rect 25872 13515 25924 13524
rect 25872 13481 25881 13515
rect 25881 13481 25915 13515
rect 25915 13481 25924 13515
rect 25872 13472 25924 13481
rect 26976 13472 27028 13524
rect 11612 13404 11664 13456
rect 13452 13404 13504 13456
rect 13728 13404 13780 13456
rect 14648 13404 14700 13456
rect 14832 13404 14884 13456
rect 20076 13404 20128 13456
rect 20996 13404 21048 13456
rect 21364 13447 21416 13456
rect 21364 13413 21373 13447
rect 21373 13413 21407 13447
rect 21407 13413 21416 13447
rect 21364 13404 21416 13413
rect 3700 13200 3752 13252
rect 5724 13200 5776 13252
rect 2964 13132 3016 13184
rect 7748 13200 7800 13252
rect 11704 13268 11756 13320
rect 11796 13268 11848 13320
rect 12348 13268 12400 13320
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 8392 13200 8444 13252
rect 8852 13200 8904 13252
rect 9404 13243 9456 13252
rect 9404 13209 9413 13243
rect 9413 13209 9447 13243
rect 9447 13209 9456 13243
rect 9404 13200 9456 13209
rect 9956 13200 10008 13252
rect 10784 13200 10836 13252
rect 14740 13336 14792 13388
rect 15108 13336 15160 13388
rect 14004 13268 14056 13320
rect 14188 13268 14240 13320
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 20168 13336 20220 13388
rect 27988 13404 28040 13456
rect 22928 13336 22980 13388
rect 24584 13379 24636 13388
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 15660 13268 15712 13320
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 18236 13311 18288 13320
rect 18236 13277 18245 13311
rect 18245 13277 18279 13311
rect 18279 13277 18288 13311
rect 18236 13268 18288 13277
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 19340 13268 19392 13320
rect 19524 13268 19576 13320
rect 21088 13268 21140 13320
rect 22744 13311 22796 13320
rect 9772 13132 9824 13184
rect 10140 13132 10192 13184
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 13452 13132 13504 13184
rect 15476 13132 15528 13184
rect 16396 13243 16448 13252
rect 16396 13209 16405 13243
rect 16405 13209 16439 13243
rect 16439 13209 16448 13243
rect 16396 13200 16448 13209
rect 16672 13200 16724 13252
rect 17040 13200 17092 13252
rect 19064 13200 19116 13252
rect 22744 13277 22753 13311
rect 22753 13277 22787 13311
rect 22787 13277 22796 13311
rect 22744 13268 22796 13277
rect 25228 13268 25280 13320
rect 23756 13200 23808 13252
rect 23940 13243 23992 13252
rect 23940 13209 23949 13243
rect 23949 13209 23983 13243
rect 23983 13209 23992 13243
rect 23940 13200 23992 13209
rect 25596 13268 25648 13320
rect 25780 13200 25832 13252
rect 16856 13132 16908 13184
rect 24768 13132 24820 13184
rect 25320 13132 25372 13184
rect 27252 13132 27304 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3700 12928 3752 12980
rect 6092 12928 6144 12980
rect 8392 12928 8444 12980
rect 10324 12928 10376 12980
rect 11336 12928 11388 12980
rect 1860 12903 1912 12912
rect 1860 12869 1869 12903
rect 1869 12869 1903 12903
rect 1903 12869 1912 12903
rect 1860 12860 1912 12869
rect 4344 12903 4396 12912
rect 4344 12869 4353 12903
rect 4353 12869 4387 12903
rect 4387 12869 4396 12903
rect 4344 12860 4396 12869
rect 6736 12860 6788 12912
rect 6920 12860 6972 12912
rect 7840 12860 7892 12912
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 5448 12792 5500 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 1584 12767 1636 12776
rect 1584 12733 1593 12767
rect 1593 12733 1627 12767
rect 1627 12733 1636 12767
rect 1584 12724 1636 12733
rect 2228 12724 2280 12776
rect 3792 12724 3844 12776
rect 6184 12724 6236 12776
rect 5816 12699 5868 12708
rect 5816 12665 5825 12699
rect 5825 12665 5859 12699
rect 5859 12665 5868 12699
rect 7380 12724 7432 12776
rect 7564 12724 7616 12776
rect 9496 12792 9548 12844
rect 10048 12792 10100 12844
rect 16212 12928 16264 12980
rect 16488 12928 16540 12980
rect 18328 12928 18380 12980
rect 19064 12971 19116 12980
rect 19064 12937 19073 12971
rect 19073 12937 19107 12971
rect 19107 12937 19116 12971
rect 19064 12928 19116 12937
rect 19984 12928 20036 12980
rect 20812 12928 20864 12980
rect 22284 12928 22336 12980
rect 13636 12860 13688 12912
rect 15200 12860 15252 12912
rect 20168 12860 20220 12912
rect 23572 12928 23624 12980
rect 24216 12971 24268 12980
rect 24216 12937 24225 12971
rect 24225 12937 24259 12971
rect 24259 12937 24268 12971
rect 24216 12928 24268 12937
rect 25596 12971 25648 12980
rect 25596 12937 25605 12971
rect 25605 12937 25639 12971
rect 25639 12937 25648 12971
rect 25596 12928 25648 12937
rect 23112 12903 23164 12912
rect 23112 12869 23121 12903
rect 23121 12869 23155 12903
rect 23155 12869 23164 12903
rect 23112 12860 23164 12869
rect 8116 12724 8168 12776
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 9312 12724 9364 12776
rect 11152 12724 11204 12776
rect 15936 12792 15988 12844
rect 18144 12792 18196 12844
rect 18512 12792 18564 12844
rect 21364 12792 21416 12844
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 24768 12792 24820 12844
rect 25412 12792 25464 12844
rect 26240 12792 26292 12844
rect 38016 12835 38068 12844
rect 38016 12801 38025 12835
rect 38025 12801 38059 12835
rect 38059 12801 38068 12835
rect 38016 12792 38068 12801
rect 5816 12656 5868 12665
rect 6184 12588 6236 12640
rect 7932 12588 7984 12640
rect 8116 12588 8168 12640
rect 8576 12588 8628 12640
rect 9772 12588 9824 12640
rect 10784 12588 10836 12640
rect 11612 12588 11664 12640
rect 12164 12588 12216 12640
rect 15200 12724 15252 12776
rect 15568 12767 15620 12776
rect 15568 12733 15577 12767
rect 15577 12733 15611 12767
rect 15611 12733 15620 12767
rect 15568 12724 15620 12733
rect 16764 12724 16816 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 23940 12724 23992 12776
rect 28264 12724 28316 12776
rect 13728 12656 13780 12708
rect 15016 12656 15068 12708
rect 25320 12656 25372 12708
rect 13084 12588 13136 12640
rect 16212 12588 16264 12640
rect 21180 12588 21232 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 2136 12384 2188 12436
rect 3424 12427 3476 12436
rect 2044 12248 2096 12300
rect 3148 12248 3200 12300
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 7472 12384 7524 12436
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 3608 12248 3660 12300
rect 3884 12044 3936 12096
rect 5540 12248 5592 12300
rect 6552 12248 6604 12300
rect 6828 12248 6880 12300
rect 10692 12384 10744 12436
rect 8116 12316 8168 12368
rect 9036 12316 9088 12368
rect 10600 12316 10652 12368
rect 16488 12384 16540 12436
rect 16580 12384 16632 12436
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 11428 12316 11480 12368
rect 12532 12316 12584 12368
rect 12716 12316 12768 12368
rect 16948 12316 17000 12368
rect 17316 12316 17368 12368
rect 7840 12248 7892 12300
rect 8392 12248 8444 12300
rect 7196 12180 7248 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 4620 12112 4672 12164
rect 6276 12112 6328 12164
rect 9496 12180 9548 12232
rect 10508 12248 10560 12300
rect 14740 12248 14792 12300
rect 8668 12112 8720 12164
rect 10048 12112 10100 12164
rect 12348 12180 12400 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 16028 12180 16080 12232
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 17500 12180 17552 12232
rect 21088 12384 21140 12436
rect 23112 12384 23164 12436
rect 23756 12384 23808 12436
rect 24860 12384 24912 12436
rect 19340 12248 19392 12300
rect 20352 12316 20404 12368
rect 20076 12248 20128 12300
rect 33968 12316 34020 12368
rect 19984 12180 20036 12232
rect 20628 12180 20680 12232
rect 22652 12180 22704 12232
rect 23204 12180 23256 12232
rect 25412 12223 25464 12232
rect 11152 12112 11204 12164
rect 12900 12112 12952 12164
rect 11612 12044 11664 12096
rect 12992 12044 13044 12096
rect 13820 12044 13872 12096
rect 14556 12112 14608 12164
rect 15016 12155 15068 12164
rect 15016 12121 15025 12155
rect 15025 12121 15059 12155
rect 15059 12121 15068 12155
rect 15016 12112 15068 12121
rect 16488 12112 16540 12164
rect 20904 12112 20956 12164
rect 20996 12155 21048 12164
rect 20996 12121 21005 12155
rect 21005 12121 21039 12155
rect 21039 12121 21048 12155
rect 21548 12155 21600 12164
rect 20996 12112 21048 12121
rect 21548 12121 21557 12155
rect 21557 12121 21591 12155
rect 21591 12121 21600 12155
rect 21548 12112 21600 12121
rect 19248 12044 19300 12096
rect 19432 12044 19484 12096
rect 25412 12189 25421 12223
rect 25421 12189 25455 12223
rect 25455 12189 25464 12223
rect 25412 12180 25464 12189
rect 38108 12180 38160 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 3516 11840 3568 11892
rect 7012 11840 7064 11892
rect 9312 11840 9364 11892
rect 9496 11840 9548 11892
rect 10324 11840 10376 11892
rect 11428 11840 11480 11892
rect 4620 11815 4672 11824
rect 4620 11781 4629 11815
rect 4629 11781 4663 11815
rect 4663 11781 4672 11815
rect 4620 11772 4672 11781
rect 1492 11704 1544 11756
rect 3976 11704 4028 11756
rect 7012 11704 7064 11756
rect 7932 11772 7984 11824
rect 9036 11772 9088 11824
rect 9404 11772 9456 11824
rect 12440 11772 12492 11824
rect 14096 11840 14148 11892
rect 14924 11840 14976 11892
rect 15292 11883 15344 11892
rect 15292 11849 15301 11883
rect 15301 11849 15335 11883
rect 15335 11849 15344 11883
rect 15292 11840 15344 11849
rect 16120 11883 16172 11892
rect 16120 11849 16129 11883
rect 16129 11849 16163 11883
rect 16163 11849 16172 11883
rect 16120 11840 16172 11849
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 18420 11840 18472 11892
rect 19340 11840 19392 11892
rect 20628 11840 20680 11892
rect 20996 11840 21048 11892
rect 15384 11772 15436 11824
rect 15476 11772 15528 11824
rect 10692 11704 10744 11756
rect 12532 11704 12584 11756
rect 1860 11679 1912 11688
rect 1860 11645 1869 11679
rect 1869 11645 1903 11679
rect 1903 11645 1912 11679
rect 1860 11636 1912 11645
rect 5172 11679 5224 11688
rect 1676 11568 1728 11620
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 5172 11500 5224 11552
rect 5632 11500 5684 11552
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 6736 11636 6788 11688
rect 8668 11636 8720 11688
rect 9220 11568 9272 11620
rect 10048 11636 10100 11688
rect 10416 11636 10468 11688
rect 11336 11636 11388 11688
rect 12900 11636 12952 11688
rect 10232 11568 10284 11620
rect 10324 11568 10376 11620
rect 15108 11704 15160 11756
rect 10048 11500 10100 11552
rect 14648 11500 14700 11552
rect 15660 11568 15712 11620
rect 17316 11568 17368 11620
rect 17592 11704 17644 11756
rect 19984 11772 20036 11824
rect 20720 11772 20772 11824
rect 19432 11704 19484 11756
rect 20628 11747 20680 11756
rect 20628 11713 20637 11747
rect 20637 11713 20671 11747
rect 20671 11713 20680 11747
rect 20628 11704 20680 11713
rect 20904 11704 20956 11756
rect 18144 11636 18196 11688
rect 19248 11636 19300 11688
rect 20996 11636 21048 11688
rect 18788 11500 18840 11552
rect 20628 11500 20680 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1952 11296 2004 11348
rect 9404 11296 9456 11348
rect 11888 11296 11940 11348
rect 12256 11296 12308 11348
rect 13912 11296 13964 11348
rect 16396 11296 16448 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 20812 11296 20864 11348
rect 7748 11228 7800 11280
rect 4620 11160 4672 11212
rect 5540 11160 5592 11212
rect 5816 11160 5868 11212
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 3700 11092 3752 11144
rect 2044 11024 2096 11076
rect 2412 11024 2464 11076
rect 5172 11067 5224 11076
rect 5172 11033 5181 11067
rect 5181 11033 5215 11067
rect 5215 11033 5224 11067
rect 5172 11024 5224 11033
rect 6184 11024 6236 11076
rect 7656 11160 7708 11212
rect 8300 11228 8352 11280
rect 8668 11228 8720 11280
rect 9496 11228 9548 11280
rect 10508 11228 10560 11280
rect 12164 11228 12216 11280
rect 7104 11092 7156 11144
rect 9220 11160 9272 11212
rect 12256 11160 12308 11212
rect 8300 11092 8352 11144
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9864 11092 9916 11144
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 8484 11067 8536 11076
rect 8484 11033 8493 11067
rect 8493 11033 8527 11067
rect 8527 11033 8536 11067
rect 8484 11024 8536 11033
rect 8576 11024 8628 11076
rect 11612 11092 11664 11144
rect 12992 11228 13044 11280
rect 21364 11228 21416 11280
rect 22468 11296 22520 11348
rect 37188 11296 37240 11348
rect 14648 11092 14700 11144
rect 18144 11203 18196 11212
rect 18144 11169 18153 11203
rect 18153 11169 18187 11203
rect 18187 11169 18196 11203
rect 18144 11160 18196 11169
rect 21732 11160 21784 11212
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 17960 11092 18012 11144
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 38292 11135 38344 11144
rect 5908 10956 5960 11008
rect 6552 10956 6604 11008
rect 7472 10956 7524 11008
rect 10508 10956 10560 11008
rect 15752 10956 15804 11008
rect 17500 10999 17552 11008
rect 17500 10965 17509 10999
rect 17509 10965 17543 10999
rect 17543 10965 17552 10999
rect 17500 10956 17552 10965
rect 19432 10956 19484 11008
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 21364 11067 21416 11076
rect 21364 11033 21373 11067
rect 21373 11033 21407 11067
rect 21407 11033 21416 11067
rect 21364 11024 21416 11033
rect 21456 11067 21508 11076
rect 21456 11033 21465 11067
rect 21465 11033 21499 11067
rect 21499 11033 21508 11067
rect 21456 11024 21508 11033
rect 21732 11024 21784 11076
rect 28356 11024 28408 11076
rect 22744 10956 22796 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1952 10752 2004 10804
rect 2780 10752 2832 10804
rect 2964 10752 3016 10804
rect 3424 10752 3476 10804
rect 4160 10752 4212 10804
rect 4988 10752 5040 10804
rect 5356 10752 5408 10804
rect 7564 10795 7616 10804
rect 7564 10761 7573 10795
rect 7573 10761 7607 10795
rect 7607 10761 7616 10795
rect 7564 10752 7616 10761
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2688 10616 2740 10668
rect 3148 10616 3200 10668
rect 10416 10752 10468 10804
rect 13176 10752 13228 10804
rect 14004 10752 14056 10804
rect 15200 10752 15252 10804
rect 15936 10795 15988 10804
rect 15936 10761 15945 10795
rect 15945 10761 15979 10795
rect 15979 10761 15988 10795
rect 15936 10752 15988 10761
rect 16764 10752 16816 10804
rect 19432 10752 19484 10804
rect 21456 10752 21508 10804
rect 21548 10752 21600 10804
rect 8576 10684 8628 10736
rect 6000 10659 6052 10668
rect 6000 10625 6009 10659
rect 6009 10625 6043 10659
rect 6043 10625 6052 10659
rect 6000 10616 6052 10625
rect 7012 10616 7064 10668
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 8944 10659 8996 10668
rect 2320 10480 2372 10532
rect 3424 10480 3476 10532
rect 7380 10548 7432 10600
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9772 10684 9824 10736
rect 9956 10684 10008 10736
rect 12256 10727 12308 10736
rect 12256 10693 12265 10727
rect 12265 10693 12299 10727
rect 12299 10693 12308 10727
rect 12256 10684 12308 10693
rect 12992 10684 13044 10736
rect 17868 10684 17920 10736
rect 13268 10616 13320 10668
rect 14648 10659 14700 10668
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 15568 10616 15620 10668
rect 17500 10616 17552 10668
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 19524 10659 19576 10668
rect 8392 10480 8444 10532
rect 11704 10548 11756 10600
rect 12532 10548 12584 10600
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 20536 10616 20588 10668
rect 21640 10616 21692 10668
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 27252 10659 27304 10668
rect 27252 10625 27261 10659
rect 27261 10625 27295 10659
rect 27295 10625 27304 10659
rect 27252 10616 27304 10625
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 13084 10480 13136 10532
rect 18512 10480 18564 10532
rect 34152 10480 34204 10532
rect 2596 10412 2648 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 8852 10412 8904 10464
rect 10876 10412 10928 10464
rect 18696 10412 18748 10464
rect 23572 10412 23624 10464
rect 36360 10412 36412 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1308 10208 1360 10260
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3700 10208 3752 10260
rect 6552 10208 6604 10260
rect 8024 10208 8076 10260
rect 8116 10208 8168 10260
rect 3792 10140 3844 10192
rect 7472 10140 7524 10192
rect 9956 10208 10008 10260
rect 10784 10208 10836 10260
rect 8576 10140 8628 10192
rect 9128 10140 9180 10192
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 5908 10072 5960 10124
rect 6276 10072 6328 10124
rect 6920 10072 6972 10124
rect 11980 10208 12032 10260
rect 12716 10208 12768 10260
rect 14464 10208 14516 10260
rect 15568 10251 15620 10260
rect 9588 10072 9640 10124
rect 14648 10140 14700 10192
rect 2688 10004 2740 10056
rect 3148 10004 3200 10056
rect 3608 10004 3660 10056
rect 7380 10004 7432 10056
rect 8300 10004 8352 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 4528 9936 4580 9988
rect 4804 9936 4856 9988
rect 5632 9936 5684 9988
rect 2044 9868 2096 9920
rect 6736 9868 6788 9920
rect 9588 9936 9640 9988
rect 10876 10004 10928 10056
rect 12716 10072 12768 10124
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 18328 10208 18380 10260
rect 18604 10208 18656 10260
rect 20536 10251 20588 10260
rect 20536 10217 20545 10251
rect 20545 10217 20579 10251
rect 20579 10217 20588 10251
rect 20536 10208 20588 10217
rect 33968 10251 34020 10260
rect 33968 10217 33977 10251
rect 33977 10217 34011 10251
rect 34011 10217 34020 10251
rect 33968 10208 34020 10217
rect 16212 10140 16264 10192
rect 17960 10072 18012 10124
rect 15108 10047 15160 10056
rect 10784 9868 10836 9920
rect 11428 9936 11480 9988
rect 12532 9936 12584 9988
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 17224 10004 17276 10056
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 19524 10004 19576 10056
rect 28264 10047 28316 10056
rect 28264 10013 28273 10047
rect 28273 10013 28307 10047
rect 28307 10013 28316 10047
rect 28264 10004 28316 10013
rect 28356 10004 28408 10056
rect 37188 10004 37240 10056
rect 14464 9868 14516 9920
rect 18512 9868 18564 9920
rect 29644 9868 29696 9920
rect 31668 9868 31720 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2596 9664 2648 9716
rect 1216 9596 1268 9648
rect 2504 9639 2556 9648
rect 2504 9605 2513 9639
rect 2513 9605 2547 9639
rect 2547 9605 2556 9639
rect 2504 9596 2556 9605
rect 1952 9528 2004 9580
rect 2596 9528 2648 9580
rect 3608 9596 3660 9648
rect 4804 9664 4856 9716
rect 5448 9664 5500 9716
rect 5540 9664 5592 9716
rect 7012 9664 7064 9716
rect 8116 9664 8168 9716
rect 8300 9664 8352 9716
rect 8944 9664 8996 9716
rect 1584 9324 1636 9376
rect 2596 9324 2648 9376
rect 3700 9460 3752 9512
rect 5264 9528 5316 9580
rect 6092 9528 6144 9580
rect 6920 9596 6972 9648
rect 8392 9596 8444 9648
rect 8760 9596 8812 9648
rect 11060 9639 11112 9648
rect 5448 9460 5500 9512
rect 5172 9392 5224 9444
rect 3792 9324 3844 9376
rect 5816 9324 5868 9376
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7564 9460 7616 9512
rect 7932 9392 7984 9444
rect 9404 9528 9456 9580
rect 10140 9528 10192 9580
rect 11060 9605 11069 9639
rect 11069 9605 11103 9639
rect 11103 9605 11112 9639
rect 11060 9596 11112 9605
rect 10876 9528 10928 9580
rect 12256 9596 12308 9648
rect 12808 9596 12860 9648
rect 14556 9639 14608 9648
rect 14556 9605 14565 9639
rect 14565 9605 14599 9639
rect 14599 9605 14608 9639
rect 14556 9596 14608 9605
rect 8760 9460 8812 9512
rect 8576 9392 8628 9444
rect 8760 9324 8812 9376
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 10784 9460 10836 9512
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 12440 9528 12492 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 14096 9460 14148 9512
rect 31668 9528 31720 9580
rect 12072 9392 12124 9444
rect 25228 9460 25280 9512
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 16580 9324 16632 9376
rect 38016 9324 38068 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3424 9120 3476 9172
rect 7104 9163 7156 9172
rect 3516 9052 3568 9104
rect 2228 8984 2280 9036
rect 2596 8984 2648 9036
rect 4620 8984 4672 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2504 8848 2556 8900
rect 5632 8848 5684 8900
rect 6368 8891 6420 8900
rect 6368 8857 6377 8891
rect 6377 8857 6411 8891
rect 6411 8857 6420 8891
rect 6368 8848 6420 8857
rect 7104 9129 7134 9163
rect 7134 9129 7156 9163
rect 7104 9120 7156 9129
rect 8116 9120 8168 9172
rect 8300 9052 8352 9104
rect 9496 9120 9548 9172
rect 9772 9120 9824 9172
rect 12624 9163 12676 9172
rect 10140 9052 10192 9104
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 14004 9120 14056 9172
rect 20260 9120 20312 9172
rect 13268 9052 13320 9104
rect 14188 9052 14240 9104
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7564 8984 7616 9036
rect 8944 8984 8996 9036
rect 9036 8916 9088 8968
rect 10968 8984 11020 9036
rect 11060 8984 11112 9036
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 17960 8984 18012 9036
rect 12808 8916 12860 8968
rect 13176 8916 13228 8968
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 6828 8780 6880 8832
rect 7012 8780 7064 8832
rect 8484 8780 8536 8832
rect 10876 8848 10928 8900
rect 11244 8848 11296 8900
rect 28632 8916 28684 8968
rect 38016 8959 38068 8968
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 12532 8780 12584 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 4896 8576 4948 8628
rect 5080 8576 5132 8628
rect 5724 8576 5776 8628
rect 6368 8576 6420 8628
rect 1860 8440 1912 8492
rect 2044 8440 2096 8492
rect 3608 8440 3660 8492
rect 3792 8440 3844 8492
rect 5080 8440 5132 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 1584 8304 1636 8356
rect 3700 8372 3752 8424
rect 8024 8508 8076 8560
rect 8484 8508 8536 8560
rect 9312 8576 9364 8628
rect 10232 8576 10284 8628
rect 11152 8576 11204 8628
rect 11520 8576 11572 8628
rect 12348 8619 12400 8628
rect 12348 8585 12357 8619
rect 12357 8585 12391 8619
rect 12391 8585 12400 8619
rect 12348 8576 12400 8585
rect 12992 8619 13044 8628
rect 12992 8585 13001 8619
rect 13001 8585 13035 8619
rect 13035 8585 13044 8619
rect 12992 8576 13044 8585
rect 14096 8576 14148 8628
rect 14740 8619 14792 8628
rect 14740 8585 14749 8619
rect 14749 8585 14783 8619
rect 14783 8585 14792 8619
rect 14740 8576 14792 8585
rect 14832 8576 14884 8628
rect 25412 8576 25464 8628
rect 17316 8508 17368 8560
rect 17500 8508 17552 8560
rect 22560 8508 22612 8560
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 10784 8440 10836 8492
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13176 8483 13228 8492
rect 13176 8449 13185 8483
rect 13185 8449 13219 8483
rect 13219 8449 13228 8483
rect 13176 8440 13228 8449
rect 13268 8440 13320 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 2320 8236 2372 8288
rect 2688 8236 2740 8288
rect 6920 8372 6972 8424
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8024 8372 8076 8424
rect 14832 8372 14884 8424
rect 7104 8347 7156 8356
rect 7104 8313 7113 8347
rect 7113 8313 7147 8347
rect 7147 8313 7156 8347
rect 7104 8304 7156 8313
rect 9312 8304 9364 8356
rect 11704 8304 11756 8356
rect 8116 8236 8168 8288
rect 8484 8236 8536 8288
rect 10140 8236 10192 8288
rect 13360 8304 13412 8356
rect 17040 8304 17092 8356
rect 22008 8440 22060 8492
rect 33968 8483 34020 8492
rect 33968 8449 33977 8483
rect 33977 8449 34011 8483
rect 34011 8449 34020 8483
rect 33968 8440 34020 8449
rect 22468 8372 22520 8424
rect 21180 8304 21232 8356
rect 22376 8304 22428 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 4804 8032 4856 8084
rect 5724 8032 5776 8084
rect 7932 8075 7984 8084
rect 3332 8007 3384 8016
rect 3332 7973 3341 8007
rect 3341 7973 3375 8007
rect 3375 7973 3384 8007
rect 3332 7964 3384 7973
rect 4988 7964 5040 8016
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 10600 8032 10652 8084
rect 12900 8032 12952 8084
rect 13176 8032 13228 8084
rect 27988 8075 28040 8084
rect 27988 8041 27997 8075
rect 27997 8041 28031 8075
rect 28031 8041 28040 8075
rect 27988 8032 28040 8041
rect 37188 8032 37240 8084
rect 10048 7964 10100 8016
rect 11704 7964 11756 8016
rect 3148 7896 3200 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 3700 7828 3752 7880
rect 6920 7896 6972 7948
rect 10600 7896 10652 7948
rect 11796 7896 11848 7948
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 2872 7760 2924 7812
rect 4068 7760 4120 7812
rect 5448 7692 5500 7744
rect 6552 7760 6604 7812
rect 10508 7760 10560 7812
rect 10876 7760 10928 7812
rect 8300 7692 8352 7744
rect 9956 7692 10008 7744
rect 33600 7828 33652 7880
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 15108 7760 15160 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4712 7488 4764 7540
rect 5724 7488 5776 7540
rect 6460 7488 6512 7540
rect 1952 7463 2004 7472
rect 1952 7429 1961 7463
rect 1961 7429 1995 7463
rect 1995 7429 2004 7463
rect 1952 7420 2004 7429
rect 2964 7420 3016 7472
rect 3884 7420 3936 7472
rect 1584 7352 1636 7404
rect 3148 7284 3200 7336
rect 5080 7352 5132 7404
rect 6460 7352 6512 7404
rect 6920 7352 6972 7404
rect 7748 7420 7800 7472
rect 8484 7420 8536 7472
rect 10048 7488 10100 7540
rect 10324 7488 10376 7540
rect 9956 7420 10008 7472
rect 11796 7488 11848 7540
rect 11152 7420 11204 7472
rect 7564 7284 7616 7336
rect 15844 7352 15896 7404
rect 36360 7395 36412 7404
rect 36360 7361 36369 7395
rect 36369 7361 36403 7395
rect 36403 7361 36412 7395
rect 36360 7352 36412 7361
rect 10968 7284 11020 7336
rect 4804 7216 4856 7268
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 10784 7148 10836 7200
rect 15660 7148 15712 7200
rect 17868 7148 17920 7200
rect 38016 7148 38068 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1952 6944 2004 6996
rect 1860 6876 1912 6928
rect 2412 6876 2464 6928
rect 1492 6808 1544 6860
rect 3792 6944 3844 6996
rect 5356 6944 5408 6996
rect 8944 6944 8996 6996
rect 14464 6944 14516 6996
rect 4620 6876 4672 6928
rect 1952 6740 2004 6792
rect 2044 6740 2096 6792
rect 3240 6808 3292 6860
rect 3056 6740 3108 6792
rect 3516 6740 3568 6792
rect 5724 6808 5776 6860
rect 6000 6851 6052 6860
rect 6000 6817 6009 6851
rect 6009 6817 6043 6851
rect 6043 6817 6052 6851
rect 6000 6808 6052 6817
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 6828 6808 6880 6860
rect 9036 6876 9088 6928
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 6092 6740 6144 6792
rect 6460 6740 6512 6792
rect 6736 6740 6788 6792
rect 9128 6740 9180 6792
rect 9864 6808 9916 6860
rect 9404 6740 9456 6792
rect 10048 6808 10100 6860
rect 11888 6808 11940 6860
rect 12532 6851 12584 6860
rect 12532 6817 12541 6851
rect 12541 6817 12575 6851
rect 12575 6817 12584 6851
rect 12532 6808 12584 6817
rect 25412 6851 25464 6860
rect 25412 6817 25421 6851
rect 25421 6817 25455 6851
rect 25455 6817 25464 6851
rect 25412 6808 25464 6817
rect 2228 6604 2280 6656
rect 3240 6604 3292 6656
rect 4804 6604 4856 6656
rect 5448 6604 5500 6656
rect 5724 6604 5776 6656
rect 7196 6604 7248 6656
rect 9036 6604 9088 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 11060 6672 11112 6724
rect 12348 6672 12400 6724
rect 9128 6604 9180 6613
rect 11980 6604 12032 6656
rect 12164 6604 12216 6656
rect 27528 6740 27580 6792
rect 34152 6783 34204 6792
rect 34152 6749 34161 6783
rect 34161 6749 34195 6783
rect 34195 6749 34204 6783
rect 34152 6740 34204 6749
rect 37004 6604 37056 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2136 6400 2188 6452
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 2228 6332 2280 6384
rect 5908 6400 5960 6452
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3148 6264 3200 6316
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 5724 6332 5776 6384
rect 7932 6400 7984 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 8668 6332 8720 6384
rect 4620 6307 4672 6316
rect 3700 6264 3752 6273
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 5264 6307 5316 6316
rect 4620 6264 4672 6273
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 6460 6264 6512 6316
rect 7196 6264 7248 6316
rect 4712 6196 4764 6248
rect 5080 6196 5132 6248
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 5448 6196 5500 6248
rect 7932 6264 7984 6316
rect 10048 6400 10100 6452
rect 9220 6332 9272 6384
rect 9680 6196 9732 6248
rect 4620 6128 4672 6180
rect 8944 6128 8996 6180
rect 4988 6060 5040 6112
rect 5724 6060 5776 6112
rect 7932 6060 7984 6112
rect 8300 6060 8352 6112
rect 11428 6400 11480 6452
rect 13452 6400 13504 6452
rect 18236 6400 18288 6452
rect 21272 6400 21324 6452
rect 38108 6443 38160 6452
rect 38108 6409 38117 6443
rect 38117 6409 38151 6443
rect 38151 6409 38160 6443
rect 38108 6400 38160 6409
rect 14924 6264 14976 6316
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 22652 6264 22704 6316
rect 32864 6264 32916 6316
rect 35624 6264 35676 6316
rect 38292 6307 38344 6316
rect 38292 6273 38301 6307
rect 38301 6273 38335 6307
rect 38335 6273 38344 6307
rect 38292 6264 38344 6273
rect 18420 6196 18472 6248
rect 24676 6128 24728 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2596 5856 2648 5908
rect 3976 5856 4028 5908
rect 4160 5856 4212 5908
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 7288 5856 7340 5908
rect 2964 5788 3016 5840
rect 6276 5788 6328 5840
rect 9220 5856 9272 5908
rect 10692 5856 10744 5908
rect 2504 5720 2556 5772
rect 2044 5652 2096 5704
rect 2412 5652 2464 5704
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 4252 5652 4304 5704
rect 5356 5652 5408 5704
rect 6000 5720 6052 5772
rect 11336 5788 11388 5840
rect 7472 5720 7524 5772
rect 6092 5652 6144 5704
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 11152 5695 11204 5704
rect 5724 5584 5776 5636
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 13728 5652 13780 5704
rect 17868 5695 17920 5704
rect 17868 5661 17877 5695
rect 17877 5661 17911 5695
rect 17911 5661 17920 5695
rect 17868 5652 17920 5661
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 21180 5695 21232 5704
rect 21180 5661 21189 5695
rect 21189 5661 21223 5695
rect 21223 5661 21232 5695
rect 21180 5652 21232 5661
rect 23572 5695 23624 5704
rect 23572 5661 23581 5695
rect 23581 5661 23615 5695
rect 23615 5661 23624 5695
rect 23572 5652 23624 5661
rect 10048 5584 10100 5636
rect 6184 5516 6236 5568
rect 6460 5516 6512 5568
rect 7748 5516 7800 5568
rect 18144 5516 18196 5568
rect 19432 5516 19484 5568
rect 23296 5516 23348 5568
rect 24768 5516 24820 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2320 5312 2372 5364
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 7104 5312 7156 5364
rect 5632 5244 5684 5296
rect 2412 5176 2464 5228
rect 2964 5219 3016 5228
rect 2964 5185 2973 5219
rect 2973 5185 3007 5219
rect 3007 5185 3016 5219
rect 2964 5176 3016 5185
rect 3516 5176 3568 5228
rect 3700 5176 3752 5228
rect 4252 5219 4304 5228
rect 4252 5185 4269 5219
rect 4269 5185 4303 5219
rect 4303 5185 4304 5219
rect 4252 5176 4304 5185
rect 4804 5176 4856 5228
rect 5080 5176 5132 5228
rect 7748 5176 7800 5228
rect 8208 5176 8260 5228
rect 29644 5176 29696 5228
rect 2412 5040 2464 5092
rect 4252 5040 4304 5092
rect 13084 5108 13136 5160
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 3884 4972 3936 5024
rect 4988 4972 5040 5024
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 11244 5040 11296 5092
rect 8852 4972 8904 5024
rect 9128 4972 9180 5024
rect 36912 4972 36964 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2872 4768 2924 4820
rect 3884 4700 3936 4752
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 2964 4632 3016 4684
rect 4712 4700 4764 4752
rect 5264 4700 5316 4752
rect 6552 4768 6604 4820
rect 7564 4768 7616 4820
rect 12808 4768 12860 4820
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 10876 4700 10928 4752
rect 2964 4496 3016 4548
rect 3700 4496 3752 4548
rect 4804 4564 4856 4616
rect 5356 4564 5408 4616
rect 5632 4564 5684 4616
rect 10968 4632 11020 4684
rect 7196 4564 7248 4616
rect 4712 4496 4764 4548
rect 22836 4564 22888 4616
rect 38016 4607 38068 4616
rect 38016 4573 38025 4607
rect 38025 4573 38059 4607
rect 38059 4573 38068 4607
rect 38016 4564 38068 4573
rect 7840 4428 7892 4480
rect 28172 4428 28224 4480
rect 38200 4471 38252 4480
rect 38200 4437 38209 4471
rect 38209 4437 38243 4471
rect 38243 4437 38252 4471
rect 38200 4428 38252 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3332 4224 3384 4276
rect 1860 4156 1912 4208
rect 2964 4156 3016 4208
rect 3884 4156 3936 4208
rect 5632 4156 5684 4208
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 4620 4088 4672 4140
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 6000 4088 6052 4140
rect 2780 4020 2832 4072
rect 3424 4020 3476 4072
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 11060 4020 11112 4072
rect 2688 3952 2740 4004
rect 3240 3952 3292 4004
rect 8116 3952 8168 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3240 3680 3292 3732
rect 5172 3680 5224 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6828 3680 6880 3732
rect 33968 3680 34020 3732
rect 3148 3612 3200 3664
rect 3976 3612 4028 3664
rect 5540 3612 5592 3664
rect 2596 3544 2648 3596
rect 2504 3476 2556 3528
rect 2872 3476 2924 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 5080 3519 5132 3528
rect 2412 3408 2464 3460
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 38292 3519 38344 3528
rect 4160 3408 4212 3460
rect 38292 3485 38301 3519
rect 38301 3485 38335 3519
rect 38335 3485 38344 3519
rect 38292 3476 38344 3485
rect 8484 3340 8536 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5172 3136 5224 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6736 3136 6788 3188
rect 35624 3136 35676 3188
rect 2964 3111 3016 3120
rect 2504 3000 2556 3052
rect 2964 3077 2973 3111
rect 2973 3077 3007 3111
rect 3007 3077 3016 3111
rect 2964 3068 3016 3077
rect 3976 3068 4028 3120
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 5172 3043 5224 3052
rect 2780 2932 2832 2984
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5356 3000 5408 3052
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 28172 3043 28224 3052
rect 28172 3009 28181 3043
rect 28181 3009 28215 3043
rect 28215 3009 28224 3043
rect 28172 3000 28224 3009
rect 15016 2932 15068 2984
rect 37004 3000 37056 3052
rect 39304 2932 39356 2984
rect 4712 2864 4764 2916
rect 20 2796 72 2848
rect 4620 2796 4672 2848
rect 7012 2796 7064 2848
rect 30196 2796 30248 2848
rect 38200 2839 38252 2848
rect 38200 2805 38209 2839
rect 38209 2805 38243 2839
rect 38243 2805 38252 2839
rect 38200 2796 38252 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2780 2592 2832 2644
rect 5448 2592 5500 2644
rect 7380 2592 7432 2644
rect 11152 2592 11204 2644
rect 14648 2592 14700 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 18328 2592 18380 2644
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 22652 2635 22704 2644
rect 22652 2601 22661 2635
rect 22661 2601 22695 2635
rect 22695 2601 22704 2635
rect 22652 2592 22704 2601
rect 28632 2592 28684 2644
rect 33600 2635 33652 2644
rect 33600 2601 33609 2635
rect 33609 2601 33643 2635
rect 33643 2601 33652 2635
rect 33600 2592 33652 2601
rect 5356 2524 5408 2576
rect 2504 2431 2556 2440
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 3884 2388 3936 2440
rect 4620 2388 4672 2440
rect 7288 2456 7340 2508
rect 27528 2524 27580 2576
rect 32864 2524 32916 2576
rect 30196 2456 30248 2508
rect 4528 2320 4580 2372
rect 7012 2388 7064 2440
rect 7104 2388 7156 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 10784 2388 10836 2440
rect 11612 2388 11664 2440
rect 13544 2388 13596 2440
rect 14832 2388 14884 2440
rect 16764 2388 16816 2440
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 21272 2388 21324 2440
rect 22560 2388 22612 2440
rect 23296 2388 23348 2440
rect 24768 2388 24820 2440
rect 27160 2388 27212 2440
rect 27068 2320 27120 2372
rect 29000 2388 29052 2440
rect 30288 2388 30340 2440
rect 33508 2388 33560 2440
rect 34796 2388 34848 2440
rect 36084 2388 36136 2440
rect 36912 2388 36964 2440
rect 1308 2252 1360 2304
rect 5816 2252 5868 2304
rect 9036 2252 9088 2304
rect 10324 2252 10376 2304
rect 18052 2252 18104 2304
rect 19340 2252 19392 2304
rect 23848 2252 23900 2304
rect 25780 2252 25832 2304
rect 31576 2252 31628 2304
rect 38016 2252 38068 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 3238 39200 3294 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 7746 39200 7802 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 15474 39200 15530 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 30286 39200 30342 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34794 39200 34850 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 39302 39200 39358 39800
rect 32 36922 60 39200
rect 1320 37126 1348 39200
rect 3146 38176 3202 38185
rect 3146 38111 3202 38120
rect 3160 37262 3188 38111
rect 3252 37262 3280 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 37726
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 1308 37120 1360 37126
rect 1308 37062 1360 37068
rect 20 36916 72 36922
rect 20 36858 72 36864
rect 1596 36650 1624 37198
rect 2320 37120 2372 37126
rect 2320 37062 2372 37068
rect 2332 36718 2360 37062
rect 2792 36825 2820 37198
rect 5632 37188 5684 37194
rect 5632 37130 5684 37136
rect 3976 37120 4028 37126
rect 3976 37062 4028 37068
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 3988 36922 4016 37062
rect 3976 36916 4028 36922
rect 3976 36858 4028 36864
rect 2778 36816 2834 36825
rect 2778 36751 2834 36760
rect 3976 36780 4028 36786
rect 3976 36722 4028 36728
rect 2320 36712 2372 36718
rect 2320 36654 2372 36660
rect 1584 36644 1636 36650
rect 1584 36586 1636 36592
rect 3988 36378 4016 36722
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 4068 36168 4120 36174
rect 4068 36110 4120 36116
rect 1768 33516 1820 33522
rect 1768 33458 1820 33464
rect 1780 33425 1808 33458
rect 1766 33416 1822 33425
rect 1766 33351 1822 33360
rect 3884 33312 3936 33318
rect 3884 33254 3936 33260
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1780 32065 1808 32370
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1768 30728 1820 30734
rect 1766 30696 1768 30705
rect 1820 30696 1822 30705
rect 1766 30631 1822 30640
rect 1492 30592 1544 30598
rect 1492 30534 1544 30540
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1216 18624 1268 18630
rect 1216 18566 1268 18572
rect 1228 9654 1256 18566
rect 1320 10266 1348 21626
rect 1504 17270 1532 30534
rect 3896 29646 3924 33254
rect 3976 32224 4028 32230
rect 3976 32166 4028 32172
rect 3884 29640 3936 29646
rect 3884 29582 3936 29588
rect 1768 29164 1820 29170
rect 1768 29106 1820 29112
rect 1780 28665 1808 29106
rect 1766 28656 1822 28665
rect 1766 28591 1822 28600
rect 3988 28082 4016 32166
rect 3976 28076 4028 28082
rect 3976 28018 4028 28024
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 27305 1808 27406
rect 1766 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 25288 1820 25294
rect 1766 25256 1768 25265
rect 1820 25256 1822 25265
rect 1766 25191 1822 25200
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 1596 23866 1624 24142
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1952 24064 2004 24070
rect 1952 24006 2004 24012
rect 1780 23905 1808 24006
rect 1766 23896 1822 23905
rect 1584 23860 1636 23866
rect 1766 23831 1822 23840
rect 1584 23802 1636 23808
rect 1964 23730 1992 24006
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1584 22568 1636 22574
rect 1584 22510 1636 22516
rect 1596 22030 1624 22510
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1596 21486 1624 21966
rect 1584 21480 1636 21486
rect 1584 21422 1636 21428
rect 1596 20942 1624 21422
rect 1584 20936 1636 20942
rect 1584 20878 1636 20884
rect 1596 20398 1624 20878
rect 1584 20392 1636 20398
rect 1584 20334 1636 20340
rect 1596 19854 1624 20334
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19310 1624 19790
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1596 18766 1624 19246
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1492 17264 1544 17270
rect 1492 17206 1544 17212
rect 1596 17066 1624 18702
rect 1688 17202 1716 22918
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1780 20505 1808 21490
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1780 18426 1808 19071
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1584 17060 1636 17066
rect 1584 17002 1636 17008
rect 1596 16590 1624 17002
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1596 16046 1624 16526
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 14940 1624 15982
rect 1780 15745 1808 16934
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1872 15586 1900 18634
rect 1964 17678 1992 21286
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1780 15558 1900 15586
rect 1676 14952 1728 14958
rect 1596 14912 1676 14940
rect 1676 14894 1728 14900
rect 1688 14414 1716 14894
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1504 11762 1532 13874
rect 1688 13326 1716 14350
rect 1780 13734 1808 15558
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1872 13938 1900 15438
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1858 13424 1914 13433
rect 1858 13359 1914 13368
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1584 12776 1636 12782
rect 1688 12764 1716 13262
rect 1872 12918 1900 13359
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 1636 12736 1716 12764
rect 1584 12718 1636 12724
rect 1688 12238 1716 12736
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1216 9648 1268 9654
rect 1216 9590 1268 9596
rect 1504 6866 1532 11698
rect 1688 11626 1716 12174
rect 1676 11620 1728 11626
rect 1676 11562 1728 11568
rect 1688 11150 1716 11562
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10985 1716 11086
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1688 9674 1716 10911
rect 1596 9646 1716 9674
rect 1596 9382 1624 9646
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8974 1624 9318
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8362 1624 8910
rect 1674 8664 1730 8673
rect 1674 8599 1676 8608
rect 1728 8599 1730 8608
rect 1676 8570 1728 8576
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1596 7886 1624 8298
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7410 1624 7822
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1780 6322 1808 12271
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1872 8498 1900 11630
rect 1964 11354 1992 16594
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2056 12306 2084 16186
rect 2148 15570 2176 23666
rect 2332 18193 2360 24142
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2318 18184 2374 18193
rect 2318 18119 2374 18128
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2148 12442 2176 15506
rect 2516 15178 2544 18226
rect 2608 16658 2636 23598
rect 2700 23118 2728 23666
rect 2872 23520 2924 23526
rect 2872 23462 2924 23468
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2700 21622 2728 21830
rect 2688 21616 2740 21622
rect 2688 21558 2740 21564
rect 2792 17785 2820 22918
rect 2884 20874 2912 23462
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2976 21865 3004 21898
rect 2962 21856 3018 21865
rect 2962 21791 3018 21800
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2778 17776 2834 17785
rect 2778 17711 2834 17720
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2516 15150 2636 15178
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1950 10840 2006 10849
rect 1950 10775 1952 10784
rect 2004 10775 2006 10784
rect 1952 10746 2004 10752
rect 2056 9926 2084 11018
rect 2134 10160 2190 10169
rect 2134 10095 2190 10104
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1964 8378 1992 9522
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1872 8350 1992 8378
rect 1872 6934 1900 8350
rect 1950 8256 2006 8265
rect 1950 8191 2006 8200
rect 1964 7478 1992 8191
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1860 6928 1912 6934
rect 1860 6870 1912 6876
rect 1964 6798 1992 6938
rect 2056 6798 2084 8434
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 2056 5710 2084 6734
rect 2148 6458 2176 10095
rect 2240 9042 2268 12718
rect 2332 10674 2360 13738
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2332 8294 2360 10474
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2424 7698 2452 11018
rect 2516 9654 2544 15030
rect 2608 10470 2636 15150
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2700 14482 2728 14758
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2792 11801 2820 17614
rect 2884 15570 2912 18362
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2976 14464 3004 16458
rect 3068 15570 3096 21286
rect 3160 19786 3188 23462
rect 3896 23254 3924 23666
rect 3884 23248 3936 23254
rect 3884 23190 3936 23196
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3252 20534 3280 22918
rect 3884 22704 3936 22710
rect 3884 22646 3936 22652
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 2884 14436 3004 14464
rect 2778 11792 2834 11801
rect 2778 11727 2834 11736
rect 2778 11248 2834 11257
rect 2778 11183 2834 11192
rect 2792 10810 2820 11183
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2700 10062 2728 10610
rect 2688 10056 2740 10062
rect 2608 10016 2688 10044
rect 2608 9722 2636 10016
rect 2688 9998 2740 10004
rect 2596 9716 2648 9722
rect 2884 9674 2912 14436
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2976 13841 3004 14282
rect 2962 13832 3018 13841
rect 2962 13767 3018 13776
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2976 13190 3004 13670
rect 2964 13184 3016 13190
rect 3160 13138 3188 19314
rect 3252 16046 3280 19654
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 3344 18970 3372 19246
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3238 14376 3294 14385
rect 3238 14311 3294 14320
rect 2964 13126 3016 13132
rect 3068 13110 3188 13138
rect 3068 12434 3096 13110
rect 2976 12406 3096 12434
rect 2976 10810 3004 12406
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3160 10674 3188 12242
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10062 3188 10610
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2596 9658 2648 9664
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2608 9586 2636 9658
rect 2700 9646 2912 9674
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 9042 2636 9318
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2700 8922 2728 9646
rect 2778 9480 2834 9489
rect 2778 9415 2834 9424
rect 3054 9480 3110 9489
rect 3054 9415 3110 9424
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2608 8894 2728 8922
rect 2332 7670 2452 7698
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2240 6390 2268 6598
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2332 5370 2360 7670
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2424 6322 2452 6870
rect 2516 6458 2544 8842
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2424 6066 2452 6258
rect 2424 6038 2544 6066
rect 2516 5778 2544 6038
rect 2608 5914 2636 8894
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2424 5234 2452 5646
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2424 5098 2452 5170
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4865 1808 4966
rect 1766 4856 1822 4865
rect 1766 4791 1822 4800
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1872 4214 1900 4558
rect 1860 4208 1912 4214
rect 1860 4150 1912 4156
rect 2424 3466 2452 5034
rect 2700 4010 2728 8230
rect 2792 4078 2820 9415
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 2884 4826 2912 7754
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2976 5846 3004 7414
rect 3068 6882 3096 9415
rect 3160 7954 3188 9998
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3160 7342 3188 7890
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3068 6854 3188 6882
rect 3252 6866 3280 14311
rect 3344 10266 3372 16118
rect 3528 15094 3556 22510
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3608 20868 3660 20874
rect 3608 20810 3660 20816
rect 3620 20466 3648 20810
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3606 18592 3662 18601
rect 3606 18527 3662 18536
rect 3620 18290 3648 18527
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 3712 17746 3740 21626
rect 3790 19952 3846 19961
rect 3790 19887 3792 19896
rect 3844 19887 3846 19896
rect 3792 19858 3844 19864
rect 3804 19446 3832 19858
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3606 16280 3662 16289
rect 3606 16215 3662 16224
rect 3620 16182 3648 16215
rect 3608 16176 3660 16182
rect 3608 16118 3660 16124
rect 3804 15366 3832 18158
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3516 15088 3568 15094
rect 3792 15088 3844 15094
rect 3516 15030 3568 15036
rect 3790 15056 3792 15065
rect 3844 15056 3846 15065
rect 3790 14991 3846 15000
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 13530 3464 14894
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3422 13016 3478 13025
rect 3528 13002 3556 13806
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3478 12974 3556 13002
rect 3422 12951 3478 12960
rect 3436 12442 3464 12951
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3620 12306 3648 13466
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3712 12986 3740 13194
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3804 12345 3832 12718
rect 3790 12336 3846 12345
rect 3608 12300 3660 12306
rect 3790 12271 3846 12280
rect 3608 12242 3660 12248
rect 3896 12220 3924 22646
rect 4080 22094 4108 36110
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4632 33998 4660 37062
rect 4620 33992 4672 33998
rect 4620 33934 4672 33940
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 5644 32910 5672 37130
rect 5828 37126 5856 39200
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 5816 37120 5868 37126
rect 5816 37062 5868 37068
rect 6564 34746 6592 37198
rect 7760 37126 7788 39200
rect 9048 37262 9076 39200
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 7748 37120 7800 37126
rect 7748 37062 7800 37068
rect 7852 34746 7880 37198
rect 10336 37126 10364 39200
rect 11612 37256 11664 37262
rect 11612 37198 11664 37204
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 9140 36854 9168 37062
rect 10232 36916 10284 36922
rect 10232 36858 10284 36864
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 8312 35290 8340 36722
rect 8852 36712 8904 36718
rect 8852 36654 8904 36660
rect 8300 35284 8352 35290
rect 8300 35226 8352 35232
rect 8208 35080 8260 35086
rect 8208 35022 8260 35028
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 7840 34740 7892 34746
rect 7840 34682 7892 34688
rect 5816 34604 5868 34610
rect 5816 34546 5868 34552
rect 6552 34604 6604 34610
rect 6552 34546 6604 34552
rect 5632 32904 5684 32910
rect 5632 32846 5684 32852
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5736 31793 5764 32710
rect 5722 31784 5778 31793
rect 5722 31719 5778 31728
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5828 28762 5856 34546
rect 6564 32026 6592 34546
rect 6552 32020 6604 32026
rect 6552 31962 6604 31968
rect 7380 31816 7432 31822
rect 7380 31758 7432 31764
rect 6552 29028 6604 29034
rect 6552 28970 6604 28976
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 4804 27872 4856 27878
rect 4804 27814 4856 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4172 23662 4200 24142
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4172 22642 4200 23054
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3988 22066 4108 22094
rect 3988 17728 4016 22066
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4448 21486 4476 21898
rect 4632 21570 4660 23462
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4724 22137 4752 22374
rect 4710 22128 4766 22137
rect 4710 22063 4766 22072
rect 4632 21542 4752 21570
rect 4436 21480 4488 21486
rect 4436 21422 4488 21428
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4172 20312 4200 20742
rect 4264 20466 4292 20946
rect 4526 20632 4582 20641
rect 4526 20567 4582 20576
rect 4540 20534 4568 20567
rect 4528 20528 4580 20534
rect 4528 20470 4580 20476
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4080 20284 4200 20312
rect 4080 19938 4108 20284
rect 4264 20262 4292 20402
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4080 19910 4200 19938
rect 4172 19174 4200 19910
rect 4160 19168 4212 19174
rect 4540 19156 4568 19994
rect 4632 19854 4660 21354
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4724 19310 4752 21542
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4540 19128 4660 19156
rect 4160 19110 4212 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18680 4660 19128
rect 4632 18652 4752 18680
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4436 17808 4488 17814
rect 4434 17776 4436 17785
rect 4488 17776 4490 17785
rect 3988 17700 4108 17728
rect 4434 17711 4490 17720
rect 4080 17610 4108 17700
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 3988 14414 4016 17546
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4068 16040 4120 16046
rect 4172 16028 4200 16458
rect 4120 16000 4200 16028
rect 4068 15982 4120 15988
rect 4080 15026 4108 15982
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14414 4108 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4526 14512 4582 14521
rect 4526 14447 4582 14456
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 13734 4108 14350
rect 4540 14346 4568 14447
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3976 13320 4028 13326
rect 4080 13308 4108 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4028 13280 4108 13308
rect 3976 13262 4028 13268
rect 4080 12850 4108 13280
rect 4344 12912 4396 12918
rect 4342 12880 4344 12889
rect 4396 12880 4398 12889
rect 4068 12844 4120 12850
rect 4342 12815 4398 12824
rect 4068 12786 4120 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4434 12336 4490 12345
rect 4632 12288 4660 15370
rect 4724 13870 4752 18652
rect 4816 18426 4844 27814
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5184 24818 5212 25094
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 4896 23588 4948 23594
rect 4896 23530 4948 23536
rect 4908 23186 4936 23530
rect 5000 23186 5028 24550
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 4896 23180 4948 23186
rect 4896 23122 4948 23128
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4908 20806 4936 21422
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4894 20632 4950 20641
rect 4894 20567 4950 20576
rect 4908 20058 4936 20567
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4894 19544 4950 19553
rect 4894 19479 4950 19488
rect 4908 19378 4936 19479
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 18834 4936 19110
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 5000 18698 5028 22374
rect 5092 21554 5120 24006
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5172 23112 5224 23118
rect 5172 23054 5224 23060
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19922 5120 20198
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5092 19689 5120 19722
rect 5078 19680 5134 19689
rect 5078 19615 5134 19624
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4896 18284 4948 18290
rect 4948 18244 5120 18272
rect 4896 18226 4948 18232
rect 5092 18154 5120 18244
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4816 14278 4844 17478
rect 4896 17128 4948 17134
rect 4894 17096 4896 17105
rect 4948 17096 4950 17105
rect 4894 17031 4950 17040
rect 4908 16794 4936 17031
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13530 4752 13670
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4724 13161 4752 13466
rect 4710 13152 4766 13161
rect 4710 13087 4766 13096
rect 4908 12730 4936 16458
rect 5000 16250 5028 18090
rect 5184 17814 5212 23054
rect 5368 22642 5396 23666
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 5172 17808 5224 17814
rect 5172 17750 5224 17756
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4434 12271 4490 12280
rect 3804 12192 3924 12220
rect 3974 12200 4030 12209
rect 3698 11928 3754 11937
rect 3516 11892 3568 11898
rect 3698 11863 3754 11872
rect 3516 11834 3568 11840
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3436 10538 3464 10746
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 8016 3384 8022
rect 3330 7984 3332 7993
rect 3384 7984 3386 7993
rect 3330 7919 3386 7928
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3160 6746 3188 6854
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3068 6322 3096 6734
rect 3160 6718 3372 6746
rect 3240 6656 3292 6662
rect 3146 6624 3202 6633
rect 3240 6598 3292 6604
rect 3146 6559 3202 6568
rect 3160 6458 3188 6559
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3252 6361 3280 6598
rect 3238 6352 3294 6361
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3148 6316 3200 6322
rect 3238 6287 3294 6296
rect 3148 6258 3200 6264
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 3160 5710 3188 6258
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2976 4706 3004 5170
rect 2884 4690 3004 4706
rect 2884 4684 3016 4690
rect 2884 4678 2964 4684
rect 2884 4146 2912 4678
rect 2964 4626 3016 4632
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 4214 3004 4490
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2516 3058 2544 3470
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 2516 2446 2544 2994
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1320 800 1348 2246
rect 2608 800 2636 3538
rect 2884 3534 2912 4082
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2976 3126 3004 4150
rect 3160 3670 3188 5646
rect 3344 4282 3372 6718
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3436 4078 3464 9114
rect 3528 9110 3556 11834
rect 3712 11150 3740 11863
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3712 10656 3740 11086
rect 3620 10628 3740 10656
rect 3620 10062 3648 10628
rect 3698 10568 3754 10577
rect 3698 10503 3754 10512
rect 3712 10266 3740 10503
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3804 10198 3832 12192
rect 3974 12135 4030 12144
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3620 9654 3648 9998
rect 3608 9648 3660 9654
rect 3660 9608 3832 9636
rect 3608 9590 3660 9596
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3620 8650 3648 9590
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3528 8622 3648 8650
rect 3528 6798 3556 8622
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3528 5234 3556 6734
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3620 4146 3648 8434
rect 3712 8430 3740 9454
rect 3804 9382 3832 9608
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3804 8276 3832 8434
rect 3712 8248 3832 8276
rect 3712 7886 3740 8248
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3712 6322 3740 7822
rect 3896 7478 3924 12038
rect 3988 11914 4016 12135
rect 3988 11886 4108 11914
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3804 6458 3832 6938
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3790 6216 3846 6225
rect 3790 6151 3846 6160
rect 3698 5536 3754 5545
rect 3698 5471 3754 5480
rect 3712 5370 3740 5471
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3712 4554 3740 5170
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 3738 3280 3946
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 3804 3058 3832 6151
rect 3988 5914 4016 11698
rect 4080 7818 4108 11886
rect 4448 11540 4476 12271
rect 4540 12260 4660 12288
rect 4724 12702 4936 12730
rect 4540 11937 4568 12260
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4632 12073 4660 12106
rect 4618 12064 4674 12073
rect 4618 11999 4674 12008
rect 4526 11928 4582 11937
rect 4526 11863 4582 11872
rect 4620 11824 4672 11830
rect 4618 11792 4620 11801
rect 4672 11792 4674 11801
rect 4618 11727 4674 11736
rect 4724 11540 4752 12702
rect 5000 11642 5028 15030
rect 4908 11614 5028 11642
rect 4448 11512 4660 11540
rect 4724 11512 4844 11540
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11370 4660 11512
rect 4632 11342 4752 11370
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4158 10976 4214 10985
rect 4158 10911 4214 10920
rect 4172 10810 4200 10911
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 11154
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 9489 4568 9930
rect 4526 9480 4582 9489
rect 4526 9415 4582 9424
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9042 4660 10066
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4618 7576 4674 7585
rect 4724 7546 4752 11342
rect 4816 9994 4844 11512
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4816 8090 4844 9658
rect 4908 8634 4936 11614
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 5000 9217 5028 10746
rect 4986 9208 5042 9217
rect 4986 9143 5042 9152
rect 5092 9058 5120 17206
rect 5184 14074 5212 17478
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5170 12744 5226 12753
rect 5170 12679 5226 12688
rect 5184 12434 5212 12679
rect 5276 12617 5304 20810
rect 5368 17610 5396 21626
rect 5460 20641 5488 25842
rect 5736 23730 5764 27270
rect 5816 25424 5868 25430
rect 5816 25366 5868 25372
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5446 20632 5502 20641
rect 5446 20567 5502 20576
rect 5552 20534 5580 23190
rect 5632 22092 5684 22098
rect 5828 22094 5856 25366
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 5632 22034 5684 22040
rect 5736 22066 5856 22094
rect 5908 22092 5960 22098
rect 5644 20777 5672 22034
rect 5736 21554 5764 22066
rect 5908 22034 5960 22040
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5920 21146 5948 22034
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 5630 20768 5686 20777
rect 5630 20703 5686 20712
rect 5540 20528 5592 20534
rect 5540 20470 5592 20476
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5920 20262 5948 20334
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5460 19514 5488 19858
rect 5630 19816 5686 19825
rect 5630 19751 5632 19760
rect 5684 19751 5686 19760
rect 5908 19780 5960 19786
rect 5632 19722 5684 19728
rect 5908 19722 5960 19728
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5446 19408 5502 19417
rect 5446 19343 5502 19352
rect 5460 19310 5488 19343
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5460 17542 5488 17750
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 16436 5488 17478
rect 5540 16448 5592 16454
rect 5460 16408 5540 16436
rect 5540 16390 5592 16396
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5184 12406 5304 12434
rect 5172 11688 5224 11694
rect 5170 11656 5172 11665
rect 5224 11656 5226 11665
rect 5170 11591 5226 11600
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11082 5212 11494
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5276 9674 5304 12406
rect 5368 10810 5396 16118
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5460 15162 5488 15370
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5644 14822 5672 18226
rect 5828 18154 5856 18702
rect 5816 18148 5868 18154
rect 5816 18090 5868 18096
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16182 5764 16390
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5828 14958 5856 16662
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5460 13841 5488 14282
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5446 13832 5502 13841
rect 5446 13767 5502 13776
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5460 12753 5488 12786
rect 5446 12744 5502 12753
rect 5446 12679 5502 12688
rect 5552 12424 5580 13942
rect 5460 12396 5580 12424
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5460 9722 5488 12396
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 11218 5580 12242
rect 5644 11558 5672 14758
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 9722 5580 11154
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5448 9716 5500 9722
rect 5276 9646 5396 9674
rect 5448 9658 5500 9664
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5000 9030 5120 9058
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4894 8528 4950 8537
rect 4894 8463 4950 8472
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4802 7576 4858 7585
rect 4618 7511 4674 7520
rect 4712 7540 4764 7546
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6934 4660 7511
rect 4802 7511 4858 7520
rect 4712 7482 4764 7488
rect 4816 7274 4844 7511
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4620 6928 4672 6934
rect 4158 6896 4214 6905
rect 4620 6870 4672 6876
rect 4158 6831 4214 6840
rect 4172 6202 4200 6831
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4802 6760 4858 6769
rect 4632 6322 4660 6734
rect 4802 6695 4858 6704
rect 4816 6662 4844 6695
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4080 6174 4200 6202
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4620 6180 4672 6186
rect 3976 5908 4028 5914
rect 4080 5896 4108 6174
rect 4620 6122 4672 6128
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5908 4212 5914
rect 4080 5868 4160 5896
rect 3976 5850 4028 5856
rect 4160 5850 4212 5856
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4264 5234 4292 5646
rect 4342 5400 4398 5409
rect 4342 5335 4344 5344
rect 4396 5335 4398 5344
rect 4344 5306 4396 5312
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4264 5098 4292 5170
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4758 3924 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 4250 4720 4306 4729
rect 4250 4655 4252 4664
rect 4304 4655 4306 4664
rect 4252 4626 4304 4632
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2792 2650 2820 2926
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3896 2446 3924 4150
rect 4632 4146 4660 6122
rect 4724 4758 4752 6190
rect 4908 5250 4936 8463
rect 5000 8022 5028 9030
rect 5078 8664 5134 8673
rect 5078 8599 5080 8608
rect 5132 8599 5134 8608
rect 5080 8570 5132 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4986 7440 5042 7449
rect 5092 7410 5120 8434
rect 4986 7375 5042 7384
rect 5080 7404 5132 7410
rect 5000 6118 5028 7375
rect 5080 7346 5132 7352
rect 5092 6254 5120 7346
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4986 5672 5042 5681
rect 4986 5607 5042 5616
rect 5000 5370 5028 5607
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4804 5228 4856 5234
rect 4908 5222 5028 5250
rect 4804 5170 4856 5176
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4816 4622 4844 5170
rect 5000 5030 5028 5222
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4528 4072 4580 4078
rect 4526 4040 4528 4049
rect 4580 4040 4582 4049
rect 4526 3975 4582 3984
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3988 3534 4016 3606
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3988 2825 4016 3062
rect 4172 2938 4200 3402
rect 4080 2910 4200 2938
rect 4724 2922 4752 4490
rect 5092 4146 5120 5170
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 5092 3534 5120 4082
rect 5184 3738 5212 9386
rect 5276 7886 5304 9522
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5368 7002 5396 9646
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 7750 5488 9454
rect 5644 9024 5672 9930
rect 5552 8996 5672 9024
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5446 7032 5502 7041
rect 5356 6996 5408 7002
rect 5446 6967 5502 6976
rect 5356 6938 5408 6944
rect 5460 6662 5488 6967
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5354 6488 5410 6497
rect 5354 6423 5410 6432
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5692 5304 6258
rect 5368 6254 5396 6423
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5354 5944 5410 5953
rect 5354 5879 5356 5888
rect 5408 5879 5410 5888
rect 5356 5850 5408 5856
rect 5356 5704 5408 5710
rect 5276 5664 5356 5692
rect 5356 5646 5408 5652
rect 5264 4752 5316 4758
rect 5264 4694 5316 4700
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5276 3194 5304 4694
rect 5368 4622 5396 5646
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5184 3058 5212 3130
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 4712 2916 4764 2922
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4080 1465 4108 2910
rect 4712 2858 4764 2864
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2446 4660 2790
rect 5368 2582 5396 2994
rect 5460 2650 5488 6190
rect 5552 3670 5580 8996
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 5302 5672 8842
rect 5736 8634 5764 13194
rect 5828 12714 5856 14894
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11218 5856 11494
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5920 11014 5948 19722
rect 6012 19514 6040 22374
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6104 16454 6132 22918
rect 6196 22001 6224 28494
rect 6564 26994 6592 28970
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6552 23044 6604 23050
rect 6552 22986 6604 22992
rect 6564 22658 6592 22986
rect 6656 22794 6684 23462
rect 6748 23186 6776 24006
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6656 22766 6776 22794
rect 6276 22636 6328 22642
rect 6564 22630 6684 22658
rect 6276 22578 6328 22584
rect 6182 21992 6238 22001
rect 6182 21927 6238 21936
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 21690 6224 21830
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6288 21570 6316 22578
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6196 21542 6316 21570
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6196 16046 6224 21542
rect 6380 21434 6408 22374
rect 6656 22234 6684 22630
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6550 21992 6606 22001
rect 6550 21927 6606 21936
rect 6380 21406 6500 21434
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6288 16522 6316 19314
rect 6276 16516 6328 16522
rect 6276 16458 6328 16464
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6012 10674 6040 15846
rect 6196 14890 6224 15982
rect 6288 15706 6316 16458
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6288 14618 6316 15030
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6380 13870 6408 21286
rect 6472 17746 6500 21406
rect 6564 19242 6592 21927
rect 6656 19310 6684 22170
rect 6748 22030 6776 22766
rect 6840 22166 6868 23598
rect 6932 23050 6960 24006
rect 7208 23730 7236 25230
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7208 23100 7236 23666
rect 7300 23254 7328 24754
rect 7288 23248 7340 23254
rect 7288 23190 7340 23196
rect 7392 23186 7420 31758
rect 8116 29504 8168 29510
rect 8116 29446 8168 29452
rect 8128 25362 8156 29446
rect 8116 25356 8168 25362
rect 8116 25298 8168 25304
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7576 24206 7604 24550
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 7380 23180 7432 23186
rect 7432 23140 7512 23168
rect 7380 23122 7432 23128
rect 7208 23072 7328 23100
rect 6920 23044 6972 23050
rect 6920 22986 6972 22992
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6736 21412 6788 21418
rect 6736 21354 6788 21360
rect 6748 20942 6776 21354
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20398 6776 20878
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6564 17814 6592 19178
rect 6642 18728 6698 18737
rect 6748 18698 6776 19654
rect 6642 18663 6644 18672
rect 6696 18663 6698 18672
rect 6736 18692 6788 18698
rect 6644 18634 6696 18640
rect 6736 18634 6788 18640
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6656 17746 6684 18294
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6748 16726 6776 18226
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6564 15706 6592 16050
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8498 5856 9318
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5736 7546 5764 8026
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6662 5764 6802
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5920 6458 5948 10066
rect 6104 9586 6132 12922
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 12646 6224 12718
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5998 6896 6054 6905
rect 5998 6831 6000 6840
rect 6052 6831 6054 6840
rect 6000 6802 6052 6808
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5736 6118 5764 6326
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4214 5672 4558
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 5736 3738 5764 5578
rect 6012 4146 6040 5714
rect 6104 5710 6132 6734
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6196 5574 6224 11018
rect 6288 10130 6316 12106
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6274 9888 6330 9897
rect 6274 9823 6330 9832
rect 6288 5846 6316 9823
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6380 8634 6408 8842
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6472 7546 6500 15370
rect 6748 15162 6776 15506
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6564 14958 6592 15098
rect 6552 14952 6604 14958
rect 6604 14912 6776 14940
rect 6552 14894 6604 14900
rect 6748 14414 6776 14912
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6748 13938 6776 14350
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6642 13696 6698 13705
rect 6642 13631 6698 13640
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12306 6592 12786
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10266 6592 10950
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6564 9353 6592 10202
rect 6550 9344 6606 9353
rect 6550 9279 6606 9288
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6472 6798 6500 7346
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6322 6500 6734
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6472 5574 6500 6258
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6564 4826 6592 7754
rect 6656 6866 6684 13631
rect 6748 13394 6776 13874
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6748 12918 6776 13330
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6748 11694 6776 12854
rect 6840 12306 6868 22102
rect 6932 21554 6960 22374
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 6932 18766 6960 19382
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6932 17270 6960 18566
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 7024 17082 7052 21966
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 18222 7144 21830
rect 7208 21010 7236 22578
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7208 20058 7236 20946
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7208 18329 7236 18702
rect 7194 18320 7250 18329
rect 7194 18255 7196 18264
rect 7248 18255 7250 18264
rect 7196 18226 7248 18232
rect 7104 18216 7156 18222
rect 7208 18195 7236 18226
rect 7104 18158 7156 18164
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7116 17649 7144 17818
rect 7196 17672 7248 17678
rect 7102 17640 7158 17649
rect 7196 17614 7248 17620
rect 7102 17575 7158 17584
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17338 7144 17478
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 6932 17054 7052 17082
rect 6932 12918 6960 17054
rect 7208 16454 7236 17614
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7300 16266 7328 23072
rect 7484 20584 7512 23140
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7576 22642 7604 22986
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 8036 22098 8064 23462
rect 7668 22066 7972 22094
rect 7668 22030 7696 22066
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 7944 21978 7972 22066
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 8116 22024 8168 22030
rect 7944 21972 8116 21978
rect 7944 21966 8168 21972
rect 7852 21690 7880 21966
rect 7944 21950 8156 21966
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7576 20777 7604 20810
rect 7562 20768 7618 20777
rect 7562 20703 7618 20712
rect 7392 20556 7512 20584
rect 7392 16658 7420 20556
rect 7564 20528 7616 20534
rect 7484 20488 7564 20516
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7208 16238 7328 16266
rect 7208 16182 7236 16238
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7104 15088 7156 15094
rect 7156 15048 7236 15076
rect 7104 15030 7156 15036
rect 7208 14958 7236 15048
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7012 14272 7064 14278
rect 7208 14249 7236 14282
rect 7288 14272 7340 14278
rect 7012 14214 7064 14220
rect 7194 14240 7250 14249
rect 7024 13870 7052 14214
rect 7288 14214 7340 14220
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7194 14175 7250 14184
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7010 11928 7066 11937
rect 7010 11863 7012 11872
rect 7064 11863 7066 11872
rect 7012 11834 7064 11840
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 7024 10674 7052 11698
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9500 6776 9862
rect 6932 9654 6960 10066
rect 7024 9722 7052 10610
rect 7116 10169 7144 11086
rect 7102 10160 7158 10169
rect 7102 10095 7158 10104
rect 7012 9716 7064 9722
rect 7064 9664 7144 9674
rect 7012 9658 7144 9664
rect 6920 9648 6972 9654
rect 7024 9646 7144 9658
rect 6920 9590 6972 9596
rect 6828 9512 6880 9518
rect 6748 9472 6828 9500
rect 6828 9454 6880 9460
rect 6828 9036 6880 9042
rect 6932 9024 6960 9590
rect 7116 9178 7144 9646
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6880 8996 6960 9024
rect 6828 8978 6880 8984
rect 6826 8936 6882 8945
rect 6826 8871 6882 8880
rect 6840 8838 6868 8871
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6932 8430 6960 8996
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8498 7052 8774
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6932 7954 6960 8366
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7410 6960 7890
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 6748 3194 6776 6734
rect 6840 3738 6868 6802
rect 7116 5370 7144 8298
rect 7208 6662 7236 12174
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5710 7236 6258
rect 7300 5914 7328 14214
rect 7392 14074 7420 14214
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7392 10606 7420 12718
rect 7484 12442 7512 20488
rect 7564 20470 7616 20476
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7576 19310 7604 20334
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7576 18902 7604 19246
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7668 16674 7696 18022
rect 7760 17610 7788 21626
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7852 19786 7880 21286
rect 8128 21010 8156 21490
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8220 20210 8248 35022
rect 8864 30258 8892 36654
rect 10244 31346 10272 36858
rect 11624 36378 11652 37198
rect 12268 37108 12296 39200
rect 13556 37262 13584 39200
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 14648 37188 14700 37194
rect 14648 37130 14700 37136
rect 12440 37120 12492 37126
rect 12268 37080 12440 37108
rect 12440 37062 12492 37068
rect 14280 37120 14332 37126
rect 14280 37062 14332 37068
rect 13820 36848 13872 36854
rect 13820 36790 13872 36796
rect 11612 36372 11664 36378
rect 11612 36314 11664 36320
rect 11796 36168 11848 36174
rect 11796 36110 11848 36116
rect 11808 32026 11836 36110
rect 11888 33856 11940 33862
rect 11888 33798 11940 33804
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 11520 31136 11572 31142
rect 11520 31078 11572 31084
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8864 24818 8892 26726
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10612 25362 10640 25638
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 11532 25294 11560 31078
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11808 25906 11836 26318
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11808 25362 11836 25638
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 9876 24818 9904 25230
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 9864 24812 9916 24818
rect 9864 24754 9916 24760
rect 11244 24812 11296 24818
rect 11244 24754 11296 24760
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9416 23322 9444 23666
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9312 23248 9364 23254
rect 9312 23190 9364 23196
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8496 22098 8524 22578
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8220 20182 8340 20210
rect 8312 19990 8340 20182
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8022 19816 8078 19825
rect 7840 19780 7892 19786
rect 8022 19751 8024 19760
rect 7840 19722 7892 19728
rect 8076 19751 8078 19760
rect 8024 19722 8076 19728
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7840 18352 7892 18358
rect 7838 18320 7840 18329
rect 7892 18320 7894 18329
rect 7838 18255 7894 18264
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7668 16646 7788 16674
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7668 16250 7696 16458
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7760 15434 7788 16646
rect 7944 15638 7972 19178
rect 8312 18902 8340 19926
rect 8404 19922 8432 21966
rect 8496 21078 8524 22034
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 8484 20936 8536 20942
rect 8484 20878 8536 20884
rect 8496 19961 8524 20878
rect 8588 20398 8616 22646
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8772 21486 8800 21558
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8576 20392 8628 20398
rect 9128 20392 9180 20398
rect 8576 20334 8628 20340
rect 9126 20360 9128 20369
rect 9180 20360 9182 20369
rect 8482 19952 8538 19961
rect 8392 19916 8444 19922
rect 8482 19887 8538 19896
rect 8392 19858 8444 19864
rect 8588 19334 8616 20334
rect 9126 20295 9182 20304
rect 8666 19544 8722 19553
rect 8666 19479 8722 19488
rect 8496 19306 8616 19334
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8312 18601 8340 18702
rect 8298 18592 8354 18601
rect 8298 18527 8354 18536
rect 8208 18148 8260 18154
rect 8208 18090 8260 18096
rect 8220 17814 8248 18090
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8036 16658 8064 17546
rect 8116 16992 8168 16998
rect 8114 16960 8116 16969
rect 8168 16960 8170 16969
rect 8114 16895 8170 16904
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 8036 15434 8064 16390
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7852 13841 7880 15030
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14550 8156 14758
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8022 14376 8078 14385
rect 8022 14311 8078 14320
rect 7838 13832 7894 13841
rect 7838 13767 7894 13776
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10674 7512 10950
rect 7576 10810 7604 12718
rect 7760 12186 7788 13194
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7852 12306 7880 12854
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7760 12158 7880 12186
rect 7654 11656 7710 11665
rect 7654 11591 7710 11600
rect 7668 11218 7696 11591
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7208 4622 7236 5646
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 7024 2446 7052 2790
rect 7300 2514 7328 4966
rect 7392 2650 7420 9998
rect 7484 5778 7512 10134
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 9042 7604 9454
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7760 7478 7788 11222
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7576 4826 7604 7278
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7760 5234 7788 5510
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7852 4486 7880 12158
rect 7944 11830 7972 12582
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 8036 10266 8064 14311
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8128 12782 8156 13942
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8128 12646 8156 12718
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8116 12368 8168 12374
rect 8114 12336 8116 12345
rect 8168 12336 8170 12345
rect 8114 12271 8170 12280
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 10266 8156 12174
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7944 8430 7972 9386
rect 8128 9178 8156 9658
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8036 8430 8064 8502
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7930 8120 7986 8129
rect 7930 8055 7932 8064
rect 7984 8055 7986 8064
rect 7932 8026 7984 8032
rect 7930 6896 7986 6905
rect 7930 6831 7986 6840
rect 7944 6458 7972 6831
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7944 6118 7972 6258
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 8128 4010 8156 8230
rect 8220 5234 8248 17750
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8312 11286 8340 17206
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16726 8432 16934
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8404 16289 8432 16390
rect 8390 16280 8446 16289
rect 8390 16215 8446 16224
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8404 14482 8432 15506
rect 8496 15178 8524 19306
rect 8574 18728 8630 18737
rect 8574 18663 8576 18672
rect 8628 18663 8630 18672
rect 8576 18634 8628 18640
rect 8680 17814 8708 19479
rect 9034 19272 9090 19281
rect 9034 19207 9036 19216
rect 9088 19207 9090 19216
rect 9036 19178 9088 19184
rect 9128 19168 9180 19174
rect 9126 19136 9128 19145
rect 9180 19136 9182 19145
rect 9126 19071 9182 19080
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8680 17202 8708 17750
rect 8864 17270 8892 18566
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8588 15337 8616 16050
rect 8956 15638 8984 18770
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9140 18290 9168 18362
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9126 17912 9182 17921
rect 9126 17847 9182 17856
rect 9140 17746 9168 17847
rect 9232 17746 9260 22442
rect 9324 22094 9352 23190
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9416 22778 9444 23054
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9600 22642 9628 23530
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23186 9720 23462
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9324 22066 9444 22094
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 9324 19854 9352 21014
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9312 19440 9364 19446
rect 9310 19408 9312 19417
rect 9364 19408 9366 19417
rect 9310 19343 9366 19352
rect 9416 18426 9444 22066
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9692 17882 9720 22918
rect 9770 21992 9826 22001
rect 9770 21927 9826 21936
rect 9784 21486 9812 21927
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9772 21344 9824 21350
rect 9876 21321 9904 24754
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 22710 10640 22918
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10244 22234 10272 22510
rect 10232 22228 10284 22234
rect 10232 22170 10284 22176
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9968 21350 9996 21966
rect 10508 21956 10560 21962
rect 10508 21898 10560 21904
rect 10416 21616 10468 21622
rect 10416 21558 10468 21564
rect 9956 21344 10008 21350
rect 9772 21286 9824 21292
rect 9862 21312 9918 21321
rect 9784 20534 9812 21286
rect 10008 21304 10272 21332
rect 9956 21286 10008 21292
rect 9862 21247 9918 21256
rect 10046 21176 10102 21185
rect 9864 21140 9916 21146
rect 9916 21120 10046 21128
rect 9916 21111 10102 21120
rect 9916 21100 10088 21111
rect 9864 21082 9916 21088
rect 9862 21040 9918 21049
rect 10244 21010 10272 21304
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 9862 20975 9918 20984
rect 9956 21004 10008 21010
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9784 19990 9812 20470
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9784 19446 9812 19926
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9784 18834 9812 19382
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9402 17776 9458 17785
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9220 17740 9272 17746
rect 9402 17711 9404 17720
rect 9220 17682 9272 17688
rect 9456 17711 9458 17720
rect 9404 17682 9456 17688
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9140 16590 9168 17138
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16114 9168 16526
rect 9416 16522 9444 17478
rect 9784 17354 9812 18226
rect 9692 17326 9812 17354
rect 9496 16992 9548 16998
rect 9494 16960 9496 16969
rect 9548 16960 9550 16969
rect 9494 16895 9550 16904
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8944 15632 8996 15638
rect 8944 15574 8996 15580
rect 8574 15328 8630 15337
rect 8574 15263 8630 15272
rect 8496 15150 8616 15178
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8496 13682 8524 13806
rect 8404 13654 8524 13682
rect 8404 13258 8432 13654
rect 8588 13546 8616 15150
rect 9140 15094 9168 16050
rect 9508 15994 9536 16458
rect 9324 15966 9536 15994
rect 9128 15088 9180 15094
rect 9048 15048 9128 15076
rect 9048 14482 9076 15048
rect 9128 15030 9180 15036
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9140 14618 9168 14894
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9324 14521 9352 15966
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9310 14512 9366 14521
rect 9036 14476 9088 14482
rect 9310 14447 9366 14456
rect 9036 14418 9088 14424
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8496 13518 8616 13546
rect 8496 13394 8524 13518
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8390 13016 8446 13025
rect 8390 12951 8392 12960
rect 8444 12951 8446 12960
rect 8392 12922 8444 12928
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8588 12434 8616 12582
rect 8496 12406 8616 12434
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10062 8340 11086
rect 8404 10538 8432 12242
rect 8496 11082 8524 12406
rect 8680 12170 8708 14214
rect 9048 14090 9076 14418
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 8772 14062 9076 14090
rect 8772 14006 8800 14062
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13705 8984 13942
rect 8942 13696 8998 13705
rect 8942 13631 8998 13640
rect 9048 13394 9076 14062
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8574 11792 8630 11801
rect 8574 11727 8630 11736
rect 8588 11082 8616 11727
rect 8680 11694 8708 12106
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8312 9110 8340 9658
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8312 8945 8340 9046
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 6118 8340 7686
rect 8404 6458 8432 9590
rect 8496 8838 8524 11018
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8588 10198 8616 10678
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9450 8616 9998
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8496 8294 8524 8502
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8496 3398 8524 7414
rect 8680 6390 8708 11222
rect 8864 10470 8892 13194
rect 9324 13138 9352 14282
rect 9416 13258 9444 15846
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9600 15366 9628 15438
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9508 14278 9536 15098
rect 9692 14464 9720 17326
rect 9772 17264 9824 17270
rect 9876 17252 9904 20975
rect 9956 20946 10008 20952
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 9968 20913 9996 20946
rect 10048 20936 10100 20942
rect 9954 20904 10010 20913
rect 10336 20890 10364 21082
rect 10100 20884 10364 20890
rect 10048 20878 10364 20884
rect 10060 20862 10364 20878
rect 9954 20839 10010 20848
rect 9954 20496 10010 20505
rect 9954 20431 10010 20440
rect 9824 17224 9904 17252
rect 9772 17206 9824 17212
rect 9784 15162 9812 17206
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9692 14436 9812 14464
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13852 9536 14214
rect 9692 13977 9720 14282
rect 9784 14006 9812 14436
rect 9968 14226 9996 20431
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10060 18970 10088 20334
rect 10152 19854 10180 20862
rect 10428 20505 10456 21558
rect 10520 21486 10548 21898
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10520 21010 10548 21286
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10520 20913 10548 20946
rect 10506 20904 10562 20913
rect 10612 20874 10640 20946
rect 10506 20839 10562 20848
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10414 20496 10470 20505
rect 10414 20431 10470 20440
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10796 19961 10824 20402
rect 10782 19952 10838 19961
rect 10782 19887 10838 19896
rect 10140 19848 10192 19854
rect 10192 19808 10272 19836
rect 10140 19790 10192 19796
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10046 18456 10102 18465
rect 10046 18391 10102 18400
rect 10060 18222 10088 18391
rect 10152 18358 10180 18702
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10152 16266 10180 18294
rect 10244 17134 10272 19808
rect 10600 19780 10652 19786
rect 10888 19768 10916 23802
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 10980 22098 11008 23666
rect 11256 23118 11284 24754
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11808 24206 11836 24550
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11520 24132 11572 24138
rect 11520 24074 11572 24080
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10980 21554 11008 22034
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 19786 11008 21490
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11072 20777 11100 20810
rect 11058 20768 11114 20777
rect 11058 20703 11114 20712
rect 11164 20602 11192 22170
rect 11256 22094 11284 23054
rect 11256 22066 11468 22094
rect 11336 21956 11388 21962
rect 11336 21898 11388 21904
rect 11348 20777 11376 21898
rect 11334 20768 11390 20777
rect 11334 20703 11390 20712
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 10652 19740 10916 19768
rect 10600 19722 10652 19728
rect 10506 19408 10562 19417
rect 10506 19343 10562 19352
rect 10782 19408 10838 19417
rect 10888 19394 10916 19740
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10888 19366 11008 19394
rect 10782 19343 10784 19352
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 17728 10364 18634
rect 10520 18290 10548 19343
rect 10836 19343 10838 19352
rect 10784 19314 10836 19320
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10980 19258 11008 19366
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10336 17700 10456 17728
rect 10322 17640 10378 17649
rect 10322 17575 10378 17584
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10060 16238 10180 16266
rect 10060 16046 10088 16238
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10152 15337 10180 16118
rect 10138 15328 10194 15337
rect 10138 15263 10194 15272
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9876 14198 9996 14226
rect 9772 14000 9824 14006
rect 9678 13968 9734 13977
rect 9772 13942 9824 13948
rect 9678 13903 9734 13912
rect 9680 13864 9732 13870
rect 9508 13824 9680 13852
rect 9680 13806 9732 13812
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9324 13110 9444 13138
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9048 12374 9076 12718
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9126 12064 9182 12073
rect 9126 11999 9182 12008
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8772 9654 8800 10406
rect 8956 9722 8984 10610
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8760 9512 8812 9518
rect 9048 9466 9076 11766
rect 9140 10690 9168 11999
rect 9324 11898 9352 12718
rect 9416 12434 9444 13110
rect 9494 12880 9550 12889
rect 9494 12815 9496 12824
rect 9548 12815 9550 12824
rect 9496 12786 9548 12792
rect 9416 12406 9628 12434
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9508 11898 9536 12174
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9404 11824 9456 11830
rect 9404 11766 9456 11772
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11218 9260 11562
rect 9416 11354 9444 11766
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9496 11280 9548 11286
rect 9416 11228 9496 11234
rect 9416 11222 9548 11228
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9416 11206 9536 11222
rect 9140 10662 9352 10690
rect 9128 10192 9180 10198
rect 9126 10160 9128 10169
rect 9180 10160 9182 10169
rect 9126 10095 9182 10104
rect 8760 9454 8812 9460
rect 8772 9382 8800 9454
rect 8864 9438 9076 9466
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8864 5030 8892 9438
rect 9036 9376 9088 9382
rect 8942 9344 8998 9353
rect 9036 9318 9088 9324
rect 8942 9279 8998 9288
rect 8956 9042 8984 9279
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 9048 8974 9076 9318
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9324 8634 9352 10662
rect 9416 9586 9444 11206
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9508 9178 9536 11086
rect 9600 10130 9628 12406
rect 9692 10169 9720 13670
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12646 9812 13126
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 10742 9812 12582
rect 9876 11257 9904 14198
rect 10060 14074 10088 14554
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10244 13841 10272 14962
rect 10230 13832 10286 13841
rect 10230 13767 10286 13776
rect 10336 13734 10364 17575
rect 10428 17134 10456 17700
rect 10520 17678 10548 18022
rect 10612 17814 10640 18634
rect 10888 18358 10916 19246
rect 10980 19230 11100 19258
rect 11072 19174 11100 19230
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10876 18352 10928 18358
rect 10782 18320 10838 18329
rect 10876 18294 10928 18300
rect 11164 18290 11192 20538
rect 11348 20369 11376 20538
rect 11334 20360 11390 20369
rect 11334 20295 11390 20304
rect 11440 19938 11468 22066
rect 11348 19910 11468 19938
rect 11348 18329 11376 19910
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11334 18320 11390 18329
rect 10782 18255 10838 18264
rect 11152 18284 11204 18290
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10520 14550 10548 17614
rect 10612 16658 10640 17750
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10704 16697 10732 17206
rect 10690 16688 10746 16697
rect 10600 16652 10652 16658
rect 10690 16623 10746 16632
rect 10600 16594 10652 16600
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10612 14385 10640 14486
rect 10598 14376 10654 14385
rect 10598 14311 10654 14320
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10322 13560 10378 13569
rect 10322 13495 10378 13504
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9862 11248 9918 11257
rect 9862 11183 9918 11192
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9678 10160 9734 10169
rect 9588 10124 9640 10130
rect 9678 10095 9734 10104
rect 9588 10066 9640 10072
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9600 9897 9628 9930
rect 9586 9888 9642 9897
rect 9586 9823 9642 9832
rect 9496 9172 9548 9178
rect 9772 9172 9824 9178
rect 9496 9114 9548 9120
rect 9692 9132 9772 9160
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9324 8362 9352 8570
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9692 7886 9720 9132
rect 9772 9114 9824 9120
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8956 7002 8984 7142
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9048 6662 9076 6870
rect 9128 6792 9180 6798
rect 9404 6792 9456 6798
rect 9180 6752 9404 6780
rect 9128 6734 9180 6740
rect 9404 6734 9456 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9140 6202 9168 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8956 6186 9168 6202
rect 8944 6180 9168 6186
rect 8996 6174 9168 6180
rect 8944 6122 8996 6128
rect 9232 5914 9260 6326
rect 9692 6254 9720 7822
rect 9876 6866 9904 11086
rect 9968 10826 9996 13194
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10046 13016 10102 13025
rect 10046 12951 10102 12960
rect 10060 12850 10088 12951
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10046 12200 10102 12209
rect 10046 12135 10048 12144
rect 10100 12135 10102 12144
rect 10048 12106 10100 12112
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10060 11558 10088 11630
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9968 10798 10088 10826
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9968 10266 9996 10678
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10060 8022 10088 10798
rect 10152 9586 10180 13126
rect 10336 12986 10364 13495
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10704 12442 10732 14894
rect 10796 14482 10824 18255
rect 11204 18244 11284 18272
rect 11334 18255 11390 18264
rect 11152 18226 11204 18232
rect 11256 17746 11284 18244
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11348 17678 11376 18022
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11072 16794 11100 17274
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16114 11192 16390
rect 11440 16153 11468 19722
rect 11532 16250 11560 24074
rect 11900 23186 11928 33798
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 11980 26240 12032 26246
rect 11980 26182 12032 26188
rect 11992 25906 12020 26182
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12360 24138 12388 24754
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23186 12112 24006
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12268 22710 12296 23462
rect 12452 23322 12480 29990
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12544 25974 12572 26318
rect 12532 25968 12584 25974
rect 12532 25910 12584 25916
rect 12440 23316 12492 23322
rect 12440 23258 12492 23264
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12360 22166 12388 22918
rect 12348 22160 12400 22166
rect 12348 22102 12400 22108
rect 12452 21894 12480 23258
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 11794 21040 11850 21049
rect 11794 20975 11850 20984
rect 11808 20806 11836 20975
rect 12254 20904 12310 20913
rect 12254 20839 12310 20848
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11624 18057 11652 18634
rect 11610 18048 11666 18057
rect 11610 17983 11666 17992
rect 11716 16998 11744 20538
rect 12268 20330 12296 20839
rect 12452 20482 12480 21558
rect 12544 20602 12572 25910
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12636 25498 12664 25842
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12636 23730 12664 24210
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12636 21978 12664 23666
rect 12820 22574 12848 24006
rect 12912 22710 12940 31758
rect 13832 31346 13860 36790
rect 14292 33998 14320 37062
rect 14660 34746 14688 37130
rect 15488 37126 15516 39200
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 14832 35080 14884 35086
rect 14832 35022 14884 35028
rect 14648 34740 14700 34746
rect 14648 34682 14700 34688
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14556 34128 14608 34134
rect 14556 34070 14608 34076
rect 14280 33992 14332 33998
rect 14280 33934 14332 33940
rect 13820 31340 13872 31346
rect 13820 31282 13872 31288
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13360 25424 13412 25430
rect 13360 25366 13412 25372
rect 13372 25158 13400 25366
rect 13556 25362 13584 25774
rect 14004 25696 14056 25702
rect 14004 25638 14056 25644
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13372 24818 13400 25094
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12898 22128 12954 22137
rect 12898 22063 12954 22072
rect 12912 22030 12940 22063
rect 12900 22024 12952 22030
rect 12636 21950 12756 21978
rect 12900 21966 12952 21972
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12636 21185 12664 21490
rect 12622 21176 12678 21185
rect 12622 21111 12678 21120
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12636 20534 12664 21111
rect 12624 20528 12676 20534
rect 12452 20454 12572 20482
rect 12624 20470 12676 20476
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11808 17882 11836 19314
rect 11900 18358 11928 19450
rect 11992 19310 12020 19994
rect 12452 19786 12480 20266
rect 12440 19780 12492 19786
rect 12440 19722 12492 19728
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 19378 12296 19654
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12162 19272 12218 19281
rect 12162 19207 12218 19216
rect 12176 19174 12204 19207
rect 12072 19168 12124 19174
rect 11978 19136 12034 19145
rect 12072 19110 12124 19116
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 11978 19071 12034 19080
rect 11992 18873 12020 19071
rect 12084 18902 12112 19110
rect 12072 18896 12124 18902
rect 11978 18864 12034 18873
rect 12072 18838 12124 18844
rect 11978 18799 12034 18808
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 12176 18154 12204 18362
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11426 16144 11482 16153
rect 11152 16108 11204 16114
rect 11426 16079 11482 16088
rect 11152 16050 11204 16056
rect 11532 16046 11560 16186
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10888 15638 10916 15846
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 14249 10824 14418
rect 10782 14240 10838 14249
rect 10782 14175 10838 14184
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10796 12646 10824 13194
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10336 11626 10364 11834
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10152 8294 10180 9046
rect 10244 8634 10272 11562
rect 10428 10810 10456 11630
rect 10520 11286 10548 12242
rect 10612 11937 10640 12310
rect 10598 11928 10654 11937
rect 10598 11863 10654 11872
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10508 11280 10560 11286
rect 10508 11222 10560 11228
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10336 7886 10364 8910
rect 10520 8498 10548 10950
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10520 7970 10548 8434
rect 10612 8090 10640 11086
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10520 7954 10640 7970
rect 10520 7948 10652 7954
rect 10520 7942 10600 7948
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9968 7478 9996 7686
rect 10336 7546 10364 7822
rect 10520 7818 10548 7942
rect 10600 7890 10652 7896
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 10060 6866 10088 7482
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6458 10088 6802
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 10704 5914 10732 11698
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10796 9926 10824 10202
rect 10888 10062 10916 10406
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10888 9586 10916 9998
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 8498 10824 9454
rect 10980 9042 11008 15982
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11164 14074 11192 15642
rect 11716 15337 11744 15982
rect 11808 15434 11836 16934
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11702 15328 11758 15337
rect 11702 15263 11758 15272
rect 11242 15192 11298 15201
rect 11242 15127 11298 15136
rect 11256 14822 11284 15127
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 9654 11100 13806
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11164 12782 11192 13670
rect 11256 13530 11284 13670
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11348 12986 11376 14758
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11440 12374 11468 13806
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10876 8900 10928 8906
rect 11072 8888 11100 8978
rect 10928 8860 11100 8888
rect 10876 8842 10928 8848
rect 11164 8634 11192 12106
rect 11440 11898 11468 12310
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 9140 2446 9168 4966
rect 10060 3058 10088 5578
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10796 2446 10824 7142
rect 10888 4758 10916 7754
rect 10980 7342 11008 8434
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11164 7154 11192 7414
rect 10980 7126 11192 7154
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10980 4690 11008 7126
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11072 4078 11100 6666
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11164 2650 11192 5646
rect 11256 5098 11284 8842
rect 11348 5846 11376 11630
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11440 6458 11468 9930
rect 11532 8634 11560 14282
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11624 12646 11652 13398
rect 11808 13326 11836 15370
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11150 11652 12038
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11716 10606 11744 13262
rect 11900 11354 11928 15982
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11992 10266 12020 15438
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12084 13841 12112 14282
rect 12070 13832 12126 13841
rect 12070 13767 12126 13776
rect 12070 13696 12126 13705
rect 12070 13631 12126 13640
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11716 8362 11744 8434
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11716 8022 11744 8298
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11808 7546 11836 7890
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11900 6866 11928 9454
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11992 6662 12020 10095
rect 12084 9450 12112 13631
rect 12176 12646 12204 16526
rect 12268 16182 12296 19314
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12360 19145 12388 19178
rect 12346 19136 12402 19145
rect 12346 19071 12402 19080
rect 12346 18184 12402 18193
rect 12346 18119 12348 18128
rect 12400 18119 12402 18128
rect 12348 18090 12400 18096
rect 12544 17678 12572 20454
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12636 19009 12664 19382
rect 12728 19378 12756 21950
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12728 19145 12756 19314
rect 12714 19136 12770 19145
rect 12714 19071 12770 19080
rect 12622 19000 12678 19009
rect 12622 18935 12678 18944
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12636 17746 12664 18022
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12544 17354 12572 17614
rect 12360 17326 12572 17354
rect 12360 16266 12388 17326
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 16454 12664 17206
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12360 16238 12480 16266
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12268 11354 12296 15438
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12360 13705 12388 15030
rect 12346 13696 12402 13705
rect 12346 13631 12402 13640
rect 12360 13326 12388 13357
rect 12348 13320 12400 13326
rect 12452 13274 12480 16238
rect 12728 15450 12756 16390
rect 12820 15570 12848 21830
rect 13004 21622 13032 24006
rect 13096 23866 13124 24142
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 13096 23186 13124 23598
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 13188 23050 13216 24550
rect 13740 24410 13768 24686
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 14016 24274 14044 25638
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 14108 23186 14136 29106
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 14280 25696 14332 25702
rect 14280 25638 14332 25644
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12912 20874 12940 21354
rect 13464 21010 13492 22646
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 13924 21962 13952 22374
rect 13912 21956 13964 21962
rect 13912 21898 13964 21904
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13096 18222 13124 19790
rect 13280 19394 13308 20946
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13280 19366 13492 19394
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18766 13400 19246
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 18272 13400 18566
rect 13188 18244 13400 18272
rect 13084 18216 13136 18222
rect 13188 18204 13216 18244
rect 13136 18176 13216 18204
rect 13084 18158 13136 18164
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17746 13124 18022
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13096 17542 13124 17682
rect 13464 17542 13492 19366
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13464 17066 13492 17274
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12636 15422 12756 15450
rect 12808 15428 12860 15434
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12400 13268 12480 13274
rect 12348 13262 12480 13268
rect 12360 13246 12480 13262
rect 12360 12764 12388 13246
rect 12360 12736 12480 12764
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12176 6662 12204 11222
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12268 10742 12296 11154
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12268 9654 12296 10678
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12360 8634 12388 12174
rect 12452 11830 12480 12736
rect 12544 12374 12572 14894
rect 12636 14618 12664 15422
rect 12808 15370 12860 15376
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 14482 12756 15302
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12820 14362 12848 15370
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12636 14334 12848 14362
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12636 13734 12664 14334
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12617 12664 13262
rect 12622 12608 12678 12617
rect 12622 12543 12678 12552
rect 12532 12368 12584 12374
rect 12716 12368 12768 12374
rect 12532 12310 12584 12316
rect 12622 12336 12678 12345
rect 12716 12310 12768 12316
rect 12622 12271 12678 12280
rect 12532 12232 12584 12238
rect 12530 12200 12532 12209
rect 12584 12200 12586 12209
rect 12530 12135 12586 12144
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12544 11762 12572 12135
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12544 9994 12572 10542
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12452 6882 12480 9522
rect 12636 9178 12664 12271
rect 12728 10266 12756 12310
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8498 12572 8774
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12452 6866 12572 6882
rect 12452 6860 12584 6866
rect 12452 6854 12532 6860
rect 12532 6802 12584 6808
rect 12728 6746 12756 10066
rect 12820 9654 12848 13806
rect 12912 12434 12940 14350
rect 13004 14006 13032 14758
rect 13280 14550 13308 14894
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13176 14408 13228 14414
rect 13372 14396 13400 16118
rect 13556 15502 13584 20402
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13636 19304 13688 19310
rect 13740 19292 13768 20266
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13832 19514 13860 19654
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13820 19304 13872 19310
rect 13740 19264 13820 19292
rect 13636 19246 13688 19252
rect 13820 19246 13872 19252
rect 13648 17338 13676 19246
rect 13924 18970 13952 21898
rect 14016 21894 14044 22374
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13740 16658 13768 18158
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13832 16250 13860 16594
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13556 15026 13584 15438
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13176 14350 13228 14356
rect 13280 14368 13400 14396
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 14074 13124 14282
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12646 13124 13126
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12912 12406 13124 12434
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12912 11801 12940 12106
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12898 11792 12954 11801
rect 12898 11727 12954 11736
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12360 6730 12756 6746
rect 12348 6724 12756 6730
rect 12400 6718 12756 6724
rect 12348 6666 12400 6672
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 12820 4826 12848 8910
rect 12912 8090 12940 11630
rect 13004 11286 13032 12038
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 13096 10690 13124 12406
rect 13188 10810 13216 14350
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13004 8634 13032 10678
rect 13096 10662 13216 10690
rect 13280 10674 13308 14368
rect 13648 13530 13676 15846
rect 13832 15162 13860 16050
rect 13924 15706 13952 18226
rect 14016 16046 14044 21830
rect 14108 21622 14136 23122
rect 14200 22094 14228 25230
rect 14292 24818 14320 25638
rect 14476 25362 14504 26454
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14476 23186 14504 24006
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14280 23112 14332 23118
rect 14278 23080 14280 23089
rect 14332 23080 14334 23089
rect 14278 23015 14334 23024
rect 14292 22234 14320 23015
rect 14568 22642 14596 34070
rect 14752 29730 14780 34546
rect 14844 29850 14872 35022
rect 15580 34746 15608 37198
rect 15844 37188 15896 37194
rect 15844 37130 15896 37136
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14752 29702 14872 29730
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14752 25498 14780 29582
rect 14844 28762 14872 29702
rect 15028 29306 15056 34546
rect 15856 33998 15884 37130
rect 16776 37126 16804 39200
rect 18064 37262 18092 39200
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16868 35290 16896 37198
rect 16856 35284 16908 35290
rect 16856 35226 16908 35232
rect 18524 34746 18552 37198
rect 19996 37126 20024 39200
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 20640 34746 20668 37198
rect 20904 37188 20956 37194
rect 20904 37130 20956 37136
rect 18512 34740 18564 34746
rect 18512 34682 18564 34688
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17500 34536 17552 34542
rect 17500 34478 17552 34484
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 15108 33856 15160 33862
rect 15108 33798 15160 33804
rect 15016 29300 15068 29306
rect 15016 29242 15068 29248
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 15120 26874 15148 33798
rect 16304 31884 16356 31890
rect 16304 31826 16356 31832
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 15844 29640 15896 29646
rect 15844 29582 15896 29588
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 14936 26846 15148 26874
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14752 24954 14780 25434
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14200 22066 14320 22094
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 14200 19446 14228 21422
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 14200 17134 14228 19382
rect 14292 18698 14320 22066
rect 14556 22024 14608 22030
rect 14608 21972 14688 21978
rect 14556 21966 14688 21972
rect 14568 21950 14688 21966
rect 14844 21962 14872 23462
rect 14660 21690 14688 21950
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14740 21480 14792 21486
rect 14740 21422 14792 21428
rect 14556 21344 14608 21350
rect 14556 21286 14608 21292
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 18970 14412 20334
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19310 14504 20198
rect 14568 19854 14596 21286
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14660 20534 14688 20878
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14752 20058 14780 21422
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14844 21078 14872 21286
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14292 17678 14320 18634
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14292 16590 14320 17138
rect 14844 17134 14872 21014
rect 14936 21010 14964 26846
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15304 25906 15332 26318
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15200 25696 15252 25702
rect 15200 25638 15252 25644
rect 15212 24886 15240 25638
rect 15200 24880 15252 24886
rect 15200 24822 15252 24828
rect 15016 23248 15068 23254
rect 15016 23190 15068 23196
rect 15028 22574 15056 23190
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15120 22710 15148 22918
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 15016 22568 15068 22574
rect 15016 22510 15068 22516
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 15028 19718 15056 21558
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15108 21072 15160 21078
rect 15106 21040 15108 21049
rect 15160 21040 15162 21049
rect 15106 20975 15162 20984
rect 15212 19990 15240 21286
rect 15304 20913 15332 25842
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15396 22778 15424 23054
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15672 22710 15700 29106
rect 15856 23798 15884 29582
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 15948 25362 15976 25774
rect 15936 25356 15988 25362
rect 15936 25298 15988 25304
rect 16224 24274 16252 31078
rect 16212 24268 16264 24274
rect 16212 24210 16264 24216
rect 15844 23792 15896 23798
rect 15844 23734 15896 23740
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15672 22094 15700 22646
rect 15856 22094 15884 23734
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 16028 22976 16080 22982
rect 16028 22918 16080 22924
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15580 22066 15700 22094
rect 15764 22066 15884 22094
rect 15290 20904 15346 20913
rect 15290 20839 15346 20848
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 15304 20534 15332 20742
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15580 20398 15608 22066
rect 15764 22030 15792 22066
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15856 21554 15884 21830
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15764 20806 15792 21422
rect 15948 20942 15976 22578
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15396 19922 15424 20198
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15120 19530 15148 19654
rect 15028 19502 15148 19530
rect 15028 19258 15056 19502
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14936 19242 15056 19258
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14924 19236 15056 19242
rect 14976 19230 15056 19236
rect 14924 19178 14976 19184
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14936 17066 14964 17682
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 15028 16538 15056 18702
rect 15120 17678 15148 19246
rect 15212 18816 15240 19314
rect 15488 19242 15516 20334
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15488 18970 15516 19178
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15292 18828 15344 18834
rect 15212 18788 15292 18816
rect 15292 18770 15344 18776
rect 15580 18465 15608 19926
rect 15764 19854 15792 20742
rect 16040 20330 16068 22918
rect 16132 22642 16160 22986
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16224 19922 16252 22374
rect 16316 20942 16344 31826
rect 17512 29306 17540 34478
rect 17880 29850 17908 34546
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 17868 29844 17920 29850
rect 17868 29786 17920 29792
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 17224 26512 17276 26518
rect 17224 26454 17276 26460
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16868 25906 16896 26250
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24750 16620 25094
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16592 24410 16620 24686
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16960 24274 16988 25638
rect 17236 25294 17264 26454
rect 17684 26240 17736 26246
rect 17684 26182 17736 26188
rect 17696 25906 17724 26182
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17512 25362 17540 25638
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 17052 24886 17080 25094
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17868 24132 17920 24138
rect 17868 24074 17920 24080
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17696 23186 17724 23462
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16500 22030 16528 22578
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16868 22098 16896 22374
rect 17880 22137 17908 24074
rect 17972 22642 18000 24142
rect 18236 22772 18288 22778
rect 18236 22714 18288 22720
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17866 22128 17922 22137
rect 16856 22092 16908 22098
rect 17866 22063 17922 22072
rect 16856 22034 16908 22040
rect 16488 22024 16540 22030
rect 16486 21992 16488 22001
rect 16540 21992 16542 22001
rect 16486 21927 16542 21936
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 21146 16436 21286
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16684 21010 16712 21830
rect 17696 21690 17724 21898
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16316 19854 16344 20878
rect 16776 20806 16804 21082
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 17236 20058 17264 21558
rect 17684 20868 17736 20874
rect 17684 20810 17736 20816
rect 17696 20602 17724 20810
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 16316 19446 16344 19790
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15672 18630 15700 18906
rect 16316 18766 16344 19110
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 15566 18456 15622 18465
rect 15566 18391 15622 18400
rect 16316 18290 16344 18566
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15212 16794 15240 18226
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13740 14006 13768 14554
rect 13832 14482 13860 14826
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13372 12434 13400 13466
rect 13452 13456 13504 13462
rect 13728 13456 13780 13462
rect 13452 13398 13504 13404
rect 13556 13404 13728 13410
rect 13556 13398 13780 13404
rect 13464 13190 13492 13398
rect 13556 13382 13768 13398
rect 13556 13326 13584 13382
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13636 12912 13688 12918
rect 13634 12880 13636 12889
rect 13688 12880 13690 12889
rect 13634 12815 13690 12824
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13372 12406 13492 12434
rect 13082 10568 13138 10577
rect 13082 10503 13084 10512
rect 13136 10503 13138 10512
rect 13084 10474 13136 10480
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13096 5166 13124 10474
rect 13188 8974 13216 10662
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13280 8498 13308 9046
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13188 8090 13216 8434
rect 13372 8362 13400 8910
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13464 6458 13492 12406
rect 13740 12238 13768 12650
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13740 5710 13768 12174
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 9382 13860 12038
rect 13924 11354 13952 14418
rect 14004 13320 14056 13326
rect 14004 13262 14056 13268
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14016 10810 14044 13262
rect 14108 11898 14136 16118
rect 14292 15201 14320 16526
rect 14648 16516 14700 16522
rect 15028 16510 15148 16538
rect 15212 16522 15240 16730
rect 15396 16697 15424 17614
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15382 16688 15438 16697
rect 15382 16623 15438 16632
rect 14648 16458 14700 16464
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14476 16182 14504 16390
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15570 14596 15914
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14660 15450 14688 16458
rect 15120 16046 15148 16510
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 14568 15422 14688 15450
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14200 13326 14228 13942
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14186 12880 14242 12889
rect 14186 12815 14242 12824
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 14016 9178 14044 9522
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14108 8634 14136 9454
rect 14200 9110 14228 12815
rect 14476 10266 14504 13262
rect 14568 12434 14596 15422
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14660 13462 14688 13670
rect 14752 13530 14780 13874
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14844 13462 14872 15438
rect 15120 14958 15148 15982
rect 15292 15428 15344 15434
rect 15212 15388 15292 15416
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14924 13864 14976 13870
rect 15108 13864 15160 13870
rect 14976 13824 15056 13852
rect 14924 13806 14976 13812
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14568 12406 14688 12434
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9586 14504 9862
rect 14568 9654 14596 12106
rect 14660 11558 14688 12406
rect 14752 12306 14780 13330
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14660 10674 14688 11086
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14660 10198 14688 10610
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14476 7002 14504 9522
rect 14752 8634 14780 12242
rect 14936 11898 14964 13466
rect 15028 13138 15056 13824
rect 15108 13806 15160 13812
rect 15120 13394 15148 13806
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15028 13110 15148 13138
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15028 12170 15056 12650
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 14660 2650 14688 8434
rect 14844 8430 14872 8570
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14936 2650 14964 6258
rect 15028 2990 15056 12106
rect 15120 11762 15148 13110
rect 15212 12918 15240 15388
rect 15292 15370 15344 15376
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 10062 15148 11698
rect 15212 10810 15240 12718
rect 15304 11898 15332 14894
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15396 11830 15424 16458
rect 15488 16454 15516 17002
rect 15856 16522 15884 17070
rect 15844 16516 15896 16522
rect 15844 16458 15896 16464
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15638 15516 15846
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 15566 14648 15622 14657
rect 15566 14583 15568 14592
rect 15620 14583 15622 14592
rect 15568 14554 15620 14560
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 13569 15516 14350
rect 15474 13560 15530 13569
rect 15474 13495 15530 13504
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 11830 15516 13126
rect 15580 12782 15608 14418
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15672 11626 15700 13262
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10266 15608 10610
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15120 7818 15148 9998
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15672 7206 15700 11562
rect 15764 11014 15792 15370
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15856 7410 15884 16458
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15948 14278 15976 14554
rect 16040 14482 16068 17070
rect 16132 16250 16160 17138
rect 16408 16590 16436 19450
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 17202 16528 18702
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16868 18222 16896 18634
rect 17052 18426 17080 19246
rect 17130 18864 17186 18873
rect 17130 18799 17186 18808
rect 17144 18426 17172 18799
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 17132 18420 17184 18426
rect 17132 18362 17184 18368
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17052 17338 17080 18158
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17144 17814 17172 18090
rect 17132 17808 17184 17814
rect 17132 17750 17184 17756
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15948 10810 15976 12786
rect 16040 12238 16068 14282
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16132 11898 16160 13806
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16224 12646 16252 12922
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16224 10198 16252 12582
rect 16408 11354 16436 13194
rect 16500 12986 16528 15438
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16592 12442 16620 14350
rect 16684 14346 16712 16934
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17052 15706 17080 15982
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16868 15162 16896 15574
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16868 14482 16896 15098
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16684 13258 16712 13942
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16776 13138 16804 13670
rect 16684 13110 16804 13138
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16500 12170 16528 12378
rect 16684 12238 16712 13110
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16592 9382 16620 11086
rect 16776 10810 16804 12718
rect 16868 11898 16896 13126
rect 16960 12374 16988 15438
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 17052 13530 17080 13942
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 17052 8362 17080 13194
rect 17236 10062 17264 15370
rect 17328 14958 17356 19246
rect 17420 16726 17448 19790
rect 17880 19378 17908 22063
rect 17972 20398 18000 22578
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18156 20874 18184 21354
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 18064 20602 18092 20810
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 18156 20058 18184 20470
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18156 19689 18184 19790
rect 18142 19680 18198 19689
rect 18142 19615 18198 19624
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17972 18766 18000 19450
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17604 17202 17632 18702
rect 18064 18358 18092 18906
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 17684 18352 17736 18358
rect 17684 18294 17736 18300
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17696 17746 17724 18294
rect 18156 18290 18184 18566
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 18064 17542 18092 18022
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 18064 15638 18092 17478
rect 18156 17338 18184 17614
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18156 16794 18184 17274
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17408 15088 17460 15094
rect 17408 15030 17460 15036
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17420 14657 17448 15030
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17406 14648 17462 14657
rect 17512 14618 17540 14758
rect 17406 14583 17462 14592
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17420 12442 17448 14282
rect 17604 14006 17632 14418
rect 17788 14074 17816 15370
rect 17880 14890 17908 15506
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17328 11626 17356 12310
rect 17500 12232 17552 12238
rect 17604 12220 17632 13262
rect 17552 12192 17632 12220
rect 17500 12174 17552 12180
rect 17604 11762 17632 12192
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17512 10674 17540 10950
rect 17880 10742 17908 14826
rect 18156 14618 18184 16594
rect 18248 16046 18276 22714
rect 18340 21962 18368 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 20180 24274 20208 33798
rect 20916 31822 20944 37130
rect 21284 37126 21312 39200
rect 22572 37262 22600 39200
rect 24504 37262 24532 39200
rect 25792 37262 25820 39200
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 27724 37126 27752 39200
rect 27804 37256 27856 37262
rect 27804 37198 27856 37204
rect 27896 37256 27948 37262
rect 27896 37198 27948 37204
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 25044 37120 25096 37126
rect 25044 37062 25096 37068
rect 27712 37120 27764 37126
rect 27712 37062 27764 37068
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20364 24818 20392 25094
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20456 24274 20484 26250
rect 20548 24818 20576 26726
rect 20640 26382 20668 27406
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 26994 20944 27270
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20444 24268 20496 24274
rect 20444 24210 20496 24216
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 18432 23050 18460 23666
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18524 23186 18552 23462
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18420 23044 18472 23050
rect 18420 22986 18472 22992
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18340 20534 18368 21898
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18432 19718 18460 22986
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18616 22778 18644 22918
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18708 22642 18736 23462
rect 20088 23322 20116 23666
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19260 22642 19288 22918
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20180 22778 20208 23054
rect 20548 23050 20576 23190
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19076 22098 19104 22510
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19352 21672 19380 22102
rect 19444 21894 19472 22374
rect 19536 22137 19564 22374
rect 19522 22128 19578 22137
rect 19522 22063 19524 22072
rect 19576 22063 19578 22072
rect 19524 22034 19576 22040
rect 19536 22003 19564 22034
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19352 21644 19472 21672
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19352 21010 19380 21490
rect 19444 21418 19472 21644
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19996 21078 20024 21490
rect 19984 21072 20036 21078
rect 19984 21014 20036 21020
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18524 19990 18552 20878
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 20466 19472 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20466 20024 21014
rect 20076 21004 20128 21010
rect 20180 20992 20208 22578
rect 20640 22094 20668 26318
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 20824 24410 20852 24550
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 21468 24138 21496 24550
rect 21928 24342 21956 35634
rect 23032 33998 23060 37062
rect 25056 33998 25084 37062
rect 27816 36922 27844 37198
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25516 35834 25544 36722
rect 25504 35828 25556 35834
rect 25504 35770 25556 35776
rect 27908 34746 27936 37198
rect 28080 37188 28132 37194
rect 28080 37130 28132 37136
rect 27896 34740 27948 34746
rect 27896 34682 27948 34688
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 25136 33856 25188 33862
rect 25136 33798 25188 33804
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23388 25152 23440 25158
rect 23388 25094 23440 25100
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21456 24132 21508 24138
rect 21456 24074 21508 24080
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21008 23186 21036 23462
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20824 22982 20852 23054
rect 21376 22982 21404 23258
rect 20812 22976 20864 22982
rect 20812 22918 20864 22924
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 20456 22066 20668 22094
rect 20456 21554 20484 22066
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20548 21622 20576 21830
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20640 21486 20668 21898
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20456 21010 20484 21286
rect 20548 21146 20576 21286
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20128 20964 20208 20992
rect 20444 21004 20496 21010
rect 20076 20946 20128 20952
rect 20444 20946 20496 20952
rect 20088 20534 20116 20946
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20548 20346 20576 21082
rect 20456 20318 20576 20346
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 18698 18736 19654
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18892 17882 18920 19790
rect 19260 19689 19288 19858
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19340 19712 19392 19718
rect 19246 19680 19302 19689
rect 19340 19654 19392 19660
rect 19246 19615 19302 19624
rect 19352 19310 19380 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19076 18834 19104 19110
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19168 18358 19196 18566
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19260 18086 19288 19110
rect 19524 18760 19576 18766
rect 19444 18720 19524 18748
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 17338 18828 17614
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18328 16176 18380 16182
rect 18328 16118 18380 16124
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18340 15162 18368 16118
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18524 15026 18552 15914
rect 18984 15065 19012 17138
rect 19260 15094 19288 18022
rect 19444 17882 19472 18720
rect 19524 18702 19576 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19352 15570 19380 16934
rect 19628 16794 19656 17138
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16182 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19248 15088 19300 15094
rect 18970 15056 19026 15065
rect 18512 15020 18564 15026
rect 19248 15030 19300 15036
rect 18970 14991 19026 15000
rect 18512 14962 18564 14968
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 19352 14074 19380 14826
rect 19444 14482 19472 15982
rect 19996 15434 20024 19790
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 19378 20392 19654
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 20088 16046 20116 18770
rect 20272 18154 20300 19246
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 17066 20300 17614
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20260 17060 20312 17066
rect 20260 17002 20312 17008
rect 20364 16590 20392 17138
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20180 16250 20208 16526
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 15706 20300 15846
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 19984 15428 20036 15434
rect 19984 15370 20036 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18142 13560 18198 13569
rect 18142 13495 18198 13504
rect 18156 12850 18184 13495
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18156 11218 18184 11630
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17972 10674 18000 11086
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17972 10130 18000 10610
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17972 9042 18000 10066
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17316 8560 17368 8566
rect 17500 8560 17552 8566
rect 17368 8508 17500 8514
rect 17316 8502 17552 8508
rect 17328 8486 17540 8502
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 5710 17908 7142
rect 18248 6458 18276 13262
rect 18340 12986 18368 13874
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18432 11898 18460 13262
rect 18510 13016 18566 13025
rect 18510 12951 18566 12960
rect 18524 12850 18552 12951
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18510 11792 18566 11801
rect 18510 11727 18566 11736
rect 18524 11354 18552 11727
rect 18800 11558 18828 13874
rect 19340 13320 19392 13326
rect 19524 13320 19576 13326
rect 19340 13262 19392 13268
rect 19444 13280 19524 13308
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 19076 12986 19104 13194
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19352 12306 19380 13262
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19444 12186 19472 13280
rect 19524 13262 19576 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12986 20024 15030
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20088 14074 20116 14894
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20180 13870 20208 15506
rect 20272 14482 20300 15642
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20088 12306 20116 13398
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20180 12918 20208 13330
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19352 12158 19472 12186
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11694 19288 12038
rect 19352 11898 19380 12158
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11762 19472 12038
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11830 20024 12174
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18340 10266 18368 11086
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 18156 2446 18184 5510
rect 18340 2650 18368 6258
rect 18432 6254 18460 10542
rect 18524 10538 18552 11290
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19444 10810 19472 10950
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18616 10266 18644 10542
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18708 10062 18736 10406
rect 19536 10062 19564 10610
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18524 5710 18552 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 20272 9178 20300 14282
rect 20364 12374 20392 16526
rect 20456 15502 20484 20318
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 19854 20576 20198
rect 20732 19922 20760 21966
rect 20824 20942 20852 22918
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21284 22098 21312 22578
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21622 20944 21830
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 21284 21486 21312 22034
rect 21652 21622 21680 24278
rect 22020 23866 22048 24754
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 22112 22574 22140 22986
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22020 21690 22048 21966
rect 22204 21962 22232 23666
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22480 21894 22508 22986
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20640 18358 20668 18566
rect 20628 18352 20680 18358
rect 20628 18294 20680 18300
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20640 14346 20668 18090
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16114 20760 16934
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20824 15502 20852 20878
rect 20916 20806 20944 21422
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 20916 19514 20944 20742
rect 21376 20466 21404 20742
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21560 20058 21588 20878
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 21560 19446 21588 19722
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21284 18426 21312 19246
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20916 17678 20944 18226
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20916 15348 20944 17614
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17202 21496 17478
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 16658 21404 16934
rect 21560 16794 21588 19382
rect 22112 18766 22140 21490
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22296 20602 22324 20878
rect 22468 20800 22520 20806
rect 22468 20742 22520 20748
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22204 19378 22232 20198
rect 22296 19786 22324 20198
rect 22388 19990 22416 20402
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22296 18834 22324 19246
rect 22388 19174 22416 19926
rect 22480 19310 22508 20742
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22388 18290 22416 19110
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 20732 15320 20944 15348
rect 20732 14822 20760 15320
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20640 11898 20668 12174
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 11830 20760 14282
rect 20824 13870 20852 14758
rect 21192 14498 21220 16594
rect 21640 16176 21692 16182
rect 21640 16118 21692 16124
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21192 14482 21312 14498
rect 21192 14476 21324 14482
rect 21192 14470 21272 14476
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20824 12986 20852 13806
rect 20916 13530 20944 13942
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20996 13456 21048 13462
rect 20996 13398 21048 13404
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20720 11824 20772 11830
rect 20720 11766 20772 11772
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20640 11558 20668 11698
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 20824 11354 20852 12718
rect 21008 12322 21036 13398
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21100 12442 21128 13262
rect 21192 12646 21220 14470
rect 21272 14418 21324 14424
rect 21376 13462 21404 15302
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21088 12436 21140 12442
rect 21376 12434 21404 12786
rect 21088 12378 21140 12384
rect 21284 12406 21404 12434
rect 21008 12294 21128 12322
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 20916 11762 20944 12106
rect 21008 11898 21036 12106
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21100 11778 21128 12294
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 21008 11750 21128 11778
rect 21008 11694 21036 11750
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20548 10266 20576 10610
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 21192 5710 21220 8298
rect 21284 6458 21312 12406
rect 21560 12170 21588 14282
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21376 11082 21404 11222
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21468 10810 21496 11018
rect 21560 10810 21588 12106
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21652 10674 21680 16118
rect 22204 15178 22232 17070
rect 22296 15570 22324 17206
rect 22388 17202 22416 18022
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22572 17066 22600 24754
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22664 23730 22692 24686
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22756 24274 22784 24550
rect 22744 24268 22796 24274
rect 22744 24210 22796 24216
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23216 23866 23244 24006
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 23216 23186 23244 23802
rect 23400 23730 23428 25094
rect 23492 24818 23520 25842
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23584 25294 23612 25638
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23204 23180 23256 23186
rect 23204 23122 23256 23128
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22664 18222 22692 22986
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22710 23520 22918
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 23124 21894 23152 22034
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22756 20466 22784 20878
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22756 19242 22784 20402
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 22940 19514 22968 19926
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22744 19236 22796 19242
rect 22744 19178 22796 19184
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22848 17338 22876 19314
rect 22940 18834 22968 19450
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22940 18290 22968 18566
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22560 16652 22612 16658
rect 22560 16594 22612 16600
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22204 15150 22416 15178
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22112 14074 22140 14350
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22204 13870 22232 14962
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 22296 12986 22324 13874
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21744 11082 21772 11154
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 19444 2446 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 22020 2650 22048 8434
rect 22388 8362 22416 15150
rect 22572 14482 22600 16594
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22756 16250 22784 16526
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 23124 16046 23152 21830
rect 23308 20058 23336 22170
rect 23584 22114 23612 23054
rect 23492 22086 23612 22114
rect 23768 22098 23796 23462
rect 23756 22092 23808 22098
rect 23492 21690 23520 22086
rect 23756 22034 23808 22040
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23676 21486 23704 21898
rect 24228 21622 24256 26930
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24412 23186 24440 23598
rect 24400 23180 24452 23186
rect 24400 23122 24452 23128
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24412 22234 24440 22510
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24504 22114 24532 29106
rect 24412 22086 24532 22114
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24044 20330 24072 20742
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23308 19854 23336 19994
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23492 18358 23520 18634
rect 23584 18426 23612 19382
rect 23940 19236 23992 19242
rect 23940 19178 23992 19184
rect 23952 18902 23980 19178
rect 23940 18896 23992 18902
rect 23940 18838 23992 18844
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 24044 18222 24072 20266
rect 24136 18766 24164 20402
rect 24228 19922 24256 21558
rect 24412 19990 24440 22086
rect 24596 22030 24624 31078
rect 24952 30592 25004 30598
rect 24952 30534 25004 30540
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24780 23798 24808 24142
rect 24768 23792 24820 23798
rect 24768 23734 24820 23740
rect 24780 22250 24808 23734
rect 24964 22438 24992 30534
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 25056 23186 25084 23462
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 25056 22778 25084 22918
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24780 22222 24900 22250
rect 24872 22030 24900 22222
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24504 21622 24532 21966
rect 24596 21706 24624 21966
rect 25148 21894 25176 33798
rect 27264 29306 27292 34546
rect 28092 33998 28120 37130
rect 29012 37126 29040 39200
rect 30300 37244 30328 39200
rect 32232 37262 32260 39200
rect 33520 37262 33548 39200
rect 30380 37256 30432 37262
rect 30300 37216 30380 37244
rect 30380 37198 30432 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 34428 37188 34480 37194
rect 34428 37130 34480 37136
rect 29000 37120 29052 37126
rect 29000 37062 29052 37068
rect 30012 37120 30064 37126
rect 30012 37062 30064 37068
rect 30656 37120 30708 37126
rect 30656 37062 30708 37068
rect 29828 36780 29880 36786
rect 29828 36722 29880 36728
rect 29840 36378 29868 36722
rect 29828 36372 29880 36378
rect 29828 36314 29880 36320
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 28080 33992 28132 33998
rect 28080 33934 28132 33940
rect 28080 33856 28132 33862
rect 28080 33798 28132 33804
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27252 29300 27304 29306
rect 27252 29242 27304 29248
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 25240 23730 25268 24006
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25516 22778 25544 23598
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25136 21888 25188 21894
rect 25136 21830 25188 21836
rect 24596 21678 24716 21706
rect 24492 21616 24544 21622
rect 24492 21558 24544 21564
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24400 19984 24452 19990
rect 24400 19926 24452 19932
rect 24216 19916 24268 19922
rect 24216 19858 24268 19864
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 23216 16998 23244 17546
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23216 16794 23244 16934
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 22572 14090 22600 14418
rect 22480 14062 22600 14090
rect 22480 11354 22508 14062
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22572 13530 22600 13942
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22756 13326 22784 15370
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 15162 22968 15302
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22572 12220 22600 12786
rect 22652 12232 22704 12238
rect 22572 12192 22652 12220
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22480 8430 22508 11290
rect 22572 8566 22600 12192
rect 22652 12174 22704 12180
rect 22756 11014 22784 13262
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22664 2650 22692 6258
rect 22848 4622 22876 13806
rect 22940 13394 22968 15098
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 23124 12918 23152 14214
rect 23112 12912 23164 12918
rect 23112 12854 23164 12860
rect 23124 12442 23152 12854
rect 23112 12436 23164 12442
rect 23112 12378 23164 12384
rect 23216 12238 23244 15098
rect 23308 14822 23336 18158
rect 24412 17814 24440 19926
rect 24596 19394 24624 21490
rect 24688 20942 24716 21678
rect 25240 21554 25268 22578
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25424 22098 25452 22510
rect 25412 22092 25464 22098
rect 25412 22034 25464 22040
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24688 20466 24716 20878
rect 24872 20602 24900 21422
rect 25516 21146 25544 21490
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25608 21146 25636 21286
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25596 21140 25648 21146
rect 25596 21082 25648 21088
rect 25976 21078 26004 21286
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25424 20602 25452 20742
rect 25792 20602 25820 20878
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 25424 19922 25452 20538
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24688 19514 24716 19790
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25148 19514 25176 19722
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 24596 19366 24716 19394
rect 24400 17808 24452 17814
rect 24400 17750 24452 17756
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23584 17202 23612 17478
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 15026 23428 15302
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23584 12986 23612 16526
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23676 16114 23704 16390
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23952 15094 23980 17138
rect 24412 16590 24440 17614
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24044 16250 24072 16390
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24504 16046 24532 16934
rect 24596 16658 24624 17070
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24124 15496 24176 15502
rect 24688 15450 24716 19366
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25240 18290 25268 19110
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25332 17610 25360 18566
rect 25424 18358 25452 19314
rect 25412 18352 25464 18358
rect 25412 18294 25464 18300
rect 25884 17678 25912 20878
rect 25964 20800 26016 20806
rect 25964 20742 26016 20748
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 25976 20466 26004 20742
rect 26528 20466 26556 20742
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 26068 19378 26096 19654
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 26344 18766 26372 19790
rect 27540 19242 27568 32846
rect 28092 23254 28120 33798
rect 28080 23248 28132 23254
rect 28080 23190 28132 23196
rect 29748 22506 29776 36110
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 29828 30592 29880 30598
rect 29828 30534 29880 30540
rect 29840 23322 29868 30534
rect 29932 27130 29960 30670
rect 30024 30666 30052 37062
rect 30668 31346 30696 37062
rect 31760 36780 31812 36786
rect 31760 36722 31812 36728
rect 31772 33114 31800 36722
rect 31760 33108 31812 33114
rect 31760 33050 31812 33056
rect 34440 31890 34468 37130
rect 34808 37126 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34888 37256 34940 37262
rect 34888 37198 34940 37204
rect 36740 37210 36768 39200
rect 37002 38176 37058 38185
rect 37002 38111 37058 38120
rect 36912 37256 36964 37262
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 34900 36922 34928 37198
rect 36740 37182 36860 37210
rect 36912 37198 36964 37204
rect 36832 37126 36860 37182
rect 36820 37120 36872 37126
rect 36820 37062 36872 37068
rect 34888 36916 34940 36922
rect 34888 36858 34940 36864
rect 36924 36825 36952 37198
rect 36910 36816 36966 36825
rect 36176 36780 36228 36786
rect 37016 36786 37044 38111
rect 37464 37256 37516 37262
rect 37464 37198 37516 37204
rect 36910 36751 36966 36760
rect 37004 36780 37056 36786
rect 36176 36722 36228 36728
rect 37004 36722 37056 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 36188 36378 36216 36722
rect 37476 36650 37504 37198
rect 37464 36644 37516 36650
rect 37464 36586 37516 36592
rect 36728 36576 36780 36582
rect 36728 36518 36780 36524
rect 36176 36372 36228 36378
rect 36176 36314 36228 36320
rect 34796 36168 34848 36174
rect 34796 36110 34848 36116
rect 34428 31884 34480 31890
rect 34428 31826 34480 31832
rect 33692 31816 33744 31822
rect 33692 31758 33744 31764
rect 30656 31340 30708 31346
rect 30656 31282 30708 31288
rect 30012 30660 30064 30666
rect 30012 30602 30064 30608
rect 33600 30252 33652 30258
rect 33600 30194 33652 30200
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 29920 27124 29972 27130
rect 29920 27066 29972 27072
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 29736 22500 29788 22506
rect 29736 22442 29788 22448
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27528 19236 27580 19242
rect 27528 19178 27580 19184
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25320 17604 25372 17610
rect 25320 17546 25372 17552
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24780 16250 24808 16526
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 24124 15438 24176 15444
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 24136 14890 24164 15438
rect 24596 15422 24716 15450
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 24596 14521 24624 15422
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24582 14512 24638 14521
rect 24688 14482 24716 15302
rect 24582 14447 24638 14456
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23860 14074 23888 14214
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23768 12442 23796 13194
rect 23952 12782 23980 13194
rect 24228 12986 24256 13806
rect 24596 13394 24624 13874
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23584 5710 23612 10406
rect 24688 6186 24716 13806
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12850 24808 13126
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24872 12442 24900 16118
rect 25700 16114 25728 16934
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 25148 13852 25176 15438
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25240 14550 25268 14758
rect 25332 14550 25360 14894
rect 25228 14544 25280 14550
rect 25228 14486 25280 14492
rect 25320 14544 25372 14550
rect 25320 14486 25372 14492
rect 25700 14498 25728 15506
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 25240 14006 25268 14486
rect 25332 14074 25360 14486
rect 25700 14482 26004 14498
rect 25700 14476 26016 14482
rect 25700 14470 25964 14476
rect 25700 14414 25728 14470
rect 26332 14476 26384 14482
rect 25964 14418 26016 14424
rect 26252 14436 26332 14464
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 26252 14346 26280 14436
rect 26332 14418 26384 14424
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 25872 14272 25924 14278
rect 25872 14214 25924 14220
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25148 13824 25268 13852
rect 25240 13326 25268 13824
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 25240 9518 25268 13262
rect 25320 13184 25372 13190
rect 25320 13126 25372 13132
rect 25332 12714 25360 13126
rect 25608 12986 25636 13262
rect 25792 13258 25820 13874
rect 25884 13530 25912 14214
rect 26528 14074 26556 14894
rect 27816 14482 27844 20878
rect 30024 18970 30052 29990
rect 33324 29028 33376 29034
rect 33324 28970 33376 28976
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 30472 27872 30524 27878
rect 30472 27814 30524 27820
rect 30484 21078 30512 27814
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 31772 21146 31800 25842
rect 32784 24682 32812 28494
rect 33336 24818 33364 28970
rect 33612 26042 33640 30194
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33324 24812 33376 24818
rect 33324 24754 33376 24760
rect 32772 24676 32824 24682
rect 32772 24618 32824 24624
rect 33416 24608 33468 24614
rect 33416 24550 33468 24556
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 31852 21956 31904 21962
rect 31852 21898 31904 21904
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 30472 21072 30524 21078
rect 30472 21014 30524 21020
rect 31864 20058 31892 21898
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 30012 18964 30064 18970
rect 30012 18906 30064 18912
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29748 16114 29776 16390
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 31680 15094 31708 15846
rect 31668 15088 31720 15094
rect 31668 15030 31720 15036
rect 27804 14476 27856 14482
rect 27804 14418 27856 14424
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26252 13734 26280 13874
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 25780 13252 25832 13258
rect 25780 13194 25832 13200
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 26252 12850 26280 13670
rect 26988 13530 27016 14350
rect 29932 14006 29960 14350
rect 32416 14346 32444 22374
rect 33428 16726 33456 24550
rect 33704 24138 33732 31758
rect 33784 29640 33836 29646
rect 33784 29582 33836 29588
rect 33796 28762 33824 29582
rect 33784 28756 33836 28762
rect 33784 28698 33836 28704
rect 33968 25152 34020 25158
rect 33968 25094 34020 25100
rect 33692 24132 33744 24138
rect 33692 24074 33744 24080
rect 33980 23118 34008 25094
rect 33968 23112 34020 23118
rect 33968 23054 34020 23060
rect 34808 23050 34836 36110
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35348 35080 35400 35086
rect 35348 35022 35400 35028
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30938 35388 35022
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 35348 30932 35400 30938
rect 35348 30874 35400 30880
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35452 29850 35480 32370
rect 36740 30326 36768 36518
rect 38028 36174 38056 39200
rect 39316 36922 39344 39200
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 38016 36168 38068 36174
rect 38016 36110 38068 36116
rect 37280 36032 37332 36038
rect 37280 35974 37332 35980
rect 37292 30802 37320 35974
rect 38200 34944 38252 34950
rect 38200 34886 38252 34892
rect 38212 34785 38240 34886
rect 38198 34776 38254 34785
rect 38198 34711 38254 34720
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 38304 33425 38332 33458
rect 38290 33416 38346 33425
rect 38290 33351 38346 33360
rect 38108 33312 38160 33318
rect 38108 33254 38160 33260
rect 37280 30796 37332 30802
rect 37280 30738 37332 30744
rect 36728 30320 36780 30326
rect 36728 30262 36780 30268
rect 35440 29844 35492 29850
rect 35440 29786 35492 29792
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 38120 28082 38148 33254
rect 38200 32224 38252 32230
rect 38200 32166 38252 32172
rect 38212 32065 38240 32166
rect 38198 32056 38254 32065
rect 38198 31991 38254 32000
rect 38200 30048 38252 30054
rect 38198 30016 38200 30025
rect 38252 30016 38254 30025
rect 38198 29951 38254 29960
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38304 28665 38332 29106
rect 38290 28656 38346 28665
rect 38290 28591 38346 28600
rect 38108 28076 38160 28082
rect 38108 28018 38160 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 36728 27464 36780 27470
rect 36728 27406 36780 27412
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 36740 26042 36768 27406
rect 38200 27328 38252 27334
rect 38198 27296 38200 27305
rect 38252 27296 38254 27305
rect 38198 27231 38254 27240
rect 36728 26036 36780 26042
rect 36728 25978 36780 25984
rect 36912 25900 36964 25906
rect 36912 25842 36964 25848
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36924 24818 36952 25842
rect 38292 25288 38344 25294
rect 38290 25256 38292 25265
rect 38344 25256 38346 25265
rect 38290 25191 38346 25200
rect 35532 24812 35584 24818
rect 35532 24754 35584 24760
rect 36912 24812 36964 24818
rect 36912 24754 36964 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 23044 34848 23050
rect 34796 22986 34848 22992
rect 34060 22976 34112 22982
rect 34060 22918 34112 22924
rect 33784 22228 33836 22234
rect 33784 22170 33836 22176
rect 33796 21690 33824 22170
rect 33784 21684 33836 21690
rect 33784 21626 33836 21632
rect 34072 19446 34100 22918
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35544 20874 35572 24754
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 37004 24064 37056 24070
rect 37004 24006 37056 24012
rect 37016 22642 37044 24006
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 37004 22636 37056 22642
rect 37004 22578 37056 22584
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 38120 21146 38148 21490
rect 38108 21140 38160 21146
rect 38108 21082 38160 21088
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 35532 20868 35584 20874
rect 35532 20810 35584 20816
rect 38304 20505 38332 20878
rect 38290 20496 38346 20505
rect 38290 20431 38346 20440
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34060 19440 34112 19446
rect 34060 19382 34112 19388
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 38292 17196 38344 17202
rect 38292 17138 38344 17144
rect 38304 17105 38332 17138
rect 38290 17096 38346 17105
rect 38290 17031 38346 17040
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33416 16720 33468 16726
rect 33416 16662 33468 16668
rect 36084 16108 36136 16114
rect 36084 16050 36136 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 36096 15162 36124 16050
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 36084 15156 36136 15162
rect 36084 15098 36136 15104
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33612 14618 33640 14962
rect 37188 14952 37240 14958
rect 37188 14894 37240 14900
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 32404 14340 32456 14346
rect 32404 14282 32456 14288
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27988 13456 28040 13462
rect 27988 13398 28040 13404
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 25412 12844 25464 12850
rect 25412 12786 25464 12792
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 25320 12708 25372 12714
rect 25320 12650 25372 12656
rect 25424 12238 25452 12786
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25424 8634 25452 12174
rect 27264 10674 27292 13126
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25410 7848 25466 7857
rect 25410 7783 25466 7792
rect 25424 6866 25452 7783
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23296 5568 23348 5574
rect 23296 5510 23348 5516
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 23308 2446 23336 5510
rect 24780 2446 24808 5510
rect 27172 2446 27200 10610
rect 28000 8090 28028 13398
rect 28264 12776 28316 12782
rect 28264 12718 28316 12724
rect 28276 10062 28304 12718
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 33968 12368 34020 12374
rect 33968 12310 34020 12316
rect 28356 11076 28408 11082
rect 28356 11018 28408 11024
rect 28368 10062 28396 11018
rect 33980 10266 34008 12310
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 37200 11354 37228 14894
rect 38016 14816 38068 14822
rect 38016 14758 38068 14764
rect 38028 12850 38056 14758
rect 38292 14408 38344 14414
rect 38290 14376 38292 14385
rect 38344 14376 38346 14385
rect 38290 14311 38346 14320
rect 38016 12844 38068 12850
rect 38016 12786 38068 12792
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 37188 11348 37240 11354
rect 37188 11290 37240 11296
rect 34152 10532 34204 10538
rect 34152 10474 34204 10480
rect 33968 10260 34020 10266
rect 33968 10202 34020 10208
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28356 10056 28408 10062
rect 28356 9998 28408 10004
rect 29644 9920 29696 9926
rect 29644 9862 29696 9868
rect 31668 9920 31720 9926
rect 31668 9862 31720 9868
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27540 2582 27568 6734
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28184 3058 28212 4422
rect 28172 3052 28224 3058
rect 28172 2994 28224 3000
rect 28644 2650 28672 8910
rect 29656 5234 29684 9862
rect 31680 9586 31708 9862
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 33968 8492 34020 8498
rect 33968 8434 34020 8440
rect 33600 7880 33652 7886
rect 33600 7822 33652 7828
rect 32864 6316 32916 6322
rect 32864 6258 32916 6264
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 27528 2576 27580 2582
rect 27528 2518 27580 2524
rect 30208 2514 30236 2790
rect 32876 2582 32904 6258
rect 33612 2650 33640 7822
rect 33980 3738 34008 8434
rect 34164 6798 34192 10474
rect 36360 10464 36412 10470
rect 36360 10406 36412 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 36372 7410 36400 10406
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37200 8090 37228 9998
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 38028 8974 38056 9318
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 37188 8084 37240 8090
rect 37188 8026 37240 8032
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 38016 7200 38068 7206
rect 38016 7142 38068 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 37004 6656 37056 6662
rect 37004 6598 37056 6604
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 33968 3732 34020 3738
rect 33968 3674 34020 3680
rect 35636 3194 35664 6258
rect 36912 5024 36964 5030
rect 36912 4966 36964 4972
rect 35624 3188 35676 3194
rect 35624 3130 35676 3136
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 32864 2576 32916 2582
rect 32864 2518 32916 2524
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 36924 2446 36952 4966
rect 37016 3058 37044 6598
rect 38028 4622 38056 7142
rect 38120 6458 38148 12174
rect 38292 11144 38344 11150
rect 38292 11086 38344 11092
rect 38304 10985 38332 11086
rect 38290 10976 38346 10985
rect 38290 10911 38346 10920
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38108 6452 38160 6458
rect 38108 6394 38160 6400
rect 38292 6316 38344 6322
rect 38292 6258 38344 6264
rect 38304 6225 38332 6258
rect 38290 6216 38346 6225
rect 38290 6151 38346 6160
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 38212 4185 38240 4422
rect 38198 4176 38254 4185
rect 38198 4111 38254 4120
rect 38292 3528 38344 3534
rect 38292 3470 38344 3476
rect 37004 3052 37056 3058
rect 37004 2994 37056 3000
rect 38200 2848 38252 2854
rect 38304 2825 38332 3470
rect 39304 2984 39356 2990
rect 39304 2926 39356 2932
rect 38200 2790 38252 2796
rect 38290 2816 38346 2825
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36912 2440 36964 2446
rect 36912 2382 36964 2388
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 4540 800 4568 2314
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 800 5856 2246
rect 7116 800 7144 2382
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 9048 800 9076 2246
rect 10336 800 10364 2246
rect 11624 800 11652 2382
rect 13556 800 13584 2382
rect 14844 800 14872 2382
rect 16776 800 16804 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 18064 800 18092 2246
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 21284 800 21312 2382
rect 22572 800 22600 2382
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 23860 800 23888 2246
rect 25792 800 25820 2246
rect 27080 800 27108 2314
rect 29012 800 29040 2382
rect 30300 800 30328 2382
rect 31576 2304 31628 2310
rect 31576 2246 31628 2252
rect 31588 800 31616 2246
rect 33520 800 33548 2382
rect 34808 800 34836 2382
rect 36096 800 36124 2382
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38028 800 38056 2246
rect 38212 1465 38240 2790
rect 38290 2751 38346 2760
rect 38198 1456 38254 1465
rect 38198 1391 38254 1400
rect 39316 800 39344 2926
rect 18 200 74 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 4526 200 4582 800
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 9034 200 9090 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23846 200 23902 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 31574 200 31630 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 36082 200 36138 800
rect 38014 200 38070 800
rect 39302 200 39358 800
<< via2 >>
rect 3146 38120 3202 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2778 36760 2834 36816
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 1766 33360 1822 33416
rect 1766 32000 1822 32056
rect 1766 30676 1768 30696
rect 1768 30676 1820 30696
rect 1820 30676 1822 30696
rect 1766 30640 1822 30676
rect 1766 28600 1822 28656
rect 1766 27240 1822 27296
rect 1766 25236 1768 25256
rect 1768 25236 1820 25256
rect 1820 25236 1822 25256
rect 1766 25200 1822 25236
rect 1766 23840 1822 23896
rect 1766 22480 1822 22536
rect 1766 20440 1822 20496
rect 1766 19080 1822 19136
rect 1766 15680 1822 15736
rect 1858 13368 1914 13424
rect 1766 12280 1822 12336
rect 1674 10920 1730 10976
rect 1674 8628 1730 8664
rect 1674 8608 1676 8628
rect 1676 8608 1728 8628
rect 1728 8608 1730 8628
rect 2318 18128 2374 18184
rect 2962 21800 3018 21856
rect 2778 17720 2834 17776
rect 1950 10804 2006 10840
rect 1950 10784 1952 10804
rect 1952 10784 2004 10804
rect 2004 10784 2006 10804
rect 2134 10104 2190 10160
rect 1950 8200 2006 8256
rect 2778 11736 2834 11792
rect 2778 11192 2834 11248
rect 2962 13776 3018 13832
rect 3238 14320 3294 14376
rect 2778 9424 2834 9480
rect 3054 9424 3110 9480
rect 1766 4800 1822 4856
rect 3606 18536 3662 18592
rect 3790 19916 3846 19952
rect 3790 19896 3792 19916
rect 3792 19896 3844 19916
rect 3844 19896 3846 19916
rect 3606 16224 3662 16280
rect 3790 15036 3792 15056
rect 3792 15036 3844 15056
rect 3844 15036 3846 15056
rect 3790 15000 3846 15036
rect 3422 12960 3478 13016
rect 3790 12280 3846 12336
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 5722 31728 5778 31784
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4710 22072 4766 22128
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4526 20576 4582 20632
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4434 17756 4436 17776
rect 4436 17756 4488 17776
rect 4488 17756 4490 17776
rect 4434 17720 4490 17756
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4526 14456 4582 14512
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4342 12860 4344 12880
rect 4344 12860 4396 12880
rect 4396 12860 4398 12880
rect 4342 12824 4398 12860
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4434 12280 4490 12336
rect 4894 20576 4950 20632
rect 4894 19488 4950 19544
rect 5078 19624 5134 19680
rect 4894 17076 4896 17096
rect 4896 17076 4948 17096
rect 4948 17076 4950 17096
rect 4894 17040 4950 17076
rect 4710 13096 4766 13152
rect 3698 11872 3754 11928
rect 3330 7964 3332 7984
rect 3332 7964 3384 7984
rect 3384 7964 3386 7984
rect 3330 7928 3386 7964
rect 3146 6568 3202 6624
rect 3238 6296 3294 6352
rect 3698 10512 3754 10568
rect 3974 12144 4030 12200
rect 3790 6160 3846 6216
rect 3698 5480 3754 5536
rect 4618 12008 4674 12064
rect 4526 11872 4582 11928
rect 4618 11772 4620 11792
rect 4620 11772 4672 11792
rect 4672 11772 4674 11792
rect 4618 11736 4674 11772
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4158 10920 4214 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4526 9424 4582 9480
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4618 7520 4674 7576
rect 4986 9152 5042 9208
rect 5170 12688 5226 12744
rect 5446 20576 5502 20632
rect 5630 20712 5686 20768
rect 5630 19780 5686 19816
rect 5630 19760 5632 19780
rect 5632 19760 5684 19780
rect 5684 19760 5686 19780
rect 5446 19352 5502 19408
rect 5262 12552 5318 12608
rect 5170 11636 5172 11656
rect 5172 11636 5224 11656
rect 5224 11636 5226 11656
rect 5170 11600 5226 11636
rect 5446 13776 5502 13832
rect 5446 12688 5502 12744
rect 4894 8472 4950 8528
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4802 7520 4858 7576
rect 4158 6840 4214 6896
rect 4802 6704 4858 6760
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4342 5364 4398 5400
rect 4342 5344 4344 5364
rect 4344 5344 4396 5364
rect 4396 5344 4398 5364
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4250 4684 4306 4720
rect 4250 4664 4252 4684
rect 4252 4664 4304 4684
rect 4304 4664 4306 4684
rect 5078 8628 5134 8664
rect 5078 8608 5080 8628
rect 5080 8608 5132 8628
rect 5132 8608 5134 8628
rect 4986 7384 5042 7440
rect 4986 5616 5042 5672
rect 4526 4020 4528 4040
rect 4528 4020 4580 4040
rect 4580 4020 4582 4040
rect 4526 3984 4582 4020
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5446 6976 5502 7032
rect 5354 6432 5410 6488
rect 5354 5908 5410 5944
rect 5354 5888 5356 5908
rect 5356 5888 5408 5908
rect 5408 5888 5410 5908
rect 3974 2760 4030 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6182 21936 6238 21992
rect 6550 21936 6606 21992
rect 6642 18692 6698 18728
rect 6642 18672 6644 18692
rect 6644 18672 6696 18692
rect 6696 18672 6698 18692
rect 5998 6860 6054 6896
rect 5998 6840 6000 6860
rect 6000 6840 6052 6860
rect 6052 6840 6054 6860
rect 6274 9832 6330 9888
rect 6642 13640 6698 13696
rect 6550 9288 6606 9344
rect 7194 18284 7250 18320
rect 7194 18264 7196 18284
rect 7196 18264 7248 18284
rect 7248 18264 7250 18284
rect 7102 17584 7158 17640
rect 7562 20712 7618 20768
rect 7194 14184 7250 14240
rect 7010 11892 7066 11928
rect 7010 11872 7012 11892
rect 7012 11872 7064 11892
rect 7064 11872 7066 11892
rect 7102 10104 7158 10160
rect 6826 8880 6882 8936
rect 8022 19780 8078 19816
rect 8022 19760 8024 19780
rect 8024 19760 8076 19780
rect 8076 19760 8078 19780
rect 7838 18300 7840 18320
rect 7840 18300 7892 18320
rect 7892 18300 7894 18320
rect 7838 18264 7894 18300
rect 9126 20340 9128 20360
rect 9128 20340 9180 20360
rect 9180 20340 9182 20360
rect 8482 19896 8538 19952
rect 9126 20304 9182 20340
rect 8666 19488 8722 19544
rect 8298 18536 8354 18592
rect 8114 16940 8116 16960
rect 8116 16940 8168 16960
rect 8168 16940 8170 16960
rect 8114 16904 8170 16940
rect 8022 14320 8078 14376
rect 7838 13776 7894 13832
rect 7654 11600 7710 11656
rect 8114 12316 8116 12336
rect 8116 12316 8168 12336
rect 8168 12316 8170 12336
rect 8114 12280 8170 12316
rect 7930 8084 7986 8120
rect 7930 8064 7932 8084
rect 7932 8064 7984 8084
rect 7984 8064 7986 8084
rect 7930 6840 7986 6896
rect 8390 16224 8446 16280
rect 8574 18692 8630 18728
rect 8574 18672 8576 18692
rect 8576 18672 8628 18692
rect 8628 18672 8630 18692
rect 9034 19236 9090 19272
rect 9034 19216 9036 19236
rect 9036 19216 9088 19236
rect 9088 19216 9090 19236
rect 9126 19116 9128 19136
rect 9128 19116 9180 19136
rect 9180 19116 9182 19136
rect 9126 19080 9182 19116
rect 9126 17856 9182 17912
rect 9310 19388 9312 19408
rect 9312 19388 9364 19408
rect 9364 19388 9366 19408
rect 9310 19352 9366 19388
rect 9770 21936 9826 21992
rect 9862 21256 9918 21312
rect 10046 21120 10102 21176
rect 9862 20984 9918 21040
rect 9402 17740 9458 17776
rect 9402 17720 9404 17740
rect 9404 17720 9456 17740
rect 9456 17720 9458 17740
rect 9494 16940 9496 16960
rect 9496 16940 9548 16960
rect 9548 16940 9550 16960
rect 9494 16904 9550 16940
rect 8574 15272 8630 15328
rect 9310 14456 9366 14512
rect 8390 12980 8446 13016
rect 8390 12960 8392 12980
rect 8392 12960 8444 12980
rect 8444 12960 8446 12980
rect 8942 13640 8998 13696
rect 8574 11736 8630 11792
rect 8298 8880 8354 8936
rect 9954 20848 10010 20904
rect 9954 20440 10010 20496
rect 10506 20848 10562 20904
rect 10414 20440 10470 20496
rect 10782 19896 10838 19952
rect 10046 18400 10102 18456
rect 11058 20712 11114 20768
rect 11334 20712 11390 20768
rect 10506 19352 10562 19408
rect 10782 19372 10838 19408
rect 10782 19352 10784 19372
rect 10784 19352 10836 19372
rect 10836 19352 10838 19372
rect 10322 17584 10378 17640
rect 10138 15272 10194 15328
rect 9678 13912 9734 13968
rect 9126 12008 9182 12064
rect 9494 12844 9550 12880
rect 9494 12824 9496 12844
rect 9496 12824 9548 12844
rect 9548 12824 9550 12844
rect 9126 10140 9128 10160
rect 9128 10140 9180 10160
rect 9180 10140 9182 10160
rect 9126 10104 9182 10140
rect 8942 9288 8998 9344
rect 10230 13776 10286 13832
rect 10782 18264 10838 18320
rect 11334 20304 11390 20360
rect 10690 16632 10746 16688
rect 10598 14320 10654 14376
rect 10322 13504 10378 13560
rect 9862 11192 9918 11248
rect 9678 10104 9734 10160
rect 9586 9832 9642 9888
rect 10046 12960 10102 13016
rect 10046 12164 10102 12200
rect 10046 12144 10048 12164
rect 10048 12144 10100 12164
rect 10100 12144 10102 12164
rect 11334 18264 11390 18320
rect 11794 20984 11850 21040
rect 12254 20848 12310 20904
rect 11610 17992 11666 18048
rect 12898 22072 12954 22128
rect 12622 21120 12678 21176
rect 12162 19216 12218 19272
rect 11978 19080 12034 19136
rect 11978 18808 12034 18864
rect 11426 16088 11482 16144
rect 10782 14184 10838 14240
rect 10598 11872 10654 11928
rect 11702 15272 11758 15328
rect 11242 15136 11298 15192
rect 12070 13776 12126 13832
rect 12070 13640 12126 13696
rect 11978 10104 12034 10160
rect 12346 19080 12402 19136
rect 12346 18148 12402 18184
rect 12346 18128 12348 18148
rect 12348 18128 12400 18148
rect 12400 18128 12402 18148
rect 12714 19080 12770 19136
rect 12622 18944 12678 19000
rect 12346 13640 12402 13696
rect 12622 12552 12678 12608
rect 12622 12280 12678 12336
rect 12530 12180 12532 12200
rect 12532 12180 12584 12200
rect 12584 12180 12586 12200
rect 12530 12144 12586 12180
rect 12898 11736 12954 11792
rect 14278 23060 14280 23080
rect 14280 23060 14332 23080
rect 14332 23060 14334 23080
rect 14278 23024 14334 23060
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 15106 21020 15108 21040
rect 15108 21020 15160 21040
rect 15160 21020 15162 21040
rect 15106 20984 15162 21020
rect 15290 20848 15346 20904
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 17866 22072 17922 22128
rect 16486 21972 16488 21992
rect 16488 21972 16540 21992
rect 16540 21972 16542 21992
rect 16486 21936 16542 21972
rect 15566 18400 15622 18456
rect 13634 12860 13636 12880
rect 13636 12860 13688 12880
rect 13688 12860 13690 12880
rect 13634 12824 13690 12860
rect 13082 10532 13138 10568
rect 13082 10512 13084 10532
rect 13084 10512 13136 10532
rect 13136 10512 13138 10532
rect 15382 16632 15438 16688
rect 14278 15136 14334 15192
rect 14186 12824 14242 12880
rect 15566 14612 15622 14648
rect 15566 14592 15568 14612
rect 15568 14592 15620 14612
rect 15620 14592 15622 14612
rect 15474 13504 15530 13560
rect 17130 18808 17186 18864
rect 18142 19624 18198 19680
rect 17406 14592 17462 14648
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19522 22092 19578 22128
rect 19522 22072 19524 22092
rect 19524 22072 19576 22092
rect 19576 22072 19578 22092
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19246 19624 19302 19680
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 18970 15000 19026 15056
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 18142 13504 18198 13560
rect 18510 12960 18566 13016
rect 18510 11736 18566 11792
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 37002 38120 37058 38176
rect 36910 36760 36966 36816
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 24582 14456 24638 14512
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 38198 34720 38254 34776
rect 38290 33360 38346 33416
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 38198 32000 38254 32056
rect 38198 29996 38200 30016
rect 38200 29996 38252 30016
rect 38252 29996 38254 30016
rect 38198 29960 38254 29996
rect 38290 28600 38346 28656
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 38198 27276 38200 27296
rect 38200 27276 38252 27296
rect 38252 27276 38254 27296
rect 38198 27240 38254 27276
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 38290 25236 38292 25256
rect 38292 25236 38344 25256
rect 38344 25236 38346 25256
rect 38290 25200 38346 25236
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 38290 23840 38346 23896
rect 38290 21800 38346 21856
rect 38290 20440 38346 20496
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 38290 17040 38346 17096
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 38198 15680 38254 15736
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 25410 7792 25466 7848
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38290 14356 38292 14376
rect 38292 14356 38344 14376
rect 38344 14356 38346 14376
rect 38290 14320 38346 14356
rect 38198 12280 38254 12336
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 10920 38346 10976
rect 38198 8880 38254 8936
rect 38290 7520 38346 7576
rect 38290 6160 38346 6216
rect 38198 4120 38254 4176
rect 4066 1400 4122 1456
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38290 2760 38346 2816
rect 38198 1400 38254 1456
<< metal3 >>
rect 200 38178 800 38208
rect 3141 38178 3207 38181
rect 200 38176 3207 38178
rect 200 38120 3146 38176
rect 3202 38120 3207 38176
rect 200 38118 3207 38120
rect 200 38088 800 38118
rect 3141 38115 3207 38118
rect 36997 38178 37063 38181
rect 39200 38178 39800 38208
rect 36997 38176 39800 38178
rect 36997 38120 37002 38176
rect 37058 38120 39800 38176
rect 36997 38118 39800 38120
rect 36997 38115 37063 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 2773 36818 2839 36821
rect 200 36816 2839 36818
rect 200 36760 2778 36816
rect 2834 36760 2839 36816
rect 200 36758 2839 36760
rect 200 36728 800 36758
rect 2773 36755 2839 36758
rect 36905 36818 36971 36821
rect 39200 36818 39800 36848
rect 36905 36816 39800 36818
rect 36905 36760 36910 36816
rect 36966 36760 39800 36816
rect 36905 36758 39800 36760
rect 36905 36755 36971 36758
rect 39200 36728 39800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35368 800 35488
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 38193 34778 38259 34781
rect 39200 34778 39800 34808
rect 38193 34776 39800 34778
rect 38193 34720 38198 34776
rect 38254 34720 39800 34776
rect 38193 34718 39800 34720
rect 38193 34715 38259 34718
rect 39200 34688 39800 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 200 33418 800 33448
rect 1761 33418 1827 33421
rect 200 33416 1827 33418
rect 200 33360 1766 33416
rect 1822 33360 1827 33416
rect 200 33358 1827 33360
rect 200 33328 800 33358
rect 1761 33355 1827 33358
rect 38285 33418 38351 33421
rect 39200 33418 39800 33448
rect 38285 33416 39800 33418
rect 38285 33360 38290 33416
rect 38346 33360 39800 33416
rect 38285 33358 39800 33360
rect 38285 33355 38351 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38193 32058 38259 32061
rect 39200 32058 39800 32088
rect 38193 32056 39800 32058
rect 38193 32000 38198 32056
rect 38254 32000 39800 32056
rect 38193 31998 39800 32000
rect 38193 31995 38259 31998
rect 39200 31968 39800 31998
rect 5717 31788 5783 31789
rect 5717 31784 5764 31788
rect 5828 31786 5834 31788
rect 5717 31728 5722 31784
rect 5717 31724 5764 31728
rect 5828 31726 5874 31786
rect 5828 31724 5834 31726
rect 5717 31723 5783 31724
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 38193 30018 38259 30021
rect 39200 30018 39800 30048
rect 38193 30016 39800 30018
rect 38193 29960 38198 30016
rect 38254 29960 39800 30016
rect 38193 29958 39800 29960
rect 38193 29955 38259 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 39800 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1761 28658 1827 28661
rect 200 28656 1827 28658
rect 200 28600 1766 28656
rect 1822 28600 1827 28656
rect 200 28598 1827 28600
rect 200 28568 800 28598
rect 1761 28595 1827 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 38193 27298 38259 27301
rect 39200 27298 39800 27328
rect 38193 27296 39800 27298
rect 38193 27240 38198 27296
rect 38254 27240 39800 27296
rect 38193 27238 39800 27240
rect 38193 27235 38259 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 38285 25258 38351 25261
rect 39200 25258 39800 25288
rect 38285 25256 39800 25258
rect 38285 25200 38290 25256
rect 38346 25200 39800 25256
rect 38285 25198 39800 25200
rect 38285 25195 38351 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1761 23898 1827 23901
rect 200 23896 1827 23898
rect 200 23840 1766 23896
rect 1822 23840 1827 23896
rect 200 23838 1827 23840
rect 200 23808 800 23838
rect 1761 23835 1827 23838
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 7966 23020 7972 23084
rect 8036 23082 8042 23084
rect 14273 23082 14339 23085
rect 8036 23080 14339 23082
rect 8036 23024 14278 23080
rect 14334 23024 14339 23080
rect 8036 23022 14339 23024
rect 8036 23020 8042 23022
rect 14273 23019 14339 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 4705 22130 4771 22133
rect 5206 22130 5212 22132
rect 4705 22128 5212 22130
rect 4705 22072 4710 22128
rect 4766 22072 5212 22128
rect 4705 22070 5212 22072
rect 4705 22067 4771 22070
rect 5206 22068 5212 22070
rect 5276 22130 5282 22132
rect 12893 22130 12959 22133
rect 5276 22128 12959 22130
rect 5276 22072 12898 22128
rect 12954 22072 12959 22128
rect 5276 22070 12959 22072
rect 5276 22068 5282 22070
rect 12893 22067 12959 22070
rect 17861 22130 17927 22133
rect 19517 22130 19583 22133
rect 17861 22128 19583 22130
rect 17861 22072 17866 22128
rect 17922 22072 19522 22128
rect 19578 22072 19583 22128
rect 17861 22070 19583 22072
rect 17861 22067 17927 22070
rect 19517 22067 19583 22070
rect 6177 21994 6243 21997
rect 6545 21994 6611 21997
rect 6177 21992 6611 21994
rect 6177 21936 6182 21992
rect 6238 21936 6550 21992
rect 6606 21936 6611 21992
rect 6177 21934 6611 21936
rect 6177 21931 6243 21934
rect 6545 21931 6611 21934
rect 9765 21994 9831 21997
rect 16481 21994 16547 21997
rect 9765 21992 16547 21994
rect 9765 21936 9770 21992
rect 9826 21936 16486 21992
rect 16542 21936 16547 21992
rect 9765 21934 16547 21936
rect 9765 21931 9831 21934
rect 16481 21931 16547 21934
rect 2814 21796 2820 21860
rect 2884 21858 2890 21860
rect 2957 21858 3023 21861
rect 2884 21856 3023 21858
rect 2884 21800 2962 21856
rect 3018 21800 3023 21856
rect 2884 21798 3023 21800
rect 2884 21796 2890 21798
rect 2957 21795 3023 21798
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 9857 21314 9923 21317
rect 9814 21312 9923 21314
rect 9814 21256 9862 21312
rect 9918 21256 9923 21312
rect 9814 21251 9923 21256
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 9814 21045 9874 21251
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 10041 21178 10107 21181
rect 12617 21178 12683 21181
rect 10041 21176 12683 21178
rect 10041 21120 10046 21176
rect 10102 21120 12622 21176
rect 12678 21120 12683 21176
rect 10041 21118 12683 21120
rect 10041 21115 10107 21118
rect 12617 21115 12683 21118
rect 9814 21040 9923 21045
rect 9814 20984 9862 21040
rect 9918 20984 9923 21040
rect 9814 20982 9923 20984
rect 9857 20979 9923 20982
rect 11789 21042 11855 21045
rect 15101 21042 15167 21045
rect 11789 21040 15167 21042
rect 11789 20984 11794 21040
rect 11850 20984 15106 21040
rect 15162 20984 15167 21040
rect 11789 20982 15167 20984
rect 11789 20979 11855 20982
rect 15101 20979 15167 20982
rect 9949 20906 10015 20909
rect 10501 20906 10567 20909
rect 9949 20904 10567 20906
rect 9949 20848 9954 20904
rect 10010 20848 10506 20904
rect 10562 20848 10567 20904
rect 9949 20846 10567 20848
rect 9949 20843 10015 20846
rect 10501 20843 10567 20846
rect 12249 20906 12315 20909
rect 15285 20906 15351 20909
rect 12249 20904 15351 20906
rect 12249 20848 12254 20904
rect 12310 20848 15290 20904
rect 15346 20848 15351 20904
rect 12249 20846 15351 20848
rect 12249 20843 12315 20846
rect 15285 20843 15351 20846
rect 5625 20772 5691 20773
rect 5574 20770 5580 20772
rect 5534 20710 5580 20770
rect 5644 20768 5691 20772
rect 5686 20712 5691 20768
rect 5574 20708 5580 20710
rect 5644 20708 5691 20712
rect 5625 20707 5691 20708
rect 7557 20772 7623 20773
rect 11053 20772 11119 20773
rect 11329 20772 11395 20773
rect 7557 20768 7604 20772
rect 7668 20770 7674 20772
rect 7557 20712 7562 20768
rect 7557 20708 7604 20712
rect 7668 20710 7714 20770
rect 11053 20768 11100 20772
rect 11164 20770 11170 20772
rect 11053 20712 11058 20768
rect 7668 20708 7674 20710
rect 11053 20708 11100 20712
rect 11164 20710 11210 20770
rect 11164 20708 11170 20710
rect 11278 20708 11284 20772
rect 11348 20770 11395 20772
rect 11348 20768 11440 20770
rect 11390 20712 11440 20768
rect 11348 20710 11440 20712
rect 11348 20708 11395 20710
rect 7557 20707 7623 20708
rect 11053 20707 11119 20708
rect 11329 20707 11395 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4521 20634 4587 20637
rect 4889 20634 4955 20637
rect 5441 20634 5507 20637
rect 4521 20632 5507 20634
rect 4521 20576 4526 20632
rect 4582 20576 4894 20632
rect 4950 20576 5446 20632
rect 5502 20576 5507 20632
rect 4521 20574 5507 20576
rect 4521 20571 4587 20574
rect 4889 20571 4955 20574
rect 5441 20571 5507 20574
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 9949 20498 10015 20501
rect 10409 20498 10475 20501
rect 9949 20496 10475 20498
rect 9949 20440 9954 20496
rect 10010 20440 10414 20496
rect 10470 20440 10475 20496
rect 9949 20438 10475 20440
rect 9949 20435 10015 20438
rect 10409 20435 10475 20438
rect 38285 20498 38351 20501
rect 39200 20498 39800 20528
rect 38285 20496 39800 20498
rect 38285 20440 38290 20496
rect 38346 20440 39800 20496
rect 38285 20438 39800 20440
rect 38285 20435 38351 20438
rect 39200 20408 39800 20438
rect 9121 20362 9187 20365
rect 11329 20362 11395 20365
rect 9121 20360 11395 20362
rect 9121 20304 9126 20360
rect 9182 20304 11334 20360
rect 11390 20304 11395 20360
rect 9121 20302 11395 20304
rect 9121 20299 9187 20302
rect 11329 20299 11395 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 3785 19954 3851 19957
rect 8477 19954 8543 19957
rect 3785 19952 8543 19954
rect 3785 19896 3790 19952
rect 3846 19896 8482 19952
rect 8538 19896 8543 19952
rect 3785 19894 8543 19896
rect 3785 19891 3851 19894
rect 8477 19891 8543 19894
rect 10777 19954 10843 19957
rect 10910 19954 10916 19956
rect 10777 19952 10916 19954
rect 10777 19896 10782 19952
rect 10838 19896 10916 19952
rect 10777 19894 10916 19896
rect 10777 19891 10843 19894
rect 10910 19892 10916 19894
rect 10980 19892 10986 19956
rect 5625 19818 5691 19821
rect 8017 19818 8083 19821
rect 5625 19816 8083 19818
rect 5625 19760 5630 19816
rect 5686 19760 8022 19816
rect 8078 19760 8083 19816
rect 5625 19758 8083 19760
rect 5625 19755 5691 19758
rect 8017 19755 8083 19758
rect 5073 19682 5139 19685
rect 18137 19682 18203 19685
rect 19241 19682 19307 19685
rect 5073 19680 19307 19682
rect 5073 19624 5078 19680
rect 5134 19624 18142 19680
rect 18198 19624 19246 19680
rect 19302 19624 19307 19680
rect 5073 19622 19307 19624
rect 5073 19619 5139 19622
rect 18137 19619 18203 19622
rect 19241 19619 19307 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4889 19546 4955 19549
rect 8661 19546 8727 19549
rect 4889 19544 8727 19546
rect 4889 19488 4894 19544
rect 4950 19488 8666 19544
rect 8722 19488 8727 19544
rect 4889 19486 8727 19488
rect 4889 19483 4955 19486
rect 8661 19483 8727 19486
rect 4838 19348 4844 19412
rect 4908 19410 4914 19412
rect 5441 19410 5507 19413
rect 9305 19410 9371 19413
rect 10501 19410 10567 19413
rect 10777 19412 10843 19413
rect 10726 19410 10732 19412
rect 4908 19408 6746 19410
rect 4908 19352 5446 19408
rect 5502 19352 6746 19408
rect 4908 19350 6746 19352
rect 4908 19348 4914 19350
rect 5441 19347 5507 19350
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 6686 19002 6746 19350
rect 9305 19408 10567 19410
rect 9305 19352 9310 19408
rect 9366 19352 10506 19408
rect 10562 19352 10567 19408
rect 9305 19350 10567 19352
rect 10686 19350 10732 19410
rect 10796 19408 10843 19412
rect 10838 19352 10843 19408
rect 9305 19347 9371 19350
rect 10501 19347 10567 19350
rect 10726 19348 10732 19350
rect 10796 19348 10843 19352
rect 10777 19347 10843 19348
rect 9029 19274 9095 19277
rect 12157 19274 12223 19277
rect 9029 19272 12223 19274
rect 9029 19216 9034 19272
rect 9090 19216 12162 19272
rect 12218 19216 12223 19272
rect 9029 19214 12223 19216
rect 9029 19211 9095 19214
rect 12157 19211 12223 19214
rect 9121 19138 9187 19141
rect 11973 19138 12039 19141
rect 9121 19136 12039 19138
rect 9121 19080 9126 19136
rect 9182 19080 11978 19136
rect 12034 19080 12039 19136
rect 9121 19078 12039 19080
rect 9121 19075 9187 19078
rect 11973 19075 12039 19078
rect 12341 19138 12407 19141
rect 12709 19138 12775 19141
rect 12341 19136 12775 19138
rect 12341 19080 12346 19136
rect 12402 19080 12714 19136
rect 12770 19080 12775 19136
rect 12341 19078 12775 19080
rect 12341 19075 12407 19078
rect 12709 19075 12775 19078
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19168
rect 34930 19007 35246 19008
rect 12617 19002 12683 19005
rect 6686 19000 12683 19002
rect 6686 18944 12622 19000
rect 12678 18944 12683 19000
rect 6686 18942 12683 18944
rect 12617 18939 12683 18942
rect 11973 18866 12039 18869
rect 17125 18866 17191 18869
rect 11973 18864 17191 18866
rect 11973 18808 11978 18864
rect 12034 18808 17130 18864
rect 17186 18808 17191 18864
rect 11973 18806 17191 18808
rect 11973 18803 12039 18806
rect 17125 18803 17191 18806
rect 6637 18730 6703 18733
rect 8569 18730 8635 18733
rect 6637 18728 8635 18730
rect 6637 18672 6642 18728
rect 6698 18672 8574 18728
rect 8630 18672 8635 18728
rect 6637 18670 8635 18672
rect 6637 18667 6703 18670
rect 8569 18667 8635 18670
rect 3601 18594 3667 18597
rect 8293 18594 8359 18597
rect 3601 18592 8359 18594
rect 3601 18536 3606 18592
rect 3662 18536 8298 18592
rect 8354 18536 8359 18592
rect 3601 18534 8359 18536
rect 3601 18531 3667 18534
rect 8293 18531 8359 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 10041 18458 10107 18461
rect 15561 18458 15627 18461
rect 10041 18456 15627 18458
rect 10041 18400 10046 18456
rect 10102 18400 15566 18456
rect 15622 18400 15627 18456
rect 10041 18398 15627 18400
rect 10041 18395 10107 18398
rect 15561 18395 15627 18398
rect 7189 18322 7255 18325
rect 7833 18322 7899 18325
rect 7189 18320 7899 18322
rect 7189 18264 7194 18320
rect 7250 18264 7838 18320
rect 7894 18264 7899 18320
rect 7189 18262 7899 18264
rect 7189 18259 7255 18262
rect 7833 18259 7899 18262
rect 10777 18322 10843 18325
rect 11329 18322 11395 18325
rect 10777 18320 11395 18322
rect 10777 18264 10782 18320
rect 10838 18264 11334 18320
rect 11390 18264 11395 18320
rect 10777 18262 11395 18264
rect 10777 18259 10843 18262
rect 11329 18259 11395 18262
rect 2313 18186 2379 18189
rect 12341 18186 12407 18189
rect 2313 18184 12407 18186
rect 2313 18128 2318 18184
rect 2374 18128 12346 18184
rect 12402 18128 12407 18184
rect 2313 18126 12407 18128
rect 2313 18123 2379 18126
rect 12341 18123 12407 18126
rect 11462 17988 11468 18052
rect 11532 18050 11538 18052
rect 11605 18050 11671 18053
rect 11532 18048 11671 18050
rect 11532 17992 11610 18048
rect 11666 17992 11671 18048
rect 11532 17990 11671 17992
rect 11532 17988 11538 17990
rect 11605 17987 11671 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 5758 17852 5764 17916
rect 5828 17914 5834 17916
rect 9121 17914 9187 17917
rect 5828 17912 9187 17914
rect 5828 17856 9126 17912
rect 9182 17856 9187 17912
rect 5828 17854 9187 17856
rect 5828 17852 5834 17854
rect 9121 17851 9187 17854
rect 200 17778 800 17808
rect 2773 17778 2839 17781
rect 200 17776 2839 17778
rect 200 17720 2778 17776
rect 2834 17720 2839 17776
rect 200 17718 2839 17720
rect 200 17688 800 17718
rect 2773 17715 2839 17718
rect 4429 17778 4495 17781
rect 9397 17778 9463 17781
rect 4429 17776 9463 17778
rect 4429 17720 4434 17776
rect 4490 17720 9402 17776
rect 9458 17720 9463 17776
rect 4429 17718 9463 17720
rect 4429 17715 4495 17718
rect 9397 17715 9463 17718
rect 7097 17642 7163 17645
rect 10317 17642 10383 17645
rect 7097 17640 10383 17642
rect 7097 17584 7102 17640
rect 7158 17584 10322 17640
rect 10378 17584 10383 17640
rect 7097 17582 10383 17584
rect 7097 17579 7163 17582
rect 10317 17579 10383 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 2078 17036 2084 17100
rect 2148 17098 2154 17100
rect 4889 17098 4955 17101
rect 2148 17096 4955 17098
rect 2148 17040 4894 17096
rect 4950 17040 4955 17096
rect 2148 17038 4955 17040
rect 2148 17036 2154 17038
rect 4889 17035 4955 17038
rect 38285 17098 38351 17101
rect 39200 17098 39800 17128
rect 38285 17096 39800 17098
rect 38285 17040 38290 17096
rect 38346 17040 39800 17096
rect 38285 17038 39800 17040
rect 38285 17035 38351 17038
rect 39200 17008 39800 17038
rect 8109 16962 8175 16965
rect 9489 16962 9555 16965
rect 8109 16960 9555 16962
rect 8109 16904 8114 16960
rect 8170 16904 9494 16960
rect 9550 16904 9555 16960
rect 8109 16902 9555 16904
rect 8109 16899 8175 16902
rect 9489 16899 9555 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 10542 16628 10548 16692
rect 10612 16690 10618 16692
rect 10685 16690 10751 16693
rect 10612 16688 10751 16690
rect 10612 16632 10690 16688
rect 10746 16632 10751 16688
rect 10612 16630 10751 16632
rect 10612 16628 10618 16630
rect 10685 16627 10751 16630
rect 15377 16690 15443 16693
rect 15510 16690 15516 16692
rect 15377 16688 15516 16690
rect 15377 16632 15382 16688
rect 15438 16632 15516 16688
rect 15377 16630 15516 16632
rect 15377 16627 15443 16630
rect 15510 16628 15516 16630
rect 15580 16628 15586 16692
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 3601 16282 3667 16285
rect 8385 16282 8451 16285
rect 3601 16280 8451 16282
rect 3601 16224 3606 16280
rect 3662 16224 8390 16280
rect 8446 16224 8451 16280
rect 3601 16222 8451 16224
rect 3601 16219 3667 16222
rect 8385 16219 8451 16222
rect 9438 16084 9444 16148
rect 9508 16146 9514 16148
rect 11421 16146 11487 16149
rect 9508 16144 11487 16146
rect 9508 16088 11426 16144
rect 11482 16088 11487 16144
rect 9508 16086 11487 16088
rect 9508 16084 9514 16086
rect 11421 16083 11487 16086
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 8569 15330 8635 15333
rect 8702 15330 8708 15332
rect 8569 15328 8708 15330
rect 8569 15272 8574 15328
rect 8630 15272 8708 15328
rect 8569 15270 8708 15272
rect 8569 15267 8635 15270
rect 8702 15268 8708 15270
rect 8772 15268 8778 15332
rect 8886 15268 8892 15332
rect 8956 15330 8962 15332
rect 10133 15330 10199 15333
rect 8956 15328 10199 15330
rect 8956 15272 10138 15328
rect 10194 15272 10199 15328
rect 8956 15270 10199 15272
rect 8956 15268 8962 15270
rect 10133 15267 10199 15270
rect 11697 15330 11763 15333
rect 11830 15330 11836 15332
rect 11697 15328 11836 15330
rect 11697 15272 11702 15328
rect 11758 15272 11836 15328
rect 11697 15270 11836 15272
rect 11697 15267 11763 15270
rect 11830 15268 11836 15270
rect 11900 15268 11906 15332
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 11237 15194 11303 15197
rect 14273 15194 14339 15197
rect 11237 15192 14339 15194
rect 11237 15136 11242 15192
rect 11298 15136 14278 15192
rect 14334 15136 14339 15192
rect 11237 15134 14339 15136
rect 11237 15131 11303 15134
rect 14273 15131 14339 15134
rect 3785 15058 3851 15061
rect 18965 15058 19031 15061
rect 3785 15056 19031 15058
rect 3785 15000 3790 15056
rect 3846 15000 18970 15056
rect 19026 15000 19031 15056
rect 3785 14998 19031 15000
rect 3785 14995 3851 14998
rect 18965 14995 19031 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 6678 14650 6684 14652
rect 4662 14590 6684 14650
rect 4521 14514 4587 14517
rect 4662 14514 4722 14590
rect 6678 14588 6684 14590
rect 6748 14650 6754 14652
rect 15561 14650 15627 14653
rect 17401 14650 17467 14653
rect 6748 14590 12450 14650
rect 6748 14588 6754 14590
rect 4521 14512 4722 14514
rect 4521 14456 4526 14512
rect 4582 14456 4722 14512
rect 4521 14454 4722 14456
rect 4521 14451 4587 14454
rect 6126 14452 6132 14516
rect 6196 14514 6202 14516
rect 9305 14514 9371 14517
rect 6196 14512 9371 14514
rect 6196 14456 9310 14512
rect 9366 14456 9371 14512
rect 6196 14454 9371 14456
rect 12390 14514 12450 14590
rect 15561 14648 17467 14650
rect 15561 14592 15566 14648
rect 15622 14592 17406 14648
rect 17462 14592 17467 14648
rect 15561 14590 17467 14592
rect 15561 14587 15627 14590
rect 17401 14587 17467 14590
rect 24577 14514 24643 14517
rect 12390 14512 24643 14514
rect 12390 14456 24582 14512
rect 24638 14456 24643 14512
rect 12390 14454 24643 14456
rect 6196 14452 6202 14454
rect 9305 14451 9371 14454
rect 24577 14451 24643 14454
rect 200 14378 800 14408
rect 3233 14378 3299 14381
rect 200 14376 3299 14378
rect 200 14320 3238 14376
rect 3294 14320 3299 14376
rect 200 14318 3299 14320
rect 200 14288 800 14318
rect 3233 14315 3299 14318
rect 8017 14378 8083 14381
rect 10593 14378 10659 14381
rect 8017 14376 10659 14378
rect 8017 14320 8022 14376
rect 8078 14320 10598 14376
rect 10654 14320 10659 14376
rect 8017 14318 10659 14320
rect 8017 14315 8083 14318
rect 10593 14315 10659 14318
rect 38285 14378 38351 14381
rect 39200 14378 39800 14408
rect 38285 14376 39800 14378
rect 38285 14320 38290 14376
rect 38346 14320 39800 14376
rect 38285 14318 39800 14320
rect 38285 14315 38351 14318
rect 39200 14288 39800 14318
rect 7189 14242 7255 14245
rect 10777 14242 10843 14245
rect 7189 14240 10843 14242
rect 7189 14184 7194 14240
rect 7250 14184 10782 14240
rect 10838 14184 10843 14240
rect 7189 14182 10843 14184
rect 7189 14179 7255 14182
rect 10777 14179 10843 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 5022 13908 5028 13972
rect 5092 13970 5098 13972
rect 9673 13970 9739 13973
rect 5092 13968 9739 13970
rect 5092 13912 9678 13968
rect 9734 13912 9739 13968
rect 5092 13910 9739 13912
rect 5092 13908 5098 13910
rect 9673 13907 9739 13910
rect 2957 13836 3023 13837
rect 5441 13836 5507 13837
rect 7833 13836 7899 13837
rect 2957 13832 3004 13836
rect 3068 13834 3074 13836
rect 5390 13834 5396 13836
rect 2957 13776 2962 13832
rect 2957 13772 3004 13776
rect 3068 13774 3114 13834
rect 5350 13774 5396 13834
rect 5460 13832 5507 13836
rect 7782 13834 7788 13836
rect 5502 13776 5507 13832
rect 3068 13772 3074 13774
rect 5390 13772 5396 13774
rect 5460 13772 5507 13776
rect 7742 13774 7788 13834
rect 7852 13832 7899 13836
rect 7894 13776 7899 13832
rect 7782 13772 7788 13774
rect 7852 13772 7899 13776
rect 2957 13771 3023 13772
rect 5441 13771 5507 13772
rect 7833 13771 7899 13772
rect 10225 13834 10291 13837
rect 10358 13834 10364 13836
rect 10225 13832 10364 13834
rect 10225 13776 10230 13832
rect 10286 13776 10364 13832
rect 10225 13774 10364 13776
rect 10225 13771 10291 13774
rect 10358 13772 10364 13774
rect 10428 13772 10434 13836
rect 12065 13834 12131 13837
rect 12566 13834 12572 13836
rect 12065 13832 12572 13834
rect 12065 13776 12070 13832
rect 12126 13776 12572 13832
rect 12065 13774 12572 13776
rect 12065 13771 12131 13774
rect 12566 13772 12572 13774
rect 12636 13772 12642 13836
rect 6637 13698 6703 13701
rect 8937 13698 9003 13701
rect 6637 13696 9003 13698
rect 6637 13640 6642 13696
rect 6698 13640 8942 13696
rect 8998 13640 9003 13696
rect 6637 13638 9003 13640
rect 6637 13635 6703 13638
rect 8937 13635 9003 13638
rect 12065 13698 12131 13701
rect 12341 13698 12407 13701
rect 12065 13696 12407 13698
rect 12065 13640 12070 13696
rect 12126 13640 12346 13696
rect 12402 13640 12407 13696
rect 12065 13638 12407 13640
rect 12065 13635 12131 13638
rect 12341 13635 12407 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 10317 13562 10383 13565
rect 15469 13562 15535 13565
rect 18137 13562 18203 13565
rect 10317 13560 18203 13562
rect 10317 13504 10322 13560
rect 10378 13504 15474 13560
rect 15530 13504 18142 13560
rect 18198 13504 18203 13560
rect 10317 13502 18203 13504
rect 10317 13499 10383 13502
rect 15469 13499 15535 13502
rect 18137 13499 18203 13502
rect 1853 13426 1919 13429
rect 5206 13426 5212 13428
rect 1853 13424 5212 13426
rect 1853 13368 1858 13424
rect 1914 13368 5212 13424
rect 1853 13366 5212 13368
rect 1853 13363 1919 13366
rect 5206 13364 5212 13366
rect 5276 13364 5282 13428
rect 4705 13156 4771 13157
rect 4654 13154 4660 13156
rect 4614 13094 4660 13154
rect 4724 13152 4771 13156
rect 4766 13096 4771 13152
rect 4654 13092 4660 13094
rect 4724 13092 4771 13096
rect 4705 13091 4771 13092
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 3417 13018 3483 13021
rect 8385 13018 8451 13021
rect 3417 13016 8451 13018
rect 3417 12960 3422 13016
rect 3478 12960 8390 13016
rect 8446 12960 8451 13016
rect 3417 12958 8451 12960
rect 3417 12955 3483 12958
rect 8385 12955 8451 12958
rect 10041 13018 10107 13021
rect 18505 13018 18571 13021
rect 10041 13016 18571 13018
rect 10041 12960 10046 13016
rect 10102 12960 18510 13016
rect 18566 12960 18571 13016
rect 10041 12958 18571 12960
rect 10041 12955 10107 12958
rect 18505 12955 18571 12958
rect 4337 12882 4403 12885
rect 9489 12882 9555 12885
rect 4337 12880 9555 12882
rect 4337 12824 4342 12880
rect 4398 12824 9494 12880
rect 9550 12824 9555 12880
rect 4337 12822 9555 12824
rect 4337 12819 4403 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 3785 12338 3851 12341
rect 4429 12338 4495 12341
rect 4616 12338 4676 12822
rect 9489 12819 9555 12822
rect 13629 12882 13695 12885
rect 14181 12882 14247 12885
rect 13629 12880 14247 12882
rect 13629 12824 13634 12880
rect 13690 12824 14186 12880
rect 14242 12824 14247 12880
rect 13629 12822 14247 12824
rect 13629 12819 13695 12822
rect 14181 12819 14247 12822
rect 5165 12746 5231 12749
rect 5441 12746 5507 12749
rect 5165 12744 5507 12746
rect 5165 12688 5170 12744
rect 5226 12688 5446 12744
rect 5502 12688 5507 12744
rect 5165 12686 5507 12688
rect 5165 12683 5231 12686
rect 5441 12683 5507 12686
rect 5257 12612 5323 12613
rect 5206 12610 5212 12612
rect 5166 12550 5212 12610
rect 5276 12608 5323 12612
rect 5318 12552 5323 12608
rect 5206 12548 5212 12550
rect 5276 12548 5323 12552
rect 5257 12547 5323 12548
rect 12617 12608 12683 12613
rect 12617 12552 12622 12608
rect 12678 12552 12683 12608
rect 12617 12547 12683 12552
rect 12620 12341 12680 12547
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 3785 12336 3986 12338
rect 3785 12280 3790 12336
rect 3846 12280 3986 12336
rect 3785 12278 3986 12280
rect 3785 12275 3851 12278
rect 3926 12205 3986 12278
rect 4429 12336 4676 12338
rect 4429 12280 4434 12336
rect 4490 12280 4676 12336
rect 4429 12278 4676 12280
rect 4429 12275 4495 12278
rect 7966 12276 7972 12340
rect 8036 12338 8042 12340
rect 8109 12338 8175 12341
rect 8036 12336 8175 12338
rect 8036 12280 8114 12336
rect 8170 12280 8175 12336
rect 8036 12278 8175 12280
rect 8036 12276 8042 12278
rect 8109 12275 8175 12278
rect 12617 12336 12683 12341
rect 12617 12280 12622 12336
rect 12678 12280 12683 12336
rect 12617 12275 12683 12280
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 3926 12200 4035 12205
rect 3926 12144 3974 12200
rect 4030 12144 4035 12200
rect 3926 12142 4035 12144
rect 3969 12139 4035 12142
rect 10041 12202 10107 12205
rect 12525 12202 12591 12205
rect 10041 12200 12591 12202
rect 10041 12144 10046 12200
rect 10102 12144 12530 12200
rect 12586 12144 12591 12200
rect 10041 12142 12591 12144
rect 10041 12139 10107 12142
rect 12525 12139 12591 12142
rect 4613 12066 4679 12069
rect 9121 12066 9187 12069
rect 4613 12064 9187 12066
rect 4613 12008 4618 12064
rect 4674 12008 9126 12064
rect 9182 12008 9187 12064
rect 4613 12006 9187 12008
rect 4613 12003 4679 12006
rect 9121 12003 9187 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 3693 11930 3759 11933
rect 4521 11930 4587 11933
rect 3693 11928 4587 11930
rect 3693 11872 3698 11928
rect 3754 11872 4526 11928
rect 4582 11872 4587 11928
rect 3693 11870 4587 11872
rect 3693 11867 3759 11870
rect 4521 11867 4587 11870
rect 7005 11930 7071 11933
rect 10593 11930 10659 11933
rect 7005 11928 10659 11930
rect 7005 11872 7010 11928
rect 7066 11872 10598 11928
rect 10654 11872 10659 11928
rect 7005 11870 10659 11872
rect 7005 11867 7071 11870
rect 10593 11867 10659 11870
rect 2773 11794 2839 11797
rect 4613 11794 4679 11797
rect 8569 11794 8635 11797
rect 2773 11792 8635 11794
rect 2773 11736 2778 11792
rect 2834 11736 4618 11792
rect 4674 11736 8574 11792
rect 8630 11736 8635 11792
rect 2773 11734 8635 11736
rect 2773 11731 2839 11734
rect 4613 11731 4679 11734
rect 8569 11731 8635 11734
rect 12893 11794 12959 11797
rect 18505 11794 18571 11797
rect 12893 11792 18571 11794
rect 12893 11736 12898 11792
rect 12954 11736 18510 11792
rect 18566 11736 18571 11792
rect 12893 11734 18571 11736
rect 12893 11731 12959 11734
rect 18505 11731 18571 11734
rect 5165 11658 5231 11661
rect 7649 11658 7715 11661
rect 5165 11656 7715 11658
rect 5165 11600 5170 11656
rect 5226 11600 7654 11656
rect 7710 11600 7715 11656
rect 5165 11598 7715 11600
rect 5165 11595 5231 11598
rect 7649 11595 7715 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 2773 11250 2839 11253
rect 9857 11250 9923 11253
rect 2773 11248 9923 11250
rect 2773 11192 2778 11248
rect 2834 11192 9862 11248
rect 9918 11192 9923 11248
rect 2773 11190 9923 11192
rect 2773 11187 2839 11190
rect 9857 11187 9923 11190
rect 200 10978 800 11008
rect 1669 10978 1735 10981
rect 200 10976 1735 10978
rect 200 10920 1674 10976
rect 1730 10920 1735 10976
rect 200 10918 1735 10920
rect 200 10888 800 10918
rect 1669 10915 1735 10918
rect 4153 10978 4219 10981
rect 5206 10978 5212 10980
rect 4153 10976 5212 10978
rect 4153 10920 4158 10976
rect 4214 10920 5212 10976
rect 4153 10918 5212 10920
rect 4153 10915 4219 10918
rect 5206 10916 5212 10918
rect 5276 10916 5282 10980
rect 38285 10978 38351 10981
rect 39200 10978 39800 11008
rect 38285 10976 39800 10978
rect 38285 10920 38290 10976
rect 38346 10920 39800 10976
rect 38285 10918 39800 10920
rect 38285 10915 38351 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 1945 10842 2011 10845
rect 5574 10842 5580 10844
rect 1945 10840 5580 10842
rect 1945 10784 1950 10840
rect 2006 10784 5580 10840
rect 1945 10782 5580 10784
rect 1945 10779 2011 10782
rect 5574 10780 5580 10782
rect 5644 10780 5650 10844
rect 3693 10570 3759 10573
rect 7598 10570 7604 10572
rect 3693 10568 7604 10570
rect 3693 10512 3698 10568
rect 3754 10512 7604 10568
rect 3693 10510 7604 10512
rect 3693 10507 3759 10510
rect 7598 10508 7604 10510
rect 7668 10508 7674 10572
rect 12566 10508 12572 10572
rect 12636 10570 12642 10572
rect 13077 10570 13143 10573
rect 12636 10568 13143 10570
rect 12636 10512 13082 10568
rect 13138 10512 13143 10568
rect 12636 10510 13143 10512
rect 12636 10508 12642 10510
rect 13077 10507 13143 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 2129 10162 2195 10165
rect 7097 10162 7163 10165
rect 2129 10160 7163 10162
rect 2129 10104 2134 10160
rect 2190 10104 7102 10160
rect 7158 10104 7163 10160
rect 2129 10102 7163 10104
rect 2129 10099 2195 10102
rect 7097 10099 7163 10102
rect 9121 10162 9187 10165
rect 9673 10162 9739 10165
rect 11973 10162 12039 10165
rect 9121 10160 12039 10162
rect 9121 10104 9126 10160
rect 9182 10104 9678 10160
rect 9734 10104 11978 10160
rect 12034 10104 12039 10160
rect 9121 10102 12039 10104
rect 9121 10099 9187 10102
rect 9673 10099 9739 10102
rect 11973 10099 12039 10102
rect 6269 9890 6335 9893
rect 9581 9890 9647 9893
rect 6269 9888 9647 9890
rect 6269 9832 6274 9888
rect 6330 9832 9586 9888
rect 9642 9832 9647 9888
rect 6269 9830 9647 9832
rect 6269 9827 6335 9830
rect 9581 9827 9647 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 200 9618 800 9648
rect 200 9558 1594 9618
rect 200 9528 800 9558
rect 1534 9482 1594 9558
rect 2773 9482 2839 9485
rect 1534 9480 2839 9482
rect 1534 9424 2778 9480
rect 2834 9424 2839 9480
rect 1534 9422 2839 9424
rect 2773 9419 2839 9422
rect 3049 9482 3115 9485
rect 4521 9482 4587 9485
rect 3049 9480 4587 9482
rect 3049 9424 3054 9480
rect 3110 9424 4526 9480
rect 4582 9424 4587 9480
rect 3049 9422 4587 9424
rect 3049 9419 3115 9422
rect 4521 9419 4587 9422
rect 6545 9346 6611 9349
rect 8937 9346 9003 9349
rect 6545 9344 9003 9346
rect 6545 9288 6550 9344
rect 6606 9288 8942 9344
rect 8998 9288 9003 9344
rect 6545 9286 9003 9288
rect 6545 9283 6611 9286
rect 8937 9283 9003 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4981 9210 5047 9213
rect 4846 9208 5047 9210
rect 4846 9152 4986 9208
rect 5042 9152 5047 9208
rect 4846 9150 5047 9152
rect 1669 8666 1735 8669
rect 2814 8666 2820 8668
rect 1669 8664 2820 8666
rect 1669 8608 1674 8664
rect 1730 8608 2820 8664
rect 1669 8606 2820 8608
rect 1669 8603 1735 8606
rect 2814 8604 2820 8606
rect 2884 8604 2890 8668
rect 4846 8533 4906 9150
rect 4981 9147 5047 9150
rect 6821 8938 6887 8941
rect 8293 8938 8359 8941
rect 6821 8936 8359 8938
rect 6821 8880 6826 8936
rect 6882 8880 8298 8936
rect 8354 8880 8359 8936
rect 6821 8878 8359 8880
rect 6821 8875 6887 8878
rect 8293 8875 8359 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 5073 8666 5139 8669
rect 9438 8666 9444 8668
rect 5073 8664 9444 8666
rect 5073 8608 5078 8664
rect 5134 8608 9444 8664
rect 5073 8606 9444 8608
rect 5073 8603 5139 8606
rect 9438 8604 9444 8606
rect 9508 8604 9514 8668
rect 4846 8528 4955 8533
rect 4846 8472 4894 8528
rect 4950 8472 4955 8528
rect 4846 8470 4955 8472
rect 4889 8467 4955 8470
rect 1945 8258 2011 8261
rect 2078 8258 2084 8260
rect 1945 8256 2084 8258
rect 1945 8200 1950 8256
rect 2006 8200 2084 8256
rect 1945 8198 2084 8200
rect 1945 8195 2011 8198
rect 2078 8196 2084 8198
rect 2148 8196 2154 8260
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 6678 8060 6684 8124
rect 6748 8122 6754 8124
rect 7925 8122 7991 8125
rect 6748 8120 7991 8122
rect 6748 8064 7930 8120
rect 7986 8064 7991 8120
rect 6748 8062 7991 8064
rect 6748 8060 6754 8062
rect 7925 8059 7991 8062
rect 3325 7986 3391 7989
rect 4654 7986 4660 7988
rect 3325 7984 4660 7986
rect 3325 7928 3330 7984
rect 3386 7928 4660 7984
rect 3325 7926 4660 7928
rect 3325 7923 3391 7926
rect 4654 7924 4660 7926
rect 4724 7924 4730 7988
rect 15510 7788 15516 7852
rect 15580 7850 15586 7852
rect 25405 7850 25471 7853
rect 15580 7848 25471 7850
rect 15580 7792 25410 7848
rect 25466 7792 25471 7848
rect 15580 7790 25471 7792
rect 15580 7788 15586 7790
rect 25405 7787 25471 7790
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4613 7578 4679 7581
rect 200 7576 4679 7578
rect 200 7520 4618 7576
rect 4674 7520 4679 7576
rect 200 7518 4679 7520
rect 200 7488 800 7518
rect 4613 7515 4679 7518
rect 4797 7578 4863 7581
rect 11278 7578 11284 7580
rect 4797 7576 11284 7578
rect 4797 7520 4802 7576
rect 4858 7520 11284 7576
rect 4797 7518 11284 7520
rect 4797 7515 4863 7518
rect 11278 7516 11284 7518
rect 11348 7516 11354 7580
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 4981 7442 5047 7445
rect 10726 7442 10732 7444
rect 4981 7440 10732 7442
rect 4981 7384 4986 7440
rect 5042 7384 10732 7440
rect 4981 7382 10732 7384
rect 4981 7379 5047 7382
rect 10726 7380 10732 7382
rect 10796 7380 10802 7444
rect 11462 7170 11468 7172
rect 4846 7110 11468 7170
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4846 7034 4906 7110
rect 11462 7108 11468 7110
rect 11532 7108 11538 7172
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4662 6974 4906 7034
rect 5441 7034 5507 7037
rect 8886 7034 8892 7036
rect 5441 7032 8892 7034
rect 5441 6976 5446 7032
rect 5502 6976 8892 7032
rect 5441 6974 8892 6976
rect 4153 6898 4219 6901
rect 4662 6898 4722 6974
rect 5441 6971 5507 6974
rect 8886 6972 8892 6974
rect 8956 6972 8962 7036
rect 4153 6896 4722 6898
rect 4153 6840 4158 6896
rect 4214 6840 4722 6896
rect 4153 6838 4722 6840
rect 5993 6898 6059 6901
rect 6126 6898 6132 6900
rect 5993 6896 6132 6898
rect 5993 6840 5998 6896
rect 6054 6840 6132 6896
rect 5993 6838 6132 6840
rect 4153 6835 4219 6838
rect 5993 6835 6059 6838
rect 6126 6836 6132 6838
rect 6196 6836 6202 6900
rect 7925 6898 7991 6901
rect 11830 6898 11836 6900
rect 7925 6896 11836 6898
rect 7925 6840 7930 6896
rect 7986 6840 11836 6896
rect 7925 6838 11836 6840
rect 7925 6835 7991 6838
rect 11830 6836 11836 6838
rect 11900 6836 11906 6900
rect 4797 6762 4863 6765
rect 10542 6762 10548 6764
rect 4797 6760 10548 6762
rect 4797 6704 4802 6760
rect 4858 6704 10548 6760
rect 4797 6702 10548 6704
rect 4797 6699 4863 6702
rect 10542 6700 10548 6702
rect 10612 6700 10618 6764
rect 3141 6626 3207 6629
rect 8702 6626 8708 6628
rect 3141 6624 8708 6626
rect 3141 6568 3146 6624
rect 3202 6568 8708 6624
rect 3141 6566 8708 6568
rect 3141 6563 3207 6566
rect 8702 6564 8708 6566
rect 8772 6564 8778 6628
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 5349 6490 5415 6493
rect 10358 6490 10364 6492
rect 5349 6488 10364 6490
rect 5349 6432 5354 6488
rect 5410 6432 10364 6488
rect 5349 6430 10364 6432
rect 5349 6427 5415 6430
rect 10358 6428 10364 6430
rect 10428 6428 10434 6492
rect 3233 6354 3299 6357
rect 10910 6354 10916 6356
rect 3233 6352 10916 6354
rect 3233 6296 3238 6352
rect 3294 6296 10916 6352
rect 3233 6294 10916 6296
rect 3233 6291 3299 6294
rect 10910 6292 10916 6294
rect 10980 6292 10986 6356
rect 200 6218 800 6248
rect 3785 6218 3851 6221
rect 200 6216 3851 6218
rect 200 6160 3790 6216
rect 3846 6160 3851 6216
rect 200 6158 3851 6160
rect 200 6128 800 6158
rect 3785 6155 3851 6158
rect 38285 6218 38351 6221
rect 39200 6218 39800 6248
rect 38285 6216 39800 6218
rect 38285 6160 38290 6216
rect 38346 6160 39800 6216
rect 38285 6158 39800 6160
rect 38285 6155 38351 6158
rect 39200 6128 39800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 5349 5948 5415 5949
rect 5349 5946 5396 5948
rect 5304 5944 5396 5946
rect 5304 5888 5354 5944
rect 5304 5886 5396 5888
rect 5349 5884 5396 5886
rect 5460 5884 5466 5948
rect 5349 5883 5415 5884
rect 2998 5612 3004 5676
rect 3068 5674 3074 5676
rect 4981 5674 5047 5677
rect 3068 5672 5047 5674
rect 3068 5616 4986 5672
rect 5042 5616 5047 5672
rect 3068 5614 5047 5616
rect 3068 5612 3074 5614
rect 4981 5611 5047 5614
rect 3693 5538 3759 5541
rect 7782 5538 7788 5540
rect 3693 5536 7788 5538
rect 3693 5480 3698 5536
rect 3754 5480 7788 5536
rect 3693 5478 7788 5480
rect 3693 5475 3759 5478
rect 7782 5476 7788 5478
rect 7852 5476 7858 5540
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4337 5402 4403 5405
rect 5022 5402 5028 5404
rect 4337 5400 5028 5402
rect 4337 5344 4342 5400
rect 4398 5344 5028 5400
rect 4337 5342 5028 5344
rect 4337 5339 4403 5342
rect 5022 5340 5028 5342
rect 5092 5340 5098 5404
rect 4210 4928 4526 4929
rect 200 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1761 4858 1827 4861
rect 200 4856 1827 4858
rect 200 4800 1766 4856
rect 1822 4800 1827 4856
rect 200 4798 1827 4800
rect 200 4768 800 4798
rect 1761 4795 1827 4798
rect 4245 4722 4311 4725
rect 11094 4722 11100 4724
rect 4245 4720 11100 4722
rect 4245 4664 4250 4720
rect 4306 4664 11100 4720
rect 4245 4662 11100 4664
rect 4245 4659 4311 4662
rect 11094 4660 11100 4662
rect 11164 4660 11170 4724
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38193 4178 38259 4181
rect 39200 4178 39800 4208
rect 38193 4176 39800 4178
rect 38193 4120 38198 4176
rect 38254 4120 39800 4176
rect 38193 4118 39800 4120
rect 38193 4115 38259 4118
rect 39200 4088 39800 4118
rect 4521 4042 4587 4045
rect 4838 4042 4844 4044
rect 4521 4040 4844 4042
rect 4521 3984 4526 4040
rect 4582 3984 4844 4040
rect 4521 3982 4844 3984
rect 4521 3979 4587 3982
rect 4838 3980 4844 3982
rect 4908 3980 4914 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 200 2818 800 2848
rect 3969 2818 4035 2821
rect 200 2816 4035 2818
rect 200 2760 3974 2816
rect 4030 2760 4035 2816
rect 200 2758 4035 2760
rect 200 2728 800 2758
rect 3969 2755 4035 2758
rect 38285 2818 38351 2821
rect 39200 2818 39800 2848
rect 38285 2816 39800 2818
rect 38285 2760 38290 2816
rect 38346 2760 39800 2816
rect 38285 2758 39800 2760
rect 38285 2755 38351 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 200 1458 800 1488
rect 4061 1458 4127 1461
rect 200 1456 4127 1458
rect 200 1400 4066 1456
rect 4122 1400 4127 1456
rect 200 1398 4127 1400
rect 200 1368 800 1398
rect 4061 1395 4127 1398
rect 38193 1458 38259 1461
rect 39200 1458 39800 1488
rect 38193 1456 39800 1458
rect 38193 1400 38198 1456
rect 38254 1400 39800 1456
rect 38193 1398 39800 1400
rect 38193 1395 38259 1398
rect 39200 1368 39800 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 5764 31784 5828 31788
rect 5764 31728 5778 31784
rect 5778 31728 5828 31784
rect 5764 31724 5828 31728
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 7972 23020 8036 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 5212 22068 5276 22132
rect 2820 21796 2884 21860
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 5580 20768 5644 20772
rect 5580 20712 5630 20768
rect 5630 20712 5644 20768
rect 5580 20708 5644 20712
rect 7604 20768 7668 20772
rect 7604 20712 7618 20768
rect 7618 20712 7668 20768
rect 7604 20708 7668 20712
rect 11100 20768 11164 20772
rect 11100 20712 11114 20768
rect 11114 20712 11164 20768
rect 11100 20708 11164 20712
rect 11284 20768 11348 20772
rect 11284 20712 11334 20768
rect 11334 20712 11348 20768
rect 11284 20708 11348 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 10916 19892 10980 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4844 19348 4908 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 10732 19408 10796 19412
rect 10732 19352 10782 19408
rect 10782 19352 10796 19408
rect 10732 19348 10796 19352
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 11468 17988 11532 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 5764 17852 5828 17916
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 2084 17036 2148 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 10548 16628 10612 16692
rect 15516 16628 15580 16692
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 9444 16084 9508 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 8708 15268 8772 15332
rect 8892 15268 8956 15332
rect 11836 15268 11900 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 6684 14588 6748 14652
rect 6132 14452 6196 14516
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 5028 13908 5092 13972
rect 3004 13832 3068 13836
rect 3004 13776 3018 13832
rect 3018 13776 3068 13832
rect 3004 13772 3068 13776
rect 5396 13832 5460 13836
rect 5396 13776 5446 13832
rect 5446 13776 5460 13832
rect 5396 13772 5460 13776
rect 7788 13832 7852 13836
rect 7788 13776 7838 13832
rect 7838 13776 7852 13832
rect 7788 13772 7852 13776
rect 10364 13772 10428 13836
rect 12572 13772 12636 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 5212 13364 5276 13428
rect 4660 13152 4724 13156
rect 4660 13096 4710 13152
rect 4710 13096 4724 13152
rect 4660 13092 4724 13096
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 5212 12608 5276 12612
rect 5212 12552 5262 12608
rect 5262 12552 5276 12608
rect 5212 12548 5276 12552
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 7972 12276 8036 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 5212 10916 5276 10980
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 5580 10780 5644 10844
rect 7604 10508 7668 10572
rect 12572 10508 12636 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 2820 8604 2884 8668
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 9444 8604 9508 8668
rect 2084 8196 2148 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 6684 8060 6748 8124
rect 4660 7924 4724 7988
rect 15516 7788 15580 7852
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 11284 7516 11348 7580
rect 10732 7380 10796 7444
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 11468 7108 11532 7172
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 8892 6972 8956 7036
rect 6132 6836 6196 6900
rect 11836 6836 11900 6900
rect 10548 6700 10612 6764
rect 8708 6564 8772 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 10364 6428 10428 6492
rect 10916 6292 10980 6356
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 5396 5944 5460 5948
rect 5396 5888 5410 5944
rect 5410 5888 5460 5944
rect 5396 5884 5460 5888
rect 3004 5612 3068 5676
rect 7788 5476 7852 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 5028 5340 5092 5404
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 11100 4660 11164 4724
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4844 3980 4908 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 5763 31788 5829 31789
rect 5763 31724 5764 31788
rect 5828 31724 5829 31788
rect 5763 31723 5829 31724
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 2819 21860 2885 21861
rect 2819 21796 2820 21860
rect 2884 21796 2885 21860
rect 2819 21795 2885 21796
rect 2083 17100 2149 17101
rect 2083 17036 2084 17100
rect 2148 17036 2149 17100
rect 2083 17035 2149 17036
rect 2086 8261 2146 17035
rect 2822 8669 2882 21795
rect 4208 21248 4528 22272
rect 5211 22132 5277 22133
rect 5211 22068 5212 22132
rect 5276 22068 5277 22132
rect 5211 22067 5277 22068
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4843 19412 4909 19413
rect 4843 19348 4844 19412
rect 4908 19348 4909 19412
rect 4843 19347 4909 19348
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 3003 13836 3069 13837
rect 3003 13772 3004 13836
rect 3068 13772 3069 13836
rect 3003 13771 3069 13772
rect 2819 8668 2885 8669
rect 2819 8604 2820 8668
rect 2884 8604 2885 8668
rect 2819 8603 2885 8604
rect 2083 8260 2149 8261
rect 2083 8196 2084 8260
rect 2148 8196 2149 8260
rect 2083 8195 2149 8196
rect 3006 5677 3066 13771
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4659 13156 4725 13157
rect 4659 13092 4660 13156
rect 4724 13092 4725 13156
rect 4659 13091 4725 13092
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4662 7989 4722 13091
rect 4659 7988 4725 7989
rect 4659 7924 4660 7988
rect 4724 7924 4725 7988
rect 4659 7923 4725 7924
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 3003 5676 3069 5677
rect 3003 5612 3004 5676
rect 3068 5612 3069 5676
rect 3003 5611 3069 5612
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4846 4045 4906 19347
rect 5027 13972 5093 13973
rect 5027 13908 5028 13972
rect 5092 13908 5093 13972
rect 5027 13907 5093 13908
rect 5030 5405 5090 13907
rect 5214 13429 5274 22067
rect 5579 20772 5645 20773
rect 5579 20708 5580 20772
rect 5644 20708 5645 20772
rect 5579 20707 5645 20708
rect 5395 13836 5461 13837
rect 5395 13772 5396 13836
rect 5460 13772 5461 13836
rect 5395 13771 5461 13772
rect 5211 13428 5277 13429
rect 5211 13364 5212 13428
rect 5276 13364 5277 13428
rect 5211 13363 5277 13364
rect 5211 12612 5277 12613
rect 5211 12548 5212 12612
rect 5276 12548 5277 12612
rect 5211 12547 5277 12548
rect 5214 10981 5274 12547
rect 5211 10980 5277 10981
rect 5211 10916 5212 10980
rect 5276 10916 5277 10980
rect 5211 10915 5277 10916
rect 5398 5949 5458 13771
rect 5582 10845 5642 20707
rect 5766 17917 5826 31723
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 7971 23084 8037 23085
rect 7971 23020 7972 23084
rect 8036 23020 8037 23084
rect 7971 23019 8037 23020
rect 7603 20772 7669 20773
rect 7603 20708 7604 20772
rect 7668 20708 7669 20772
rect 7603 20707 7669 20708
rect 5763 17916 5829 17917
rect 5763 17852 5764 17916
rect 5828 17852 5829 17916
rect 5763 17851 5829 17852
rect 6683 14652 6749 14653
rect 6683 14588 6684 14652
rect 6748 14588 6749 14652
rect 6683 14587 6749 14588
rect 6131 14516 6197 14517
rect 6131 14452 6132 14516
rect 6196 14452 6197 14516
rect 6131 14451 6197 14452
rect 5579 10844 5645 10845
rect 5579 10780 5580 10844
rect 5644 10780 5645 10844
rect 5579 10779 5645 10780
rect 6134 6901 6194 14451
rect 6686 8125 6746 14587
rect 7606 10573 7666 20707
rect 7787 13836 7853 13837
rect 7787 13772 7788 13836
rect 7852 13772 7853 13836
rect 7787 13771 7853 13772
rect 7603 10572 7669 10573
rect 7603 10508 7604 10572
rect 7668 10508 7669 10572
rect 7603 10507 7669 10508
rect 6683 8124 6749 8125
rect 6683 8060 6684 8124
rect 6748 8060 6749 8124
rect 6683 8059 6749 8060
rect 6131 6900 6197 6901
rect 6131 6836 6132 6900
rect 6196 6836 6197 6900
rect 6131 6835 6197 6836
rect 5395 5948 5461 5949
rect 5395 5884 5396 5948
rect 5460 5884 5461 5948
rect 5395 5883 5461 5884
rect 7790 5541 7850 13771
rect 7974 12341 8034 23019
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 11099 20772 11165 20773
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 11283 20772 11349 20773
rect 11283 20708 11284 20772
rect 11348 20708 11349 20772
rect 11283 20707 11349 20708
rect 10915 19956 10981 19957
rect 10915 19892 10916 19956
rect 10980 19892 10981 19956
rect 10915 19891 10981 19892
rect 10731 19412 10797 19413
rect 10731 19348 10732 19412
rect 10796 19348 10797 19412
rect 10731 19347 10797 19348
rect 10547 16692 10613 16693
rect 10547 16628 10548 16692
rect 10612 16628 10613 16692
rect 10547 16627 10613 16628
rect 9443 16148 9509 16149
rect 9443 16084 9444 16148
rect 9508 16084 9509 16148
rect 9443 16083 9509 16084
rect 8707 15332 8773 15333
rect 8707 15268 8708 15332
rect 8772 15268 8773 15332
rect 8707 15267 8773 15268
rect 8891 15332 8957 15333
rect 8891 15268 8892 15332
rect 8956 15268 8957 15332
rect 8891 15267 8957 15268
rect 7971 12340 8037 12341
rect 7971 12276 7972 12340
rect 8036 12276 8037 12340
rect 7971 12275 8037 12276
rect 8710 6629 8770 15267
rect 8894 7037 8954 15267
rect 9446 8669 9506 16083
rect 10363 13836 10429 13837
rect 10363 13772 10364 13836
rect 10428 13772 10429 13836
rect 10363 13771 10429 13772
rect 9443 8668 9509 8669
rect 9443 8604 9444 8668
rect 9508 8604 9509 8668
rect 9443 8603 9509 8604
rect 8891 7036 8957 7037
rect 8891 6972 8892 7036
rect 8956 6972 8957 7036
rect 8891 6971 8957 6972
rect 8707 6628 8773 6629
rect 8707 6564 8708 6628
rect 8772 6564 8773 6628
rect 8707 6563 8773 6564
rect 10366 6493 10426 13771
rect 10550 6765 10610 16627
rect 10734 7445 10794 19347
rect 10731 7444 10797 7445
rect 10731 7380 10732 7444
rect 10796 7380 10797 7444
rect 10731 7379 10797 7380
rect 10547 6764 10613 6765
rect 10547 6700 10548 6764
rect 10612 6700 10613 6764
rect 10547 6699 10613 6700
rect 10363 6492 10429 6493
rect 10363 6428 10364 6492
rect 10428 6428 10429 6492
rect 10363 6427 10429 6428
rect 10918 6357 10978 19891
rect 10915 6356 10981 6357
rect 10915 6292 10916 6356
rect 10980 6292 10981 6356
rect 10915 6291 10981 6292
rect 7787 5540 7853 5541
rect 7787 5476 7788 5540
rect 7852 5476 7853 5540
rect 7787 5475 7853 5476
rect 5027 5404 5093 5405
rect 5027 5340 5028 5404
rect 5092 5340 5093 5404
rect 5027 5339 5093 5340
rect 11102 4725 11162 20707
rect 11286 7581 11346 20707
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 11467 18052 11533 18053
rect 11467 17988 11468 18052
rect 11532 17988 11533 18052
rect 11467 17987 11533 17988
rect 11283 7580 11349 7581
rect 11283 7516 11284 7580
rect 11348 7516 11349 7580
rect 11283 7515 11349 7516
rect 11470 7173 11530 17987
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 15515 16692 15581 16693
rect 15515 16628 15516 16692
rect 15580 16628 15581 16692
rect 15515 16627 15581 16628
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11467 7172 11533 7173
rect 11467 7108 11468 7172
rect 11532 7108 11533 7172
rect 11467 7107 11533 7108
rect 11838 6901 11898 15267
rect 12571 13836 12637 13837
rect 12571 13772 12572 13836
rect 12636 13772 12637 13836
rect 12571 13771 12637 13772
rect 12574 10573 12634 13771
rect 12571 10572 12637 10573
rect 12571 10508 12572 10572
rect 12636 10508 12637 10572
rect 12571 10507 12637 10508
rect 15518 7853 15578 16627
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 15515 7852 15581 7853
rect 15515 7788 15516 7852
rect 15580 7788 15581 7852
rect 15515 7787 15581 7788
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 11835 6900 11901 6901
rect 11835 6836 11836 6900
rect 11900 6836 11901 6900
rect 11835 6835 11901 6836
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 11099 4724 11165 4725
rect 11099 4660 11100 4724
rect 11164 4660 11165 4724
rect 11099 4659 11165 4660
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 4843 4044 4909 4045
rect 4843 3980 4844 4044
rect 4908 3980 4909 4044
rect 4843 3979 4909 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 3956 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21
timestamp 1667941163
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91
timestamp 1667941163
transform 1 0 9476 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1667941163
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1667941163
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1667941163
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_118
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 1667941163
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_182
timestamp 1667941163
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1667941163
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1667941163
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1667941163
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259
timestamp 1667941163
transform 1 0 24932 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_267
timestamp 1667941163
transform 1 0 25668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1667941163
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1667941163
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1667941163
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1667941163
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1667941163
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1667941163
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_370
timestamp 1667941163
transform 1 0 35144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_378
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1667941163
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1667941163
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_37
timestamp 1667941163
transform 1 0 4508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_62
timestamp 1667941163
transform 1 0 6808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_74
timestamp 1667941163
transform 1 0 7912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_86
timestamp 1667941163
transform 1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_98
timestamp 1667941163
transform 1 0 10120 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1667941163
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_289
timestamp 1667941163
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_295
timestamp 1667941163
transform 1 0 28244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_307
timestamp 1667941163
transform 1 0 29348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_319
timestamp 1667941163
transform 1 0 30452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1667941163
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1667941163
transform 1 0 2852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_34
timestamp 1667941163
transform 1 0 4232 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_42
timestamp 1667941163
transform 1 0 4968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1667941163
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_60
timestamp 1667941163
transform 1 0 6624 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_72
timestamp 1667941163
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1667941163
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1667941163
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_29
timestamp 1667941163
transform 1 0 3772 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1667941163
transform 1 0 4324 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1667941163
transform 1 0 5336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1667941163
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1667941163
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1667941163
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_19
timestamp 1667941163
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1667941163
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1667941163
transform 1 0 4784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1667941163
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1667941163
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_58
timestamp 1667941163
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1667941163
transform 1 0 9660 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_99
timestamp 1667941163
transform 1 0 10212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_111
timestamp 1667941163
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_123
timestamp 1667941163
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1667941163
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_276
timestamp 1667941163
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_288
timestamp 1667941163
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1667941163
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1667941163
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1667941163
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1667941163
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1667941163
transform 1 0 4508 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1667941163
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1667941163
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_76
timestamp 1667941163
transform 1 0 8096 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1667941163
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1667941163
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_356
timestamp 1667941163
transform 1 0 33856 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_368
timestamp 1667941163
transform 1 0 34960 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_380
timestamp 1667941163
transform 1 0 36064 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1667941163
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_16
timestamp 1667941163
transform 1 0 2576 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1667941163
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1667941163
transform 1 0 4232 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1667941163
transform 1 0 5520 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_55
timestamp 1667941163
transform 1 0 6164 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1667941163
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_69
timestamp 1667941163
transform 1 0 7452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1667941163
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_112
timestamp 1667941163
transform 1 0 11408 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_183
timestamp 1667941163
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190
timestamp 1667941163
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_215
timestamp 1667941163
transform 1 0 20884 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_219
timestamp 1667941163
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_231
timestamp 1667941163
transform 1 0 22356 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_239
timestamp 1667941163
transform 1 0 23092 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_8
timestamp 1667941163
transform 1 0 1840 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_17
timestamp 1667941163
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1667941163
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_31
timestamp 1667941163
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1667941163
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1667941163
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1667941163
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1667941163
transform 1 0 6808 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1667941163
transform 1 0 7544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1667941163
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_141
timestamp 1667941163
transform 1 0 14076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1667941163
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_190
timestamp 1667941163
transform 1 0 18584 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_202
timestamp 1667941163
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_214
timestamp 1667941163
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_230
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_242
timestamp 1667941163
transform 1 0 23368 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_254
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_266
timestamp 1667941163
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1667941163
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1667941163
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_345
timestamp 1667941163
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_401
timestamp 1667941163
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_8
timestamp 1667941163
transform 1 0 1840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_12
timestamp 1667941163
transform 1 0 2208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1667941163
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1667941163
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1667941163
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1667941163
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_55
timestamp 1667941163
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_62
timestamp 1667941163
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1667941163
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1667941163
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_90
timestamp 1667941163
transform 1 0 9384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_118
timestamp 1667941163
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_122
timestamp 1667941163
transform 1 0 12328 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_126
timestamp 1667941163
transform 1 0 12696 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_261
timestamp 1667941163
transform 1 0 25116 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_266
timestamp 1667941163
transform 1 0 25576 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_278
timestamp 1667941163
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_290
timestamp 1667941163
transform 1 0 27784 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_302
timestamp 1667941163
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1667941163
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_34
timestamp 1667941163
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1667941163
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1667941163
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1667941163
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1667941163
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1667941163
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_135
timestamp 1667941163
transform 1 0 13524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_147
timestamp 1667941163
transform 1 0 14628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_159
timestamp 1667941163
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_174
timestamp 1667941163
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_186
timestamp 1667941163
transform 1 0 18216 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_198
timestamp 1667941163
transform 1 0 19320 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_210
timestamp 1667941163
transform 1 0 20424 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_384
timestamp 1667941163
transform 1 0 36432 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1667941163
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_34
timestamp 1667941163
transform 1 0 4232 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_48
timestamp 1667941163
transform 1 0 5520 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_54
timestamp 1667941163
transform 1 0 6072 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1667941163
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_96
timestamp 1667941163
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1667941163
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1667941163
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_294
timestamp 1667941163
transform 1 0 28152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1667941163
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_8
timestamp 1667941163
transform 1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_33
timestamp 1667941163
transform 1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1667941163
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_47
timestamp 1667941163
transform 1 0 5428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1667941163
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1667941163
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_91
timestamp 1667941163
transform 1 0 9476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1667941163
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1667941163
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1667941163
transform 1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1667941163
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_143
timestamp 1667941163
transform 1 0 14260 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_150
timestamp 1667941163
transform 1 0 14904 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1667941163
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_210
timestamp 1667941163
transform 1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1667941163
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_360
timestamp 1667941163
transform 1 0 34224 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_372
timestamp 1667941163
transform 1 0 35328 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1667941163
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1667941163
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_96
timestamp 1667941163
transform 1 0 9936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1667941163
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1667941163
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1667941163
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_146
timestamp 1667941163
transform 1 0 14536 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1667941163
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_288
timestamp 1667941163
transform 1 0 27600 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1667941163
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_10
timestamp 1667941163
transform 1 0 2024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_17
timestamp 1667941163
transform 1 0 2668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_44
timestamp 1667941163
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_80
timestamp 1667941163
transform 1 0 8464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_89
timestamp 1667941163
transform 1 0 9292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_96
timestamp 1667941163
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1667941163
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_132
timestamp 1667941163
transform 1 0 13248 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1667941163
transform 1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1667941163
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_155
timestamp 1667941163
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_364
timestamp 1667941163
transform 1 0 34592 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_376
timestamp 1667941163
transform 1 0 35696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1667941163
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_12
timestamp 1667941163
transform 1 0 2208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_19
timestamp 1667941163
transform 1 0 2852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1667941163
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_58
timestamp 1667941163
transform 1 0 6440 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1667941163
transform 1 0 6992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1667941163
transform 1 0 7360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_75
timestamp 1667941163
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_108
timestamp 1667941163
transform 1 0 11040 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_112
timestamp 1667941163
transform 1 0 11408 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_116
timestamp 1667941163
transform 1 0 11776 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1667941163
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1667941163
transform 1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1667941163
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1667941163
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_160
timestamp 1667941163
transform 1 0 15824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1667941163
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1667941163
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_202
timestamp 1667941163
transform 1 0 19688 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_210
timestamp 1667941163
transform 1 0 20424 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_214
timestamp 1667941163
transform 1 0 20792 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_226
timestamp 1667941163
transform 1 0 21896 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_238
timestamp 1667941163
transform 1 0 23000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1667941163
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1667941163
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_314
timestamp 1667941163
transform 1 0 29992 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_326
timestamp 1667941163
transform 1 0 31096 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_338
timestamp 1667941163
transform 1 0 32200 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_350
timestamp 1667941163
transform 1 0 33304 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1667941163
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1667941163
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_16
timestamp 1667941163
transform 1 0 2576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_23
timestamp 1667941163
transform 1 0 3220 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_34
timestamp 1667941163
transform 1 0 4232 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_42
timestamp 1667941163
transform 1 0 4968 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_47
timestamp 1667941163
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1667941163
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_65
timestamp 1667941163
transform 1 0 7084 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_72
timestamp 1667941163
transform 1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1667941163
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1667941163
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1667941163
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1667941163
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1667941163
transform 1 0 13340 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1667941163
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_150
timestamp 1667941163
transform 1 0 14904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1667941163
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_174
timestamp 1667941163
transform 1 0 17112 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_180
timestamp 1667941163
transform 1 0 17664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1667941163
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1667941163
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_203
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_215
timestamp 1667941163
transform 1 0 20884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1667941163
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_233
timestamp 1667941163
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_238
timestamp 1667941163
transform 1 0 23000 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_250
timestamp 1667941163
transform 1 0 24104 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_262
timestamp 1667941163
transform 1 0 25208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1667941163
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_301
timestamp 1667941163
transform 1 0 28796 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_313
timestamp 1667941163
transform 1 0 29900 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1667941163
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1667941163
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_358
timestamp 1667941163
transform 1 0 34040 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_370
timestamp 1667941163
transform 1 0 35144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_382
timestamp 1667941163
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1667941163
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_33
timestamp 1667941163
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_37
timestamp 1667941163
transform 1 0 4508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1667941163
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1667941163
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1667941163
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_116
timestamp 1667941163
transform 1 0 11776 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1667941163
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 1667941163
transform 1 0 12972 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1667941163
transform 1 0 14536 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1667941163
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_162
timestamp 1667941163
transform 1 0 16008 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1667941163
transform 1 0 17112 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_181
timestamp 1667941163
transform 1 0 17756 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 1667941163
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1667941163
transform 1 0 20240 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1667941163
transform 1 0 22080 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_235
timestamp 1667941163
transform 1 0 22724 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1667941163
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_405
timestamp 1667941163
transform 1 0 38364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_12
timestamp 1667941163
transform 1 0 2208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 1667941163
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_47
timestamp 1667941163
transform 1 0 5428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1667941163
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_92
timestamp 1667941163
transform 1 0 9568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1667941163
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1667941163
transform 1 0 12420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 1667941163
transform 1 0 13156 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_135
timestamp 1667941163
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_142
timestamp 1667941163
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_156
timestamp 1667941163
transform 1 0 15456 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_162
timestamp 1667941163
transform 1 0 16008 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1667941163
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1667941163
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1667941163
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_204
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_213
timestamp 1667941163
transform 1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1667941163
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1667941163
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1667941163
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_34
timestamp 1667941163
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_38
timestamp 1667941163
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_62
timestamp 1667941163
transform 1 0 6808 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_66
timestamp 1667941163
transform 1 0 7176 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1667941163
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1667941163
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1667941163
transform 1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1667941163
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1667941163
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1667941163
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_152
timestamp 1667941163
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1667941163
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1667941163
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_176
timestamp 1667941163
transform 1 0 17296 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1667941163
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1667941163
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_203
timestamp 1667941163
transform 1 0 19780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1667941163
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_223
timestamp 1667941163
transform 1 0 21620 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_239
timestamp 1667941163
transform 1 0 23092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1667941163
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1667941163
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1667941163
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_317
timestamp 1667941163
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_323
timestamp 1667941163
transform 1 0 30820 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_335
timestamp 1667941163
transform 1 0 31924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_347
timestamp 1667941163
transform 1 0 33028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1667941163
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_28
timestamp 1667941163
transform 1 0 3680 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1667941163
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_80
timestamp 1667941163
transform 1 0 8464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_94
timestamp 1667941163
transform 1 0 9752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1667941163
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1667941163
transform 1 0 11960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_131
timestamp 1667941163
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_144
timestamp 1667941163
transform 1 0 14352 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1667941163
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1667941163
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1667941163
transform 1 0 17204 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_183
timestamp 1667941163
transform 1 0 17940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_188
timestamp 1667941163
transform 1 0 18400 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_194
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1667941163
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_211
timestamp 1667941163
transform 1 0 20516 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1667941163
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_234
timestamp 1667941163
transform 1 0 22632 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1667941163
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1667941163
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1667941163
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1667941163
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1667941163
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1667941163
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1667941163
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1667941163
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1667941163
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_54
timestamp 1667941163
transform 1 0 6072 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_60
timestamp 1667941163
transform 1 0 6624 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_107
timestamp 1667941163
transform 1 0 10948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1667941163
transform 1 0 12052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1667941163
transform 1 0 13156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_151
timestamp 1667941163
transform 1 0 14996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_160
timestamp 1667941163
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1667941163
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_180
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1667941163
transform 1 0 20148 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1667941163
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_229
timestamp 1667941163
transform 1 0 22172 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1667941163
transform 1 0 22816 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1667941163
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_265
timestamp 1667941163
transform 1 0 25484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_272
timestamp 1667941163
transform 1 0 26128 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_279
timestamp 1667941163
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1667941163
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1667941163
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1667941163
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1667941163
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1667941163
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1667941163
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1667941163
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_19
timestamp 1667941163
transform 1 0 2852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_46
timestamp 1667941163
transform 1 0 5336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_50
timestamp 1667941163
transform 1 0 5704 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_71
timestamp 1667941163
transform 1 0 7636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1667941163
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1667941163
transform 1 0 12420 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1667941163
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1667941163
transform 1 0 14628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1667941163
transform 1 0 14996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1667941163
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1667941163
transform 1 0 18032 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1667941163
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_195
timestamp 1667941163
transform 1 0 19044 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_202
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1667941163
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_231
timestamp 1667941163
transform 1 0 22356 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_239
timestamp 1667941163
transform 1 0 23092 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_248
timestamp 1667941163
transform 1 0 23920 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_264
timestamp 1667941163
transform 1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_271
timestamp 1667941163
transform 1 0 26036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1667941163
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1667941163
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1667941163
transform 1 0 4416 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_58
timestamp 1667941163
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1667941163
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_120
timestamp 1667941163
transform 1 0 12144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_128
timestamp 1667941163
transform 1 0 12880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1667941163
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_151
timestamp 1667941163
transform 1 0 14996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_155
timestamp 1667941163
transform 1 0 15364 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_159
timestamp 1667941163
transform 1 0 15732 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1667941163
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_184
timestamp 1667941163
transform 1 0 18032 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_203
timestamp 1667941163
transform 1 0 19780 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1667941163
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_232
timestamp 1667941163
transform 1 0 22448 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1667941163
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_263
timestamp 1667941163
transform 1 0 25300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_275
timestamp 1667941163
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_282
timestamp 1667941163
transform 1 0 27048 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_294
timestamp 1667941163
transform 1 0 28152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_316
timestamp 1667941163
transform 1 0 30176 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_328
timestamp 1667941163
transform 1 0 31280 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_340
timestamp 1667941163
transform 1 0 32384 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_352
timestamp 1667941163
transform 1 0 33488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1667941163
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1667941163
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_401
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1667941163
transform 1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1667941163
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_83
timestamp 1667941163
transform 1 0 8740 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1667941163
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1667941163
transform 1 0 12420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1667941163
transform 1 0 13524 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_143
timestamp 1667941163
transform 1 0 14260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_148
timestamp 1667941163
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1667941163
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1667941163
transform 1 0 18032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_188
timestamp 1667941163
transform 1 0 18400 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_192
timestamp 1667941163
transform 1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1667941163
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1667941163
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1667941163
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_238
timestamp 1667941163
transform 1 0 23000 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1667941163
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_252
timestamp 1667941163
transform 1 0 24288 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_259
timestamp 1667941163
transform 1 0 24932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1667941163
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1667941163
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_355
timestamp 1667941163
transform 1 0 33764 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_363
timestamp 1667941163
transform 1 0 34500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_368
timestamp 1667941163
transform 1 0 34960 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_375
timestamp 1667941163
transform 1 0 35604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1667941163
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1667941163
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_14
timestamp 1667941163
transform 1 0 2392 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_37
timestamp 1667941163
transform 1 0 4508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_62
timestamp 1667941163
transform 1 0 6808 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1667941163
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1667941163
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_100
timestamp 1667941163
transform 1 0 10304 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_106
timestamp 1667941163
transform 1 0 10856 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1667941163
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_127
timestamp 1667941163
transform 1 0 12788 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1667941163
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1667941163
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1667941163
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_166
timestamp 1667941163
transform 1 0 16376 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_175
timestamp 1667941163
transform 1 0 17204 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1667941163
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_221
timestamp 1667941163
transform 1 0 21436 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_229
timestamp 1667941163
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1667941163
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1667941163
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_270
timestamp 1667941163
transform 1 0 25944 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_282
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_294
timestamp 1667941163
transform 1 0 28152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1667941163
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1667941163
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1667941163
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1667941163
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1667941163
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_28
timestamp 1667941163
transform 1 0 3680 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1667941163
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1667941163
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_86
timestamp 1667941163
transform 1 0 9016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1667941163
transform 1 0 12420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1667941163
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1667941163
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_148
timestamp 1667941163
transform 1 0 14720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1667941163
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_179
timestamp 1667941163
transform 1 0 17572 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1667941163
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1667941163
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1667941163
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1667941163
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_234
timestamp 1667941163
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_238
timestamp 1667941163
transform 1 0 23000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1667941163
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_257
timestamp 1667941163
transform 1 0 24748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1667941163
transform 1 0 25852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_277
timestamp 1667941163
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_314
timestamp 1667941163
transform 1 0 29992 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_326
timestamp 1667941163
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1667941163
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1667941163
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1667941163
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_51
timestamp 1667941163
transform 1 0 5796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_64
timestamp 1667941163
transform 1 0 6992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_68
timestamp 1667941163
transform 1 0 7360 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_78
timestamp 1667941163
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1667941163
transform 1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1667941163
transform 1 0 11316 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_115
timestamp 1667941163
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_127
timestamp 1667941163
transform 1 0 12788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1667941163
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 1667941163
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_173
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1667941163
transform 1 0 17756 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1667941163
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1667941163
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_217
timestamp 1667941163
transform 1 0 21068 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_226
timestamp 1667941163
transform 1 0 21896 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_232
timestamp 1667941163
transform 1 0 22448 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1667941163
transform 1 0 23276 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1667941163
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_263
timestamp 1667941163
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_275
timestamp 1667941163
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_287
timestamp 1667941163
transform 1 0 27508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_299
timestamp 1667941163
transform 1 0 28612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1667941163
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1667941163
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1667941163
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1667941163
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1667941163
transform 1 0 2668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_42
timestamp 1667941163
transform 1 0 4968 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1667941163
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1667941163
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1667941163
transform 1 0 8372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_86
timestamp 1667941163
transform 1 0 9016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1667941163
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp 1667941163
transform 1 0 12972 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_142
timestamp 1667941163
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_155
timestamp 1667941163
transform 1 0 15364 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1667941163
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_186
timestamp 1667941163
transform 1 0 18216 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_195
timestamp 1667941163
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1667941163
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_209
timestamp 1667941163
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1667941163
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_256
timestamp 1667941163
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_263
timestamp 1667941163
transform 1 0 25300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 1667941163
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1667941163
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1667941163
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1667941163
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1667941163
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_353
timestamp 1667941163
transform 1 0 33580 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_357
timestamp 1667941163
transform 1 0 33948 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_369
timestamp 1667941163
transform 1 0 35052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1667941163
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1667941163
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_401
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_12
timestamp 1667941163
transform 1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1667941163
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1667941163
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_57
timestamp 1667941163
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1667941163
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1667941163
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_95
timestamp 1667941163
transform 1 0 9844 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_101
timestamp 1667941163
transform 1 0 10396 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 1667941163
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1667941163
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_119
timestamp 1667941163
transform 1 0 12052 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1667941163
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 1667941163
transform 1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1667941163
transform 1 0 16100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_176
timestamp 1667941163
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1667941163
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_209
timestamp 1667941163
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_217
timestamp 1667941163
transform 1 0 21068 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1667941163
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_233
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_258
timestamp 1667941163
transform 1 0 24840 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_270
timestamp 1667941163
transform 1 0 25944 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_282
timestamp 1667941163
transform 1 0 27048 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_294
timestamp 1667941163
transform 1 0 28152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1667941163
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1667941163
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1667941163
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1667941163
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1667941163
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1667941163
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1667941163
transform 1 0 3496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1667941163
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1667941163
transform 1 0 4784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1667941163
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1667941163
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1667941163
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_65
timestamp 1667941163
transform 1 0 7084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_78
timestamp 1667941163
transform 1 0 8280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1667941163
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_103
timestamp 1667941163
transform 1 0 10580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1667941163
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_124
timestamp 1667941163
transform 1 0 12512 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_138
timestamp 1667941163
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_142
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_146
timestamp 1667941163
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1667941163
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1667941163
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1667941163
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1667941163
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_208
timestamp 1667941163
transform 1 0 20240 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_216
timestamp 1667941163
transform 1 0 20976 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1667941163
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1667941163
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_243
timestamp 1667941163
transform 1 0 23460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_250
timestamp 1667941163
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_257
timestamp 1667941163
transform 1 0 24748 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_277
timestamp 1667941163
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1667941163
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1667941163
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1667941163
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1667941163
transform 1 0 5888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1667941163
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_66
timestamp 1667941163
transform 1 0 7176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1667941163
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_96
timestamp 1667941163
transform 1 0 9936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_120
timestamp 1667941163
transform 1 0 12144 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1667941163
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1667941163
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1667941163
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_160
timestamp 1667941163
transform 1 0 15824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_164
timestamp 1667941163
transform 1 0 16192 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_168
timestamp 1667941163
transform 1 0 16560 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_175
timestamp 1667941163
transform 1 0 17204 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_182
timestamp 1667941163
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_207
timestamp 1667941163
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_214
timestamp 1667941163
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_230
timestamp 1667941163
transform 1 0 22264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_234
timestamp 1667941163
transform 1 0 22632 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_240
timestamp 1667941163
transform 1 0 23184 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1667941163
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1667941163
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1667941163
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1667941163
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1667941163
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1667941163
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_30
timestamp 1667941163
transform 1 0 3864 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_38
timestamp 1667941163
transform 1 0 4600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_42
timestamp 1667941163
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_68
timestamp 1667941163
transform 1 0 7360 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1667941163
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_86
timestamp 1667941163
transform 1 0 9016 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_124
timestamp 1667941163
transform 1 0 12512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_133
timestamp 1667941163
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_145
timestamp 1667941163
transform 1 0 14444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_151
timestamp 1667941163
transform 1 0 14996 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1667941163
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_179
timestamp 1667941163
transform 1 0 17572 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_187
timestamp 1667941163
transform 1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_197
timestamp 1667941163
transform 1 0 19228 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_201
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1667941163
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1667941163
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1667941163
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1667941163
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_258
timestamp 1667941163
transform 1 0 24840 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_265
timestamp 1667941163
transform 1 0 25484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_272
timestamp 1667941163
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1667941163
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1667941163
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1667941163
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1667941163
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_39
timestamp 1667941163
transform 1 0 4692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_64
timestamp 1667941163
transform 1 0 6992 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_70
timestamp 1667941163
transform 1 0 7544 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1667941163
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1667941163
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1667941163
transform 1 0 12972 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1667941163
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1667941163
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1667941163
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1667941163
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1667941163
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1667941163
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_202
timestamp 1667941163
transform 1 0 19688 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_208
timestamp 1667941163
transform 1 0 20240 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_216
timestamp 1667941163
transform 1 0 20976 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_220
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1667941163
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1667941163
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_268
timestamp 1667941163
transform 1 0 25760 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_275
timestamp 1667941163
transform 1 0 26404 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_287
timestamp 1667941163
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1667941163
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1667941163
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1667941163
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_28
timestamp 1667941163
transform 1 0 3680 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_89
timestamp 1667941163
transform 1 0 9292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1667941163
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1667941163
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_121
timestamp 1667941163
transform 1 0 12236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_128
timestamp 1667941163
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1667941163
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_142
timestamp 1667941163
transform 1 0 14168 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1667941163
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_175
timestamp 1667941163
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_188
timestamp 1667941163
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_195
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_208
timestamp 1667941163
transform 1 0 20240 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1667941163
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_231
timestamp 1667941163
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1667941163
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_244
timestamp 1667941163
transform 1 0 23552 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_248
timestamp 1667941163
transform 1 0 23920 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_256
timestamp 1667941163
transform 1 0 24656 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1667941163
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1667941163
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1667941163
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1667941163
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1667941163
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1667941163
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_54
timestamp 1667941163
transform 1 0 6072 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1667941163
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_95
timestamp 1667941163
transform 1 0 9844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_119
timestamp 1667941163
transform 1 0 12052 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1667941163
transform 1 0 12604 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_157
timestamp 1667941163
transform 1 0 15548 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1667941163
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_173
timestamp 1667941163
transform 1 0 17020 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_188
timestamp 1667941163
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_202
timestamp 1667941163
transform 1 0 19688 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_216
timestamp 1667941163
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1667941163
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_227
timestamp 1667941163
transform 1 0 21988 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1667941163
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_238
timestamp 1667941163
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1667941163
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1667941163
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_272
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_279
timestamp 1667941163
transform 1 0 26772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_286
timestamp 1667941163
transform 1 0 27416 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_293
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1667941163
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1667941163
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1667941163
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_405
timestamp 1667941163
transform 1 0 38364 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_8
timestamp 1667941163
transform 1 0 1840 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_37
timestamp 1667941163
transform 1 0 4508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_44
timestamp 1667941163
transform 1 0 5152 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_50
timestamp 1667941163
transform 1 0 5704 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1667941163
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_76
timestamp 1667941163
transform 1 0 8096 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_100
timestamp 1667941163
transform 1 0 10304 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_106
timestamp 1667941163
transform 1 0 10856 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_122
timestamp 1667941163
transform 1 0 12328 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_129
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1667941163
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1667941163
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_182
timestamp 1667941163
transform 1 0 17848 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_188
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_192
timestamp 1667941163
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_196
timestamp 1667941163
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_200
timestamp 1667941163
transform 1 0 19504 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1667941163
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_237
timestamp 1667941163
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_252
timestamp 1667941163
transform 1 0 24288 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_259
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1667941163
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1667941163
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1667941163
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_353
timestamp 1667941163
transform 1 0 33580 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_357
timestamp 1667941163
transform 1 0 33948 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_369
timestamp 1667941163
transform 1 0 35052 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_381
timestamp 1667941163
transform 1 0 36156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1667941163
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_58
timestamp 1667941163
transform 1 0 6440 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_69
timestamp 1667941163
transform 1 0 7452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1667941163
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_96
timestamp 1667941163
transform 1 0 9936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_132
timestamp 1667941163
transform 1 0 13248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_156
timestamp 1667941163
transform 1 0 15456 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_170
timestamp 1667941163
transform 1 0 16744 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_187
timestamp 1667941163
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1667941163
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1667941163
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_221
timestamp 1667941163
transform 1 0 21436 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_225
timestamp 1667941163
transform 1 0 21804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_229
timestamp 1667941163
transform 1 0 22172 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_235
timestamp 1667941163
transform 1 0 22724 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1667941163
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_263
timestamp 1667941163
transform 1 0 25300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1667941163
transform 1 0 25944 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1667941163
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1667941163
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1667941163
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1667941163
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_329
timestamp 1667941163
transform 1 0 31372 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_335
timestamp 1667941163
transform 1 0 31924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_347
timestamp 1667941163
transform 1 0 33028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 1667941163
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_37
timestamp 1667941163
transform 1 0 4508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_44
timestamp 1667941163
transform 1 0 5152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1667941163
transform 1 0 6808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_66
timestamp 1667941163
transform 1 0 7176 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_70
timestamp 1667941163
transform 1 0 7544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_89
timestamp 1667941163
transform 1 0 9292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_128
timestamp 1667941163
transform 1 0 12880 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_136
timestamp 1667941163
transform 1 0 13616 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1667941163
transform 1 0 14536 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_159
timestamp 1667941163
transform 1 0 15732 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_174
timestamp 1667941163
transform 1 0 17112 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1667941163
transform 1 0 17848 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1667941163
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_203
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_210
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_218
timestamp 1667941163
transform 1 0 21160 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1667941163
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1667941163
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1667941163
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_261
timestamp 1667941163
transform 1 0 25116 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_268
timestamp 1667941163
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1667941163
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1667941163
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1667941163
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_342
timestamp 1667941163
transform 1 0 32568 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_354
timestamp 1667941163
transform 1 0 33672 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_366
timestamp 1667941163
transform 1 0 34776 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_378
timestamp 1667941163
transform 1 0 35880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1667941163
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_8
timestamp 1667941163
transform 1 0 1840 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_17
timestamp 1667941163
transform 1 0 2668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_21
timestamp 1667941163
transform 1 0 3036 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1667941163
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_34
timestamp 1667941163
transform 1 0 4232 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_40
timestamp 1667941163
transform 1 0 4784 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_49
timestamp 1667941163
transform 1 0 5612 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_56
timestamp 1667941163
transform 1 0 6256 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_69
timestamp 1667941163
transform 1 0 7452 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1667941163
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_106
timestamp 1667941163
transform 1 0 10856 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_113
timestamp 1667941163
transform 1 0 11500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_125
timestamp 1667941163
transform 1 0 12604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_151
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_158
timestamp 1667941163
transform 1 0 15640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_173
timestamp 1667941163
transform 1 0 17020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1667941163
transform 1 0 17848 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1667941163
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1667941163
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1667941163
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_222
timestamp 1667941163
transform 1 0 21528 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1667941163
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_263
timestamp 1667941163
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_275
timestamp 1667941163
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_287
timestamp 1667941163
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1667941163
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1667941163
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1667941163
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1667941163
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1667941163
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_10
timestamp 1667941163
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_14
timestamp 1667941163
transform 1 0 2392 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_18
timestamp 1667941163
transform 1 0 2760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_25
timestamp 1667941163
transform 1 0 3404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_29
timestamp 1667941163
transform 1 0 3772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_33
timestamp 1667941163
transform 1 0 4140 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_40
timestamp 1667941163
transform 1 0 4784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1667941163
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_63
timestamp 1667941163
transform 1 0 6900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_67
timestamp 1667941163
transform 1 0 7268 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_74
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_86
timestamp 1667941163
transform 1 0 9016 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_91
timestamp 1667941163
transform 1 0 9476 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_99
timestamp 1667941163
transform 1 0 10212 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_103
timestamp 1667941163
transform 1 0 10580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1667941163
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_120
timestamp 1667941163
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_127
timestamp 1667941163
transform 1 0 12788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_134
timestamp 1667941163
transform 1 0 13432 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1667941163
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_148
timestamp 1667941163
transform 1 0 14720 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_174
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_178
timestamp 1667941163
transform 1 0 17480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_182
timestamp 1667941163
transform 1 0 17848 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_191
timestamp 1667941163
transform 1 0 18676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_198
timestamp 1667941163
transform 1 0 19320 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_206
timestamp 1667941163
transform 1 0 20056 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_212
timestamp 1667941163
transform 1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_219
timestamp 1667941163
transform 1 0 21252 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1667941163
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1667941163
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_242
timestamp 1667941163
transform 1 0 23368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1667941163
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1667941163
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_263
timestamp 1667941163
transform 1 0 25300 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1667941163
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1667941163
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1667941163
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1667941163
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_9
timestamp 1667941163
transform 1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_16
timestamp 1667941163
transform 1 0 2576 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_46
timestamp 1667941163
transform 1 0 5336 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_58
timestamp 1667941163
transform 1 0 6440 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_64
timestamp 1667941163
transform 1 0 6992 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_71
timestamp 1667941163
transform 1 0 7636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_113
timestamp 1667941163
transform 1 0 11500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_117
timestamp 1667941163
transform 1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1667941163
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_131
timestamp 1667941163
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_157
timestamp 1667941163
transform 1 0 15548 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_163
timestamp 1667941163
transform 1 0 16100 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_172
timestamp 1667941163
transform 1 0 16928 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_184
timestamp 1667941163
transform 1 0 18032 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_205
timestamp 1667941163
transform 1 0 19964 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1667941163
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1667941163
transform 1 0 22080 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_232
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_241
timestamp 1667941163
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1667941163
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_258
timestamp 1667941163
transform 1 0 24840 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_270
timestamp 1667941163
transform 1 0 25944 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_282
timestamp 1667941163
transform 1 0 27048 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_294
timestamp 1667941163
transform 1 0 28152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1667941163
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1667941163
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1667941163
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1667941163
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_401
timestamp 1667941163
transform 1 0 37996 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1667941163
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_68
timestamp 1667941163
transform 1 0 7360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1667941163
transform 1 0 8464 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_92
timestamp 1667941163
transform 1 0 9568 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1667941163
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_119
timestamp 1667941163
transform 1 0 12052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1667941163
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_133
timestamp 1667941163
transform 1 0 13340 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_145
timestamp 1667941163
transform 1 0 14444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp 1667941163
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_180
timestamp 1667941163
transform 1 0 17664 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_192
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_204
timestamp 1667941163
transform 1 0 19872 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_208
timestamp 1667941163
transform 1 0 20240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_244
timestamp 1667941163
transform 1 0 23552 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_256
timestamp 1667941163
transform 1 0 24656 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_268
timestamp 1667941163
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1667941163
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1667941163
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1667941163
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1667941163
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_353
timestamp 1667941163
transform 1 0 33580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_365
timestamp 1667941163
transform 1 0 34684 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_377
timestamp 1667941163
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1667941163
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_8
timestamp 1667941163
transform 1 0 1840 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1667941163
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_45
timestamp 1667941163
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_57
timestamp 1667941163
transform 1 0 6348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_69
timestamp 1667941163
transform 1 0 7452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1667941163
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_93
timestamp 1667941163
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1667941163
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_151
timestamp 1667941163
transform 1 0 14996 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_169
timestamp 1667941163
transform 1 0 16652 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_176
timestamp 1667941163
transform 1 0 17296 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1667941163
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_212
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_224
timestamp 1667941163
transform 1 0 21712 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_236
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1667941163
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1667941163
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1667941163
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1667941163
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1667941163
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1667941163
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1667941163
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1667941163
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_401
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_101
timestamp 1667941163
transform 1 0 10396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1667941163
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_119
timestamp 1667941163
transform 1 0 12052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_126
timestamp 1667941163
transform 1 0 12696 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_134
timestamp 1667941163
transform 1 0 13432 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_138
timestamp 1667941163
transform 1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_145
timestamp 1667941163
transform 1 0 14444 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_153
timestamp 1667941163
transform 1 0 15180 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_157
timestamp 1667941163
transform 1 0 15548 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1667941163
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_174
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1667941163
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1667941163
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_241
timestamp 1667941163
transform 1 0 23276 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_245
timestamp 1667941163
transform 1 0 23644 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_257
timestamp 1667941163
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1667941163
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1667941163
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1667941163
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1667941163
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_356
timestamp 1667941163
transform 1 0 33856 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_368
timestamp 1667941163
transform 1 0 34960 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_380
timestamp 1667941163
transform 1 0 36064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_386
timestamp 1667941163
transform 1 0 36616 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1667941163
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_117
timestamp 1667941163
transform 1 0 11868 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_122
timestamp 1667941163
transform 1 0 12328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_129
timestamp 1667941163
transform 1 0 12972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1667941163
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_164
timestamp 1667941163
transform 1 0 16192 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_172
timestamp 1667941163
transform 1 0 16928 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_176
timestamp 1667941163
transform 1 0 17296 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1667941163
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_215
timestamp 1667941163
transform 1 0 20884 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_219
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_231
timestamp 1667941163
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1667941163
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1667941163
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_62
timestamp 1667941163
transform 1 0 6808 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_74
timestamp 1667941163
transform 1 0 7912 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_86
timestamp 1667941163
transform 1 0 9016 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_98
timestamp 1667941163
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1667941163
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_205
timestamp 1667941163
transform 1 0 19964 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_216
timestamp 1667941163
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_293
timestamp 1667941163
transform 1 0 28060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_301
timestamp 1667941163
transform 1 0 28796 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_307
timestamp 1667941163
transform 1 0 29348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_319
timestamp 1667941163
transform 1 0 30452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1667941163
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1667941163
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_8
timestamp 1667941163
transform 1 0 1840 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1667941163
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1667941163
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1667941163
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1667941163
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_217
timestamp 1667941163
transform 1 0 21068 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_229
timestamp 1667941163
transform 1 0 22172 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_241
timestamp 1667941163
transform 1 0 23276 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1667941163
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1667941163
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1667941163
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_33
timestamp 1667941163
transform 1 0 4140 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_37
timestamp 1667941163
transform 1 0 4508 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_49
timestamp 1667941163
transform 1 0 5612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1667941163
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1667941163
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1667941163
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1667941163
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1667941163
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1667941163
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1667941163
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1667941163
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1667941163
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1667941163
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_317
timestamp 1667941163
transform 1 0 30268 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_321
timestamp 1667941163
transform 1 0 30636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_333
timestamp 1667941163
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_47
timestamp 1667941163
transform 1 0 5428 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_51
timestamp 1667941163
transform 1 0 5796 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_63
timestamp 1667941163
transform 1 0 6900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_75
timestamp 1667941163
transform 1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_176
timestamp 1667941163
transform 1 0 17296 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_188
timestamp 1667941163
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1667941163
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1667941163
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1667941163
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1667941163
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_341
timestamp 1667941163
transform 1 0 32476 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_347
timestamp 1667941163
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_359
timestamp 1667941163
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1667941163
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_8
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_20
timestamp 1667941163
transform 1 0 2944 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_32
timestamp 1667941163
transform 1 0 4048 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_44
timestamp 1667941163
transform 1 0 5152 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_144
timestamp 1667941163
transform 1 0 14352 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_156
timestamp 1667941163
transform 1 0 15456 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_180
timestamp 1667941163
transform 1 0 17664 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_192
timestamp 1667941163
transform 1 0 18768 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_204
timestamp 1667941163
transform 1 0 19872 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1667941163
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1667941163
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1667941163
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_286
timestamp 1667941163
transform 1 0 27416 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_298
timestamp 1667941163
transform 1 0 28520 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_310
timestamp 1667941163
transform 1 0 29624 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_322
timestamp 1667941163
transform 1 0 30728 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1667941163
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_58
timestamp 1667941163
transform 1 0 6440 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_70
timestamp 1667941163
transform 1 0 7544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1667941163
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1667941163
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_151
timestamp 1667941163
transform 1 0 14996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_163
timestamp 1667941163
transform 1 0 16100 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_174
timestamp 1667941163
transform 1 0 17112 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_186
timestamp 1667941163
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1667941163
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1667941163
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1667941163
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1667941163
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1667941163
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_371
timestamp 1667941163
transform 1 0 35236 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_383
timestamp 1667941163
transform 1 0 36340 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_395
timestamp 1667941163
transform 1 0 37444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_87
timestamp 1667941163
transform 1 0 9108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_99
timestamp 1667941163
transform 1 0 10212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1667941163
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1667941163
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1667941163
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_316
timestamp 1667941163
transform 1 0 30176 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_328
timestamp 1667941163
transform 1 0 31280 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_8
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1667941163
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1667941163
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1667941163
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1667941163
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1667941163
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1667941163
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_257
timestamp 1667941163
transform 1 0 24748 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_261
timestamp 1667941163
transform 1 0 25116 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_273
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_285
timestamp 1667941163
transform 1 0 27324 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_297
timestamp 1667941163
transform 1 0 28428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1667941163
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_314
timestamp 1667941163
transform 1 0 29992 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_326
timestamp 1667941163
transform 1 0 31096 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_338
timestamp 1667941163
transform 1 0 32200 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_350
timestamp 1667941163
transform 1 0 33304 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1667941163
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_370
timestamp 1667941163
transform 1 0 35144 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_382
timestamp 1667941163
transform 1 0 36248 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_394
timestamp 1667941163
transform 1 0 37352 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1667941163
transform 1 0 38456 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_102
timestamp 1667941163
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1667941163
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_141
timestamp 1667941163
transform 1 0 14076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_153
timestamp 1667941163
transform 1 0 15180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_165
timestamp 1667941163
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1667941163
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1667941163
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_286
timestamp 1667941163
transform 1 0 27416 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_298
timestamp 1667941163
transform 1 0 28520 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_310
timestamp 1667941163
transform 1 0 29624 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_322
timestamp 1667941163
transform 1 0 30728 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_334
timestamp 1667941163
transform 1 0 31832 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1667941163
transform 1 0 6348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_61
timestamp 1667941163
transform 1 0 6716 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_73
timestamp 1667941163
transform 1 0 7820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_81
timestamp 1667941163
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_117
timestamp 1667941163
transform 1 0 11868 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_122
timestamp 1667941163
transform 1 0 12328 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1667941163
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_218
timestamp 1667941163
transform 1 0 21160 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_230
timestamp 1667941163
transform 1 0 22264 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_242
timestamp 1667941163
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1667941163
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1667941163
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1667941163
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1667941163
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_20
timestamp 1667941163
transform 1 0 2944 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1667941163
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1667941163
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_52
timestamp 1667941163
transform 1 0 5888 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_64
timestamp 1667941163
transform 1 0 6992 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_76
timestamp 1667941163
transform 1 0 8096 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_285
timestamp 1667941163
transform 1 0 27324 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_290
timestamp 1667941163
transform 1 0 27784 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1667941163
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_8
timestamp 1667941163
transform 1 0 1840 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_20
timestamp 1667941163
transform 1 0 2944 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_32
timestamp 1667941163
transform 1 0 4048 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_44
timestamp 1667941163
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1667941163
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1667941163
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1667941163
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1667941163
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_401
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1667941163
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1667941163
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1667941163
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1667941163
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1667941163
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_146
timestamp 1667941163
transform 1 0 14536 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_158
timestamp 1667941163
transform 1 0 15640 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_162
timestamp 1667941163
transform 1 0 16008 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_174
timestamp 1667941163
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1667941163
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1667941163
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_237
timestamp 1667941163
transform 1 0 22908 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_241
timestamp 1667941163
transform 1 0 23276 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1667941163
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_259
timestamp 1667941163
transform 1 0 24932 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_263
timestamp 1667941163
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_275
timestamp 1667941163
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_287
timestamp 1667941163
transform 1 0 27508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_291
timestamp 1667941163
transform 1 0 27876 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_295
timestamp 1667941163
transform 1 0 28244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1667941163
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_47
timestamp 1667941163
transform 1 0 5428 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_61
timestamp 1667941163
transform 1 0 6716 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_65
timestamp 1667941163
transform 1 0 7084 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_77
timestamp 1667941163
transform 1 0 8188 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_89
timestamp 1667941163
transform 1 0 9292 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_101
timestamp 1667941163
transform 1 0 10396 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1667941163
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_145
timestamp 1667941163
transform 1 0 14444 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_150
timestamp 1667941163
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1667941163
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1667941163
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_177
timestamp 1667941163
transform 1 0 17388 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_183
timestamp 1667941163
transform 1 0 17940 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_191
timestamp 1667941163
transform 1 0 18676 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_195
timestamp 1667941163
transform 1 0 19044 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_207
timestamp 1667941163
transform 1 0 20148 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1667941163
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_285
timestamp 1667941163
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_289
timestamp 1667941163
transform 1 0 27692 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_301
timestamp 1667941163
transform 1 0 28796 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_313
timestamp 1667941163
transform 1 0 29900 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_325
timestamp 1667941163
transform 1 0 31004 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1667941163
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1667941163
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_159
timestamp 1667941163
transform 1 0 15732 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_171
timestamp 1667941163
transform 1 0 16836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_183
timestamp 1667941163
transform 1 0 17940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_256
timestamp 1667941163
transform 1 0 24656 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_268
timestamp 1667941163
transform 1 0 25760 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_35
timestamp 1667941163
transform 1 0 4324 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_47
timestamp 1667941163
transform 1 0 5428 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_59
timestamp 1667941163
transform 1 0 6532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_71
timestamp 1667941163
transform 1 0 7636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_113
timestamp 1667941163
transform 1 0 11500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_117
timestamp 1667941163
transform 1 0 11868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_129
timestamp 1667941163
transform 1 0 12972 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 1667941163
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_314
timestamp 1667941163
transform 1 0 29992 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_326
timestamp 1667941163
transform 1 0 31096 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_338
timestamp 1667941163
transform 1 0 32200 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_350
timestamp 1667941163
transform 1 0 33304 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1667941163
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_370
timestamp 1667941163
transform 1 0 35144 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_382
timestamp 1667941163
transform 1 0 36248 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_394
timestamp 1667941163
transform 1 0 37352 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_21
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_25
timestamp 1667941163
transform 1 0 3404 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_29
timestamp 1667941163
transform 1 0 3772 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_37
timestamp 1667941163
transform 1 0 4508 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_42
timestamp 1667941163
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1667941163
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_266
timestamp 1667941163
transform 1 0 25576 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1667941163
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_333
timestamp 1667941163
transform 1 0 31740 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_345
timestamp 1667941163
transform 1 0 32844 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_382
timestamp 1667941163
transform 1 0 36248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_386
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1667941163
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1667941163
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_71
timestamp 1667941163
transform 1 0 7636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1667941163
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_90
timestamp 1667941163
transform 1 0 9384 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_98
timestamp 1667941163
transform 1 0 10120 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_121
timestamp 1667941163
transform 1 0 12236 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1667941163
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1667941163
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_238
timestamp 1667941163
transform 1 0 23000 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1667941163
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1667941163
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_289
timestamp 1667941163
transform 1 0 27692 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1667941163
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_322
timestamp 1667941163
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1667941163
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_350
timestamp 1667941163
transform 1 0 33304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_356
timestamp 1667941163
transform 1 0 33856 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_383
timestamp 1667941163
transform 1 0 36340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1667941163
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0416_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0417_
timestamp 1667941163
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0419_
timestamp 1667941163
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 18492 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 18400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 20056 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 10948 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0429_
timestamp 1667941163
transform 1 0 11776 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0431_
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0432_
timestamp 1667941163
transform 1 0 10304 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0434_
timestamp 1667941163
transform 1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0435_
timestamp 1667941163
transform 1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 9752 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0437_
timestamp 1667941163
transform 1 0 12420 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 12696 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 24380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 24656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 25484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 23736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 25668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 19504 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1667941163
transform 1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0449_
timestamp 1667941163
transform 1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0450_
timestamp 1667941163
transform 1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1667941163
transform 1 0 12880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1667941163
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0455_
timestamp 1667941163
transform 1 0 11960 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 19044 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0458_
timestamp 1667941163
transform 1 0 12420 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0459_
timestamp 1667941163
transform 1 0 13064 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0460_
timestamp 1667941163
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0461_
timestamp 1667941163
transform 1 0 21160 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 21160 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0464_
timestamp 1667941163
transform 1 0 22724 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 25300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0466_
timestamp 1667941163
transform 1 0 13800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0468_
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 9660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 13156 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 14444 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 4508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 4876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0476_
timestamp 1667941163
transform 1 0 7084 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0477_
timestamp 1667941163
transform 1 0 7360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0480_
timestamp 1667941163
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0481_
timestamp 1667941163
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0482_
timestamp 1667941163
transform 1 0 15088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0483_
timestamp 1667941163
transform 1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 18768 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0486_
timestamp 1667941163
transform 1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0487_
timestamp 1667941163
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0488_
timestamp 1667941163
transform 1 0 15548 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0489_
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 13248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 11224 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0492_
timestamp 1667941163
transform 1 0 11776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0493_
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0494_
timestamp 1667941163
transform 1 0 12328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0495_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 10488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0498_
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0499_
timestamp 1667941163
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0500_
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0501_
timestamp 1667941163
transform 1 0 8740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 5520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 7636 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0504_
timestamp 1667941163
transform 1 0 4968 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0505_
timestamp 1667941163
transform 1 0 4968 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0506_
timestamp 1667941163
transform 1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0507_
timestamp 1667941163
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0510_
timestamp 1667941163
transform 1 0 9568 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0511_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0512_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0513_
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0516_
timestamp 1667941163
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0517_
timestamp 1667941163
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0518_
timestamp 1667941163
transform 1 0 18032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0519_
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0521_
timestamp 1667941163
transform 1 0 13156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0522_
timestamp 1667941163
transform 1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0525_
timestamp 1667941163
transform 1 0 17480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0526_
timestamp 1667941163
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0527_
timestamp 1667941163
transform 1 0 11500 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0528_
timestamp 1667941163
transform 1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 13524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0530_
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0531_
timestamp 1667941163
transform 1 0 14536 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 15364 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 11592 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0534_
timestamp 1667941163
transform 1 0 12512 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0535_
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0536_
timestamp 1667941163
transform 1 0 16008 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0537_
timestamp 1667941163
transform 1 0 13892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 13064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0539_
timestamp 1667941163
transform 1 0 14444 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0540_
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 23828 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 22080 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0543_
timestamp 1667941163
transform 1 0 21068 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0544_
timestamp 1667941163
transform 1 0 21344 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0545_
timestamp 1667941163
transform 1 0 25208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0546_
timestamp 1667941163
transform 1 0 24472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 24564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0548_
timestamp 1667941163
transform 1 0 22080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0549_
timestamp 1667941163
transform 1 0 22080 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 15272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 10580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0552_
timestamp 1667941163
transform 1 0 12052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1667941163
transform 1 0 11776 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0554_
timestamp 1667941163
transform 1 0 15916 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1667941163
transform 1 0 17020 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0558_
timestamp 1667941163
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 13432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_
timestamp 1667941163
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0563_
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1667941163
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1667941163
transform 1 0 20056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0570_
timestamp 1667941163
transform 1 0 23644 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0571_
timestamp 1667941163
transform 1 0 25944 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0572_
timestamp 1667941163
transform 1 0 20516 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0573_
timestamp 1667941163
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 19228 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0575_
timestamp 1667941163
transform 1 0 20148 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0576_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 25208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1667941163
transform 1 0 23644 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1667941163
transform 1 0 22724 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0581_
timestamp 1667941163
transform 1 0 26128 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0582_
timestamp 1667941163
transform 1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0584_
timestamp 1667941163
transform 1 0 26496 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0585_
timestamp 1667941163
transform 1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 26404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0588_
timestamp 1667941163
transform 1 0 26496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0589_
timestamp 1667941163
transform 1 0 26772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0590_
timestamp 1667941163
transform 1 0 25576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0591_
timestamp 1667941163
transform 1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0593_
timestamp 1667941163
transform 1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0594_
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1667941163
transform 1 0 22356 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1667941163
transform 1 0 22080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0599_
timestamp 1667941163
transform 1 0 25208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0600_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0602_
timestamp 1667941163
transform 1 0 24656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0603_
timestamp 1667941163
transform 1 0 23368 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 6808 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0606_
timestamp 1667941163
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0607_
timestamp 1667941163
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0608_
timestamp 1667941163
transform 1 0 8740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0609_
timestamp 1667941163
transform 1 0 10304 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0611_
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0612_
timestamp 1667941163
transform 1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 7176 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0615_
timestamp 1667941163
transform 1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0616_
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 1667941163
transform 1 0 8280 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1667941163
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 7268 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0620_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1667941163
transform 1 0 9200 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 7820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 16468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0624_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0625_
timestamp 1667941163
transform 1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0626_
timestamp 1667941163
transform 1 0 7176 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0627_
timestamp 1667941163
transform 1 0 4416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0629_
timestamp 1667941163
transform 1 0 2576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0630_
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0633_
timestamp 1667941163
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0634_
timestamp 1667941163
transform 1 0 19412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0635_
timestamp 1667941163
transform 1 0 22632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0636_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 18952 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0638_
timestamp 1667941163
transform 1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0639_
timestamp 1667941163
transform 1 0 19596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 20516 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 17572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0642_
timestamp 1667941163
transform 1 0 18768 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0643_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0645_
timestamp 1667941163
transform 1 0 21896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 23276 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0647_
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0648_
timestamp 1667941163
transform 1 0 23368 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0651_
timestamp 1667941163
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0652_
timestamp 1667941163
transform 1 0 13248 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0654_
timestamp 1667941163
transform 1 0 11408 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 1667941163
transform 1 0 12696 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0657_
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 20056 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0660_
timestamp 1667941163
transform 1 0 19964 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0661_
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0663_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 20976 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 1667941163
transform 1 0 20792 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0666_
timestamp 1667941163
transform 1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0669_
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0670_
timestamp 1667941163
transform 1 0 20976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 1667941163
transform 1 0 22632 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0672_
timestamp 1667941163
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 26312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0674_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0675_
timestamp 1667941163
transform 1 0 25024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 13064 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0678_
timestamp 1667941163
transform 1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0679_
timestamp 1667941163
transform 1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0680_
timestamp 1667941163
transform 1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0681_
timestamp 1667941163
transform 1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 12420 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0683_
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0684_
timestamp 1667941163
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0687_
timestamp 1667941163
transform 1 0 17480 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0688_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0689_
timestamp 1667941163
transform 1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0690_
timestamp 1667941163
transform 1 0 13800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0692_
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0696_
timestamp 1667941163
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 1667941163
transform 1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 8096 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 1667941163
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 1667941163
transform 1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0702_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0706_
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0707_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0708_
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0709_
timestamp 1667941163
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 29900 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 26220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0714_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 32936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 29716 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 33672 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 24380 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 25116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 29716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 23000 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 14260 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 30544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 33580 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 33764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 30360 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 5612 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 28244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 33856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 29900 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 31004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 27140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 33672 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 17020 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 33488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 28520 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 9936 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 10212 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 32752 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 6164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 13800 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 27508 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 33948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0760_
timestamp 1667941163
transform 1 0 31556 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 33672 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 27784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 35512 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 5520 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 3864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 2300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 33304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 8832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 15732 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 27876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 6440 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 4232 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 16836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 6992 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 29072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 33948 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 14076 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 6532 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 32292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 29716 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 25024 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 27140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 14720 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 6532 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 12052 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 25300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 22724 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 27968 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0806_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0807_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1656 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 4508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1667941163
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0818_
timestamp 1667941163
transform 1 0 2300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 5520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 3956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 2392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0829_
timestamp 1667941163
transform 1 0 3956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0840_
timestamp 1667941163
transform 1 0 1840 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 3128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 3956 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 3128 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 4876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0851_
timestamp 1667941163
transform 1 0 2668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 7176 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 2208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0862_
timestamp 1667941163
transform 1 0 2300 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 4600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1667941163
transform 1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0873_
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 5244 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 4600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1667941163
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1667941163
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1667941163
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1667941163
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1667941163
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1667941163
transform 1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1667941163
transform 1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1667941163
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1667941163
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1667941163
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1667941163
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _0890_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1656 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0891_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2852 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0892_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4232 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0893_
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 4600 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0896_
timestamp 1667941163
transform 1 0 7636 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0897_
timestamp 1667941163
transform 1 0 6532 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0898_
timestamp 1667941163
transform 1 0 1656 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0899_
timestamp 1667941163
transform 1 0 4692 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 4140 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0901_
timestamp 1667941163
transform 1 0 2392 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0902_
timestamp 1667941163
transform 1 0 1656 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0904_
timestamp 1667941163
transform 1 0 2576 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0905_
timestamp 1667941163
transform 1 0 1748 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0906_
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0907_
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0908_
timestamp 1667941163
transform 1 0 8464 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 2576 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0910_
timestamp 1667941163
transform 1 0 6808 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0911_
timestamp 1667941163
transform 1 0 5060 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0913_
timestamp 1667941163
transform 1 0 6532 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0914_
timestamp 1667941163
transform 1 0 2208 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0915_
timestamp 1667941163
transform 1 0 4324 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0916_
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0917_
timestamp 1667941163
transform 1 0 3036 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0918_
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0919_
timestamp 1667941163
transform 1 0 3956 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0920_
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0921_
timestamp 1667941163
transform 1 0 1748 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 1656 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0923_
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0925_
timestamp 1667941163
transform 1 0 3220 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0926_
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0927_
timestamp 1667941163
transform 1 0 1564 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1667941163
transform 1 0 6716 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0929_
timestamp 1667941163
transform 1 0 3956 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0930_
timestamp 1667941163
transform 1 0 9384 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0931_
timestamp 1667941163
transform 1 0 6716 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0933_
timestamp 1667941163
transform 1 0 10304 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0934_
timestamp 1667941163
transform 1 0 6532 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 10212 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0936_
timestamp 1667941163
transform 1 0 4048 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 3956 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0938_
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 1656 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1667941163
transform 1 0 6808 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0942_
timestamp 1667941163
transform 1 0 7176 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0943_
timestamp 1667941163
transform 1 0 7728 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0944_
timestamp 1667941163
transform 1 0 9200 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 10120 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0946_
timestamp 1667941163
transform 1 0 1656 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0947_
timestamp 1667941163
transform 1 0 1656 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0948_
timestamp 1667941163
transform 1 0 10304 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0950_
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0951_
timestamp 1667941163
transform 1 0 8188 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1667941163
transform 1 0 9384 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 9384 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1667941163
transform 1 0 8924 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1667941163
transform 1 0 10304 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 4600 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0957_
timestamp 1667941163
transform 1 0 6164 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1667941163
transform 1 0 9384 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1667941163
transform 1 0 8832 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1667941163
transform 1 0 10304 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1667941163
transform 1 0 9384 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1667941163
transform 1 0 7176 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1667941163
transform 1 0 10396 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1667941163
transform 1 0 9108 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 33580 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1667941163
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 23368 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 11592 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1667941163
transform 1 0 15456 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 35328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 15272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1667941163
transform 1 0 34868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 18768 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1667941163
transform 1 0 32936 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1667941163
transform 1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 14628 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1667941163
transform 1 0 27416 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1667941163
transform 1 0 34684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 33580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 2392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 17664 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 6808 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1667941163
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 5520 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1667941163
transform 1 0 36708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 36156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 35972 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 17664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 25300 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 31464 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1667941163
transform 1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1667941163
transform 1 0 3496 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 27968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1043_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1043__100 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20056 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1044_
timestamp 1667941163
transform 1 0 17940 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1045_
timestamp 1667941163
transform 1 0 19136 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1046_
timestamp 1667941163
transform 1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1047_
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1048_
timestamp 1667941163
transform 1 0 12420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1049__101
timestamp 1667941163
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1049_
timestamp 1667941163
transform 1 0 12236 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1050_
timestamp 1667941163
transform 1 0 7544 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 7452 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1052_
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1053_
timestamp 1667941163
transform 1 0 13064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1054_
timestamp 1667941163
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1055__102
timestamp 1667941163
transform 1 0 18216 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1055_
timestamp 1667941163
transform 1 0 18124 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1056_
timestamp 1667941163
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1057_
timestamp 1667941163
transform 1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1058_
timestamp 1667941163
transform 1 0 18400 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1059_
timestamp 1667941163
transform 1 0 12420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1060_
timestamp 1667941163
transform 1 0 12144 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1061_
timestamp 1667941163
transform 1 0 9292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1061__103
timestamp 1667941163
transform 1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1062_
timestamp 1667941163
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1063_
timestamp 1667941163
transform 1 0 11316 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1064_
timestamp 1667941163
transform 1 0 11868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1065_
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1066_
timestamp 1667941163
transform 1 0 23184 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1067__104
timestamp 1667941163
transform 1 0 24380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1067_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1068_
timestamp 1667941163
transform 1 0 20792 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1069_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1070_
timestamp 1667941163
transform 1 0 24380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1071_
timestamp 1667941163
transform 1 0 17112 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1072_
timestamp 1667941163
transform 1 0 21252 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1073__105
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1073_
timestamp 1667941163
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1074_
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1075_
timestamp 1667941163
transform 1 0 20700 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1076_
timestamp 1667941163
transform 1 0 20148 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1077_
timestamp 1667941163
transform 1 0 20240 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1078_
timestamp 1667941163
transform 1 0 14536 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1079_
timestamp 1667941163
transform 1 0 14536 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1079__106
timestamp 1667941163
transform 1 0 12052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1080_
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1081_
timestamp 1667941163
transform 1 0 15088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1082_
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1083_
timestamp 1667941163
transform 1 0 14904 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1084_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22264 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1085__107
timestamp 1667941163
transform 1 0 22632 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1085_
timestamp 1667941163
transform 1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1086_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1087_
timestamp 1667941163
transform 1 0 19044 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_1  _1088_
timestamp 1667941163
transform 1 0 22540 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1089_
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1090_
timestamp 1667941163
transform 1 0 20792 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1091_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1091__108
timestamp 1667941163
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1092_
timestamp 1667941163
transform 1 0 19596 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1093_
timestamp 1667941163
transform 1 0 20516 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1094_
timestamp 1667941163
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1095_
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1096_
timestamp 1667941163
transform 1 0 7544 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1097__109
timestamp 1667941163
transform 1 0 2576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1097_
timestamp 1667941163
transform 1 0 9568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1098_
timestamp 1667941163
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 7636 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1100_
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1101_
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1102_
timestamp 1667941163
transform 1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1103_
timestamp 1667941163
transform 1 0 9476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1103__110
timestamp 1667941163
transform 1 0 9384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1104_
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1105_
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1106_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1107_
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1108_
timestamp 1667941163
transform 1 0 12788 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1109_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1109__111
timestamp 1667941163
transform 1 0 7268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1110_
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1111_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1112_
timestamp 1667941163
transform 1 0 10120 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1113_
timestamp 1667941163
transform 1 0 9936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1114_
timestamp 1667941163
transform 1 0 23184 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1115__112
timestamp 1667941163
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1115_
timestamp 1667941163
transform 1 0 22264 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1116_
timestamp 1667941163
transform 1 0 21712 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 23000 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1118_
timestamp 1667941163
transform 1 0 22264 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1119_
timestamp 1667941163
transform 1 0 22356 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1120_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1121_
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1121__113
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1122_
timestamp 1667941163
transform 1 0 25668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1123_
timestamp 1667941163
transform 1 0 25300 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1124_
timestamp 1667941163
transform 1 0 23000 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1125_
timestamp 1667941163
transform 1 0 24656 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 24932 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1127__114
timestamp 1667941163
transform 1 0 27140 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1127_
timestamp 1667941163
transform 1 0 24748 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1128_
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1130_
timestamp 1667941163
transform 1 0 24748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1131_
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 17480 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1133_
timestamp 1667941163
transform 1 0 19044 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1133__115
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1134_
timestamp 1667941163
transform 1 0 23368 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 17572 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1136_
timestamp 1667941163
transform 1 0 19412 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1137_
timestamp 1667941163
transform 1 0 22724 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 17572 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1139__116
timestamp 1667941163
transform 1 0 14260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1139_
timestamp 1667941163
transform 1 0 17664 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1140_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 17204 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1142_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1143_
timestamp 1667941163
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1145__117
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1145_
timestamp 1667941163
transform 1 0 15916 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1146_
timestamp 1667941163
transform 1 0 12512 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 14996 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1148_
timestamp 1667941163
transform 1 0 16192 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1149_
timestamp 1667941163
transform 1 0 10396 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1150_
timestamp 1667941163
transform 1 0 23276 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1151_
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1151__118
timestamp 1667941163
transform 1 0 22356 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1152_
timestamp 1667941163
transform 1 0 20608 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1154_
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1155_
timestamp 1667941163
transform 1 0 22172 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1157_
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1157__119
timestamp 1667941163
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1158_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 14904 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1160_
timestamp 1667941163
transform 1 0 15088 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1161_
timestamp 1667941163
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1162_
timestamp 1667941163
transform 1 0 10948 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1163__120
timestamp 1667941163
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1163_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1164_
timestamp 1667941163
transform 1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1165_
timestamp 1667941163
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1166_
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 16100 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 17204 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1169_
timestamp 1667941163
transform 1 0 16468 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1169__121
timestamp 1667941163
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1170_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1171_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1172_
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1173_
timestamp 1667941163
transform 1 0 11684 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1174__122
timestamp 1667941163
transform 1 0 16928 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 17572 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 11776 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1176_
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1177_
timestamp 1667941163
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform 1 0 5152 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1178__123
timestamp 1667941163
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1180_
timestamp 1667941163
transform 1 0 6532 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1181_
timestamp 1667941163
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1182__124
timestamp 1667941163
transform 1 0 8096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1182_
timestamp 1667941163
transform 1 0 11684 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 17940 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 16468 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 17480 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1186_
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1186__125
timestamp 1667941163
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1187_
timestamp 1667941163
transform 1 0 13800 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1188_
timestamp 1667941163
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 12512 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1190_
timestamp 1667941163
transform 1 0 13524 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1190__126
timestamp 1667941163
transform 1 0 15272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 20792 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1192_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 20700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1194_
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1194__127
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 6900 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 13800 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 12052 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1198__128
timestamp 1667941163
transform 1 0 6716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1198_
timestamp 1667941163
transform 1 0 6624 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1199_
timestamp 1667941163
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1200_
timestamp 1667941163
transform 1 0 6164 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1201_
timestamp 1667941163
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1202__129
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1202_
timestamp 1667941163
transform 1 0 15088 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 10028 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1204_
timestamp 1667941163
transform 1 0 14628 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1206__130
timestamp 1667941163
transform 1 0 25668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1206_
timestamp 1667941163
transform 1 0 23460 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 21160 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1208_
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1210__131
timestamp 1667941163
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1210_
timestamp 1667941163
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1212_
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 6440 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1214__132
timestamp 1667941163
transform 1 0 22448 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 21252 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 16376 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1216_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1667941163
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1218__133
timestamp 1667941163
transform 1 0 25024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1220_
timestamp 1667941163
transform 1 0 23368 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 22816 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1222__134
timestamp 1667941163
transform 1 0 13524 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1222_
timestamp 1667941163
transform 1 0 14260 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1223_
timestamp 1667941163
transform 1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1224_
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1225_
timestamp 1667941163
transform 1 0 8832 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1226__135
timestamp 1667941163
transform 1 0 10580 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1226_
timestamp 1667941163
transform 1 0 12052 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1228_
timestamp 1667941163
transform 1 0 12696 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1667941163
transform 1 0 15364 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1230__136
timestamp 1667941163
transform 1 0 19504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1667941163
transform 1 0 17940 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1232_
timestamp 1667941163
transform 1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1667941163
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1234__137
timestamp 1667941163
transform 1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1234_
timestamp 1667941163
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1667941163
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1236_
timestamp 1667941163
transform 1 0 9016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1237_
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 38088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 38088 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 22724 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 36708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 1564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 38088 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 9108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 1564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 1564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 38088 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 36708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1667941163
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 38088 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 38088 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1667941163
transform 1 0 38088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1667941163
transform 1 0 38088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1667941163
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 1564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1667941163
transform 1 0 30452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1667941163
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1667941163
transform 1 0 37996 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 7820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 27784 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 6128 39800 6248 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 2 nsew signal input
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 3 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
port 6 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
port 8 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
port 9 nsew signal input
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 ccff_head
port 10 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal3 s 200 38088 800 38208 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 12 nsew signal input
flabel metal2 s 4526 200 4582 800 0 FreeSans 224 90 0 0 chanx_left_in[10]
port 13 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 14 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 15 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 16 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[14]
port 17 nsew signal input
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 18 nsew signal input
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 19 nsew signal input
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 20 nsew signal input
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 21 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 chanx_left_in[1]
port 22 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_left_in[2]
port 23 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 24 nsew signal input
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 25 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 26 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_left_in[6]
port 27 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_left_in[7]
port 28 nsew signal input
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 29 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chanx_left_in[9]
port 30 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 31 nsew signal tristate
flabel metal3 s 39200 34688 39800 34808 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 32 nsew signal tristate
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chanx_left_out[11]
port 33 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 34 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 35 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chanx_left_out[14]
port 36 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 37 nsew signal tristate
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 38 nsew signal tristate
flabel metal2 s 9034 200 9090 800 0 FreeSans 224 90 0 0 chanx_left_out[17]
port 39 nsew signal tristate
flabel metal3 s 39200 29928 39800 30048 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 40 nsew signal tristate
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 41 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 42 nsew signal tristate
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 43 nsew signal tristate
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 44 nsew signal tristate
flabel metal3 s 39200 1368 39800 1488 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 45 nsew signal tristate
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 46 nsew signal tristate
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chanx_left_out[7]
port 47 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 48 nsew signal tristate
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 49 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal3 s 200 9528 800 9648 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal2 s 36082 200 36138 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal3 s 200 33328 800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal2 s 31574 200 31630 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal2 s 7746 39200 7802 39800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal3 s 200 4768 800 4888 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal2 s 34794 39200 34850 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 88 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 89 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 90 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 91 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 92 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 93 nsew signal input
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
port 94 nsew signal input
flabel metal2 s 30286 39200 30342 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
port 95 nsew signal input
flabel metal2 s 3238 39200 3294 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
port 96 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
port 97 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 pReset
port 98 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 prog_clk
port 99 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 100 nsew signal bidirectional
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 vssd1
port 101 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 101 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 4692 11050 4692 11050 0 _0000_
rlabel metal1 3220 4046 3220 4046 0 _0001_
rlabel metal1 4094 6800 4094 6800 0 _0002_
rlabel metal2 3634 6290 3634 6290 0 _0003_
rlabel metal1 4370 5270 4370 5270 0 _0004_
rlabel metal2 2898 6290 2898 6290 0 _0005_
rlabel metal1 4278 3706 4278 3706 0 _0006_
rlabel metal1 1610 18598 1610 18598 0 _0007_
rlabel metal1 5842 8602 5842 8602 0 _0008_
rlabel metal1 3135 19754 3135 19754 0 _0009_
rlabel metal2 3128 13124 3128 13124 0 _0010_
rlabel metal1 4002 7446 4002 7446 0 _0011_
rlabel metal1 3227 16150 3227 16150 0 _0012_
rlabel metal1 4830 23222 4830 23222 0 _0013_
rlabel metal1 4784 8058 4784 8058 0 _0014_
rlabel metal1 2760 23494 2760 23494 0 _0015_
rlabel metal1 3181 20502 3181 20502 0 _0016_
rlabel metal1 5796 12410 5796 12410 0 _0017_
rlabel metal2 5014 20536 5014 20536 0 _0018_
rlabel metal1 7406 5746 7406 5746 0 _0019_
rlabel metal1 6440 4454 6440 4454 0 _0020_
rlabel metal1 7268 4794 7268 4794 0 _0021_
rlabel metal1 8602 4726 8602 4726 0 _0022_
rlabel metal1 8195 17238 8195 17238 0 _0023_
rlabel via3 11109 20740 11109 20740 0 _0024_
rlabel metal2 3910 4862 3910 4862 0 _0025_
rlabel metal1 2852 4250 2852 4250 0 _0026_
rlabel via3 7843 13804 7843 13804 0 _0027_
rlabel via3 3013 13804 3013 13804 0 _0028_
rlabel metal1 7314 14280 7314 14280 0 _0029_
rlabel metal3 7383 13940 7383 13940 0 _0030_
rlabel metal1 6854 3366 6854 3366 0 _0031_
rlabel metal1 6394 4998 6394 4998 0 _0032_
rlabel metal1 6486 5814 6486 5814 0 _0033_
rlabel metal1 8142 4046 8142 4046 0 _0034_
rlabel metal1 2530 5882 2530 5882 0 _0035_
rlabel metal1 2392 5338 2392 5338 0 _0036_
rlabel metal3 11569 18020 11569 18020 0 _0037_
rlabel metal3 7751 14484 7751 14484 0 _0038_
rlabel metal1 6447 15402 6447 15402 0 _0039_
rlabel metal3 7820 13668 7820 13668 0 _0040_
rlabel metal3 9545 15300 9545 15300 0 _0041_
rlabel via3 10787 19380 10787 19380 0 _0042_
rlabel metal1 5934 4114 5934 4114 0 _0043_
rlabel metal1 9614 5066 9614 5066 0 _0044_
rlabel via3 5451 13804 5451 13804 0 _0045_
rlabel metal1 6118 4794 6118 4794 0 _0046_
rlabel metal3 10649 16660 10649 16660 0 _0047_
rlabel metal3 10327 13804 10327 13804 0 _0048_
rlabel via3 11339 20740 11339 20740 0 _0049_
rlabel metal3 10879 19924 10879 19924 0 _0050_
rlabel metal3 8671 15300 8671 15300 0 _0051_
rlabel metal3 10465 16116 10465 16116 0 _0052_
rlabel metal1 4462 4794 4462 4794 0 _0053_
rlabel metal1 5566 7514 5566 7514 0 _0054_
rlabel metal2 2990 6630 2990 6630 0 _0055_
rlabel metal1 4745 17238 4745 17238 0 _0056_
rlabel metal1 4784 8602 4784 8602 0 _0057_
rlabel metal3 5336 12716 5336 12716 0 _0058_
rlabel metal1 4830 3638 4830 3638 0 _0059_
rlabel metal1 4048 5610 4048 5610 0 _0060_
rlabel metal2 3266 3842 3266 3842 0 _0061_
rlabel metal2 8418 8024 8418 8024 0 _0062_
rlabel via2 1702 8619 1702 8619 0 _0063_
rlabel metal1 2346 6630 2346 6630 0 _0064_
rlabel metal1 1886 10778 1886 10778 0 _0065_
rlabel metal1 1702 10234 1702 10234 0 _0066_
rlabel metal1 4922 12954 4922 12954 0 _0067_
rlabel metal1 4140 10778 4140 10778 0 _0068_
rlabel metal2 3818 11186 3818 11186 0 _0069_
rlabel metal2 2530 12342 2530 12342 0 _0070_
rlabel metal2 2530 7650 2530 7650 0 _0071_
rlabel metal1 3818 12818 3818 12818 0 _0072_
rlabel metal2 9936 14212 9936 14212 0 _0073_
rlabel metal1 4048 5882 4048 5882 0 _0074_
rlabel via3 7613 20740 7613 20740 0 _0075_
rlabel metal1 9154 9418 9154 9418 0 _0076_
rlabel metal1 10304 8602 10304 8602 0 _0077_
rlabel metal2 20102 23494 20102 23494 0 _0078_
rlabel metal1 21114 16218 21114 16218 0 _0079_
rlabel metal2 11362 17850 11362 17850 0 _0080_
rlabel metal1 11178 23732 11178 23732 0 _0081_
rlabel metal2 12650 25670 12650 25670 0 _0082_
rlabel metal1 13570 26384 13570 26384 0 _0083_
rlabel metal2 25530 23188 25530 23188 0 _0084_
rlabel metal1 25208 16082 25208 16082 0 _0085_
rlabel metal1 14076 8602 14076 8602 0 _0086_
rlabel metal2 20562 10438 20562 10438 0 _0087_
rlabel metal1 9890 18938 9890 18938 0 _0088_
rlabel metal1 22126 13260 22126 13260 0 _0089_
rlabel metal1 13294 24752 13294 24752 0 _0090_
rlabel metal2 21482 17340 21482 17340 0 _0091_
rlabel metal1 24150 21114 24150 21114 0 _0092_
rlabel metal1 5106 19482 5106 19482 0 _0093_
rlabel metal1 14306 23698 14306 23698 0 _0094_
rlabel metal1 4554 24038 4554 24038 0 _0095_
rlabel metal2 7590 24378 7590 24378 0 _0096_
rlabel metal1 4002 17646 4002 17646 0 _0097_
rlabel metal1 15962 11152 15962 11152 0 _0098_
rlabel metal1 20562 11866 20562 11866 0 _0099_
rlabel metal2 15594 10438 15594 10438 0 _0100_
rlabel metal2 11822 24378 11822 24378 0 _0101_
rlabel metal2 13018 11662 13018 11662 0 _0102_
rlabel metal1 18630 14314 18630 14314 0 _0103_
rlabel metal2 5842 18428 5842 18428 0 _0104_
rlabel metal2 5198 24956 5198 24956 0 _0105_
rlabel metal1 6578 21998 6578 21998 0 _0106_
rlabel metal2 9338 20434 9338 20434 0 _0107_
rlabel metal1 19228 20434 19228 20434 0 _0108_
rlabel metal1 14720 10030 14720 10030 0 _0109_
rlabel metal1 17848 12206 17848 12206 0 _0110_
rlabel metal1 14582 14314 14582 14314 0 _0111_
rlabel metal1 16928 11730 16928 11730 0 _0112_
rlabel metal1 12374 10064 12374 10064 0 _0113_
rlabel metal1 16146 13430 16146 13430 0 _0114_
rlabel metal1 12834 23834 12834 23834 0 _0115_
rlabel metal1 15364 20298 15364 20298 0 _0116_
rlabel metal1 14444 18938 14444 18938 0 _0117_
rlabel metal1 21344 20026 21344 20026 0 _0118_
rlabel metal1 24978 18258 24978 18258 0 _0119_
rlabel metal1 22218 20570 22218 20570 0 _0120_
rlabel metal2 12006 26044 12006 26044 0 _0121_
rlabel metal2 17250 25874 17250 25874 0 _0122_
rlabel metal2 17710 26044 17710 26044 0 _0123_
rlabel metal2 16330 18428 16330 18428 0 _0124_
rlabel metal1 18262 12954 18262 12954 0 _0125_
rlabel metal1 17710 16966 17710 16966 0 _0126_
rlabel metal1 24288 20570 24288 20570 0 _0127_
rlabel metal2 20562 21726 20562 21726 0 _0128_
rlabel metal2 20194 22916 20194 22916 0 _0129_
rlabel metal2 23690 16252 23690 16252 0 _0130_
rlabel metal2 26082 19516 26082 19516 0 _0131_
rlabel metal2 26542 20604 26542 20604 0 _0132_
rlabel metal1 26772 13498 26772 13498 0 _0133_
rlabel metal2 25622 13124 25622 13124 0 _0134_
rlabel metal1 24610 12818 24610 12818 0 _0135_
rlabel metal1 22356 12954 22356 12954 0 _0136_
rlabel metal1 25024 12206 25024 12206 0 _0137_
rlabel metal1 23598 14960 23598 14960 0 _0138_
rlabel metal2 12558 8636 12558 8636 0 _0139_
rlabel metal1 10534 9588 10534 9588 0 _0140_
rlabel metal1 12742 9928 12742 9928 0 _0141_
rlabel metal1 14766 20468 14766 20468 0 _0142_
rlabel metal1 6854 21522 6854 21522 0 _0143_
rlabel metal1 8924 23290 8924 23290 0 _0144_
rlabel metal1 16468 22066 16468 22066 0 _0145_
rlabel metal2 4646 20604 4646 20604 0 _0146_
rlabel metal1 2691 17510 2691 17510 0 _0147_
rlabel metal1 19872 16762 19872 16762 0 _0148_
rlabel metal1 22448 11730 22448 11730 0 _0149_
rlabel metal1 19642 11730 19642 11730 0 _0150_
rlabel metal2 18814 17476 18814 17476 0 _0151_
rlabel metal2 22034 21828 22034 21828 0 _0152_
rlabel metal2 23598 25466 23598 25466 0 _0153_
rlabel metal1 14168 15130 14168 15130 0 _0154_
rlabel metal2 14674 15963 14674 15963 0 _0155_
rlabel metal1 14674 19822 14674 19822 0 _0156_
rlabel metal2 20562 20026 20562 20026 0 _0157_
rlabel metal2 22034 24310 22034 24310 0 _0158_
rlabel metal2 20930 27132 20930 27132 0 _0159_
rlabel metal1 21206 23732 21206 23732 0 _0160_
rlabel metal1 23092 21658 23092 21658 0 _0161_
rlabel metal2 25254 23868 25254 23868 0 _0162_
rlabel metal2 11638 11594 11638 11594 0 _0163_
rlabel metal1 13248 8058 13248 8058 0 _0164_
rlabel metal1 9476 8942 9476 8942 0 _0165_
rlabel metal1 17296 10642 17296 10642 0 _0166_
rlabel metal1 14490 9146 14490 9146 0 _0167_
rlabel metal2 18722 10234 18722 10234 0 _0168_
rlabel metal1 4830 18258 4830 18258 0 _0169_
rlabel metal1 6026 17204 6026 17204 0 _0170_
rlabel metal1 9200 18258 9200 18258 0 _0171_
rlabel metal1 17158 18700 17158 18700 0 _0172_
rlabel metal2 22586 13736 22586 13736 0 _0173_
rlabel metal1 1610 11730 1610 11730 0 _0174_
rlabel metal1 2208 6766 2208 6766 0 _0175_
rlabel metal2 2530 5899 2530 5899 0 _0176_
rlabel metal1 1794 9520 1794 9520 0 _0177_
rlabel metal1 2346 23698 2346 23698 0 _0178_
rlabel metal1 2254 4148 2254 4148 0 _0179_
rlabel metal1 2392 5202 2392 5202 0 _0180_
rlabel metal1 5750 4148 5750 4148 0 _0181_
rlabel metal1 21436 13498 21436 13498 0 _0182_
rlabel metal1 19412 14042 19412 14042 0 _0183_
rlabel metal2 18170 18428 18170 18428 0 _0184_
rlabel metal1 19918 12954 19918 12954 0 _0185_
rlabel metal1 19044 19278 19044 19278 0 _0186_
rlabel metal1 20792 11322 20792 11322 0 _0187_
rlabel metal2 12650 17884 12650 17884 0 _0188_
rlabel metal1 12466 17068 12466 17068 0 _0189_
rlabel metal2 7774 16031 7774 16031 0 _0190_
rlabel metal2 7682 16354 7682 16354 0 _0191_
rlabel metal1 11638 13294 11638 13294 0 _0192_
rlabel metal1 13294 18326 13294 18326 0 _0193_
rlabel metal2 13846 10710 13846 10710 0 _0194_
rlabel metal1 18446 10234 18446 10234 0 _0195_
rlabel metal1 16284 12750 16284 12750 0 _0196_
rlabel metal3 13938 12852 13938 12852 0 _0197_
rlabel metal1 19090 10234 19090 10234 0 _0198_
rlabel metal3 12650 12444 12650 12444 0 _0199_
rlabel metal2 13018 9656 13018 9656 0 _0200_
rlabel metal1 9614 9146 9614 9146 0 _0201_
rlabel metal1 12328 11322 12328 11322 0 _0202_
rlabel metal1 11684 8602 11684 8602 0 _0203_
rlabel via1 12558 6851 12558 6851 0 _0204_
rlabel metal1 14214 14450 14214 14450 0 _0205_
rlabel metal1 23460 22678 23460 22678 0 _0206_
rlabel metal1 24932 23154 24932 23154 0 _0207_
rlabel metal2 21022 23324 21022 23324 0 _0208_
rlabel metal1 21804 22678 21804 22678 0 _0209_
rlabel metal2 25438 22304 25438 22304 0 _0210_
rlabel metal1 17526 23154 17526 23154 0 _0211_
rlabel metal2 21482 24344 21482 24344 0 _0212_
rlabel metal2 20562 25772 20562 25772 0 _0213_
rlabel metal1 20148 19346 20148 19346 0 _0214_
rlabel metal2 20930 21726 20930 21726 0 _0215_
rlabel metal1 20424 24242 20424 24242 0 _0216_
rlabel metal2 20470 21148 20470 21148 0 _0217_
rlabel metal2 12650 16830 12650 16830 0 _0218_
rlabel metal1 14674 20026 14674 20026 0 _0219_
rlabel metal1 13570 16218 13570 16218 0 _0220_
rlabel metal1 15364 16490 15364 16490 0 _0221_
rlabel metal1 14030 20502 14030 20502 0 _0222_
rlabel metal1 13800 15674 13800 15674 0 _0223_
rlabel metal2 22494 22440 22494 22440 0 _0224_
rlabel metal1 23138 23698 23138 23698 0 _0225_
rlabel metal2 19458 18292 19458 18292 0 _0226_
rlabel metal1 19964 18326 19964 18326 0 _0227_
rlabel metal2 22770 24412 22770 24412 0 _0228_
rlabel metal1 18078 18802 18078 18802 0 _0229_
rlabel metal1 21528 11866 21528 11866 0 _0230_
rlabel metal2 19504 13294 19504 13294 0 _0231_
rlabel metal1 19596 15538 19596 15538 0 _0232_
rlabel metal1 20976 11798 20976 11798 0 _0233_
rlabel metal1 18768 11866 18768 11866 0 _0234_
rlabel metal2 20746 16524 20746 16524 0 _0235_
rlabel viali 7770 18666 7770 18666 0 _0236_
rlabel metal1 3818 14484 3818 14484 0 _0237_
rlabel metal2 15870 21692 15870 21692 0 _0238_
rlabel metal2 7866 20536 7866 20536 0 _0239_
rlabel metal1 11776 11322 11776 11322 0 _0240_
rlabel metal1 16606 20978 16606 20978 0 _0241_
rlabel metal2 7774 19618 7774 19618 0 _0242_
rlabel metal2 9706 23324 9706 23324 0 _0243_
rlabel metal2 15410 20060 15410 20060 0 _0244_
rlabel metal1 7544 18326 7544 18326 0 _0245_
rlabel metal1 9292 17714 9292 17714 0 _0246_
rlabel metal1 16376 19890 16376 19890 0 _0247_
rlabel metal1 13018 15028 13018 15028 0 _0248_
rlabel metal1 12788 10234 12788 10234 0 _0249_
rlabel metal2 12374 10404 12374 10404 0 _0250_
rlabel metal1 12972 9622 12972 9622 0 _0251_
rlabel metal1 9844 12750 9844 12750 0 _0252_
rlabel metal1 7728 10710 7728 10710 0 _0253_
rlabel metal1 24196 12410 24196 12410 0 _0254_
rlabel metal1 22954 14926 22954 14926 0 _0255_
rlabel metal2 22126 14212 22126 14212 0 _0256_
rlabel metal1 24104 12886 24104 12886 0 _0257_
rlabel metal2 24150 15164 24150 15164 0 _0258_
rlabel metal1 23092 12274 23092 12274 0 _0259_
rlabel metal2 25898 13872 25898 13872 0 _0260_
rlabel metal2 24242 13396 24242 13396 0 _0261_
rlabel metal1 26542 14314 26542 14314 0 _0262_
rlabel metal2 26542 14484 26542 14484 0 _0263_
rlabel metal1 23966 14450 23966 14450 0 _0264_
rlabel metal1 25392 13838 25392 13838 0 _0265_
rlabel metal1 25530 19482 25530 19482 0 _0266_
rlabel metal1 25852 20570 25852 20570 0 _0267_
rlabel metal2 22770 16388 22770 16388 0 _0268_
rlabel metal1 24426 17578 24426 17578 0 _0269_
rlabel metal1 25484 20434 25484 20434 0 _0270_
rlabel metal1 23552 17170 23552 17170 0 _0271_
rlabel metal1 18124 21658 18124 21658 0 _0272_
rlabel metal2 19274 22780 19274 22780 0 _0273_
rlabel metal1 23598 21012 23598 21012 0 _0274_
rlabel metal2 18170 20264 18170 20264 0 _0275_
rlabel metal1 19412 21386 19412 21386 0 _0276_
rlabel metal2 22954 18428 22954 18428 0 _0277_
rlabel metal1 17986 14042 17986 14042 0 _0278_
rlabel metal1 17894 17748 17894 17748 0 _0279_
rlabel metal1 16606 18394 16606 18394 0 _0280_
rlabel via2 15594 14603 15594 14603 0 _0281_
rlabel metal1 16652 17306 16652 17306 0 _0282_
rlabel metal1 13386 10778 13386 10778 0 _0283_
rlabel metal2 17066 24990 17066 24990 0 _0284_
rlabel metal1 16836 25330 16836 25330 0 _0285_
rlabel metal2 11822 25500 11822 25500 0 _0286_
rlabel metal2 15226 25262 15226 25262 0 _0287_
rlabel metal1 16698 24242 16698 24242 0 _0288_
rlabel metal2 10626 25500 10626 25500 0 _0289_
rlabel metal1 24518 18360 24518 18360 0 _0290_
rlabel metal2 22494 20026 22494 20026 0 _0291_
rlabel metal1 21114 20434 21114 20434 0 _0292_
rlabel metal1 23782 18394 23782 18394 0 _0293_
rlabel metal2 24702 19652 24702 19652 0 _0294_
rlabel metal2 22402 17612 22402 17612 0 _0295_
rlabel metal1 15410 20536 15410 20536 0 _0296_
rlabel metal1 15318 19244 15318 19244 0 _0297_
rlabel metal2 14490 23596 14490 23596 0 _0298_
rlabel metal2 15134 22814 15134 22814 0 _0299_
rlabel metal2 15272 18802 15272 18802 0 _0300_
rlabel metal2 12098 23596 12098 23596 0 _0301_
rlabel metal1 11592 15470 11592 15470 0 _0302_
rlabel metal1 15824 15674 15824 15674 0 _0303_
rlabel metal1 15732 13838 15732 13838 0 _0304_
rlabel metal1 10902 13838 10902 13838 0 _0305_
rlabel metal2 13662 14688 13662 14688 0 _0306_
rlabel metal1 16468 14382 16468 14382 0 _0307_
rlabel metal2 17434 13362 17434 13362 0 _0308_
rlabel metal1 16836 15470 16836 15470 0 _0309_
rlabel metal1 14398 10234 14398 10234 0 _0310_
rlabel metal1 16376 13498 16376 13498 0 _0311_
rlabel metal2 15318 13396 15318 13396 0 _0312_
rlabel metal1 12834 8058 12834 8058 0 _0313_
rlabel metal1 18446 20570 18446 20570 0 _0314_
rlabel metal2 12006 19652 12006 19652 0 _0315_
rlabel metal1 17388 20026 17388 20026 0 _0316_
rlabel metal1 13294 19958 13294 19958 0 _0317_
rlabel metal2 6210 21760 6210 21760 0 _0318_
rlabel metal1 5060 23154 5060 23154 0 _0319_
rlabel metal1 6670 19414 6670 19414 0 _0320_
rlabel metal1 7912 23494 7912 23494 0 _0321_
rlabel metal2 11914 18904 11914 18904 0 _0322_
rlabel metal1 18308 14586 18308 14586 0 _0323_
rlabel metal1 16146 17544 16146 17544 0 _0324_
rlabel metal1 15042 16422 15042 16422 0 _0325_
rlabel metal1 15042 10982 15042 10982 0 _0326_
rlabel metal2 12834 23290 12834 23290 0 _0327_
rlabel metal1 13754 11866 13754 11866 0 _0328_
rlabel viali 12742 22066 12742 22066 0 _0329_
rlabel metal1 15410 12818 15410 12818 0 _0330_
rlabel metal1 21068 13294 21068 13294 0 _0331_
rlabel metal2 14582 10880 14582 10880 0 _0332_
rlabel metal1 19550 13838 19550 13838 0 _0333_
rlabel metal1 16100 11322 16100 11322 0 _0334_
rlabel metal1 7084 13838 7084 13838 0 _0335_
rlabel metal1 14122 13294 14122 13294 0 _0336_
rlabel metal1 12006 12614 12006 12614 0 _0337_
rlabel metal1 6900 23018 6900 23018 0 _0338_
rlabel metal1 3036 15538 3036 15538 0 _0339_
rlabel metal1 6256 16422 6256 16422 0 _0340_
rlabel metal2 4692 21556 4692 21556 0 _0341_
rlabel metal1 15318 23800 15318 23800 0 _0342_
rlabel metal1 9982 22202 9982 22202 0 _0343_
rlabel metal1 14398 23494 14398 23494 0 _0344_
rlabel metal1 13294 18666 13294 18666 0 _0345_
rlabel metal1 23690 21624 23690 21624 0 _0346_
rlabel metal2 21390 16796 21390 16796 0 _0347_
rlabel metal2 22310 19992 22310 19992 0 _0348_
rlabel metal2 21298 18836 21298 18836 0 _0349_
rlabel metal2 13202 23800 13202 23800 0 _0350_
rlabel metal1 12558 20264 12558 20264 0 _0351_
rlabel metal1 13294 21590 13294 21590 0 _0352_
rlabel metal2 6670 18020 6670 18020 0 _0353_
rlabel metal1 21298 10778 21298 10778 0 _0354_
rlabel metal1 15870 9350 15870 9350 0 _0355_
rlabel metal1 19550 10778 19550 10778 0 _0356_
rlabel metal1 10212 8058 10212 8058 0 _0357_
rlabel metal1 24656 16218 24656 16218 0 _0358_
rlabel metal1 24288 22066 24288 22066 0 _0359_
rlabel metal1 24058 16014 24058 16014 0 _0360_
rlabel metal1 24656 21590 24656 21590 0 _0361_
rlabel metal2 14490 25908 14490 25908 0 _0362_
rlabel metal1 14536 24242 14536 24242 0 _0363_
rlabel metal1 14122 24786 14122 24786 0 _0364_
rlabel metal1 9568 24718 9568 24718 0 _0365_
rlabel metal2 12282 23086 12282 23086 0 _0366_
rlabel metal1 14490 17748 14490 17748 0 _0367_
rlabel metal2 12926 21114 12926 21114 0 _0368_
rlabel metal1 15594 17782 15594 17782 0 _0369_
rlabel metal1 19504 16150 19504 16150 0 _0370_
rlabel metal1 18446 22610 18446 22610 0 _0371_
rlabel metal1 18492 15130 18492 15130 0 _0372_
rlabel metal1 18492 23154 18492 23154 0 _0373_
rlabel metal1 8050 11118 8050 11118 0 _0374_
rlabel metal1 8280 10234 8280 10234 0 _0375_
rlabel metal1 7820 12750 7820 12750 0 _0376_
rlabel metal1 11132 8602 11132 8602 0 _0377_
rlabel metal2 38318 6239 38318 6239 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 38318 33439 38318 33439 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal1 22770 37230 22770 37230 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 36984 36754 36984 36754 0 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1234 12308 1234 12308 0 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 34822 1588 34822 1588 0 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 1740 36788 1740 36788 0 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 38180 36142 38180 36142 0 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal2 29026 1588 29026 1588 0 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 2660 7548 2660 7548 0 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal3 1234 30668 1234 30668 0 ccff_head
rlabel metal2 10350 1520 10350 1520 0 ccff_tail
rlabel metal3 1924 38148 1924 38148 0 chanx_left_in[0]
rlabel metal2 4554 1554 4554 1554 0 chanx_left_in[10]
rlabel metal3 1234 20468 1234 20468 0 chanx_left_in[11]
rlabel metal1 2530 23018 2530 23018 0 chanx_left_in[12]
rlabel metal2 38318 28883 38318 28883 0 chanx_left_in[13]
rlabel metal1 18216 37230 18216 37230 0 chanx_left_in[14]
rlabel metal2 33534 1588 33534 1588 0 chanx_left_in[15]
rlabel metal3 1234 25228 1234 25228 0 chanx_left_in[16]
rlabel metal3 1234 32028 1234 32028 0 chanx_left_in[17]
rlabel metal3 1234 27268 1234 27268 0 chanx_left_in[18]
rlabel metal2 22586 1588 22586 1588 0 chanx_left_in[1]
rlabel metal2 14858 1588 14858 1588 0 chanx_left_in[2]
rlabel metal2 39330 1860 39330 1860 0 chanx_left_in[3]
rlabel metal3 2384 1428 2384 1428 0 chanx_left_in[4]
rlabel metal2 38318 20689 38318 20689 0 chanx_left_in[5]
rlabel metal1 24656 37230 24656 37230 0 chanx_left_in[6]
rlabel metal1 14030 37230 14030 37230 0 chanx_left_in[7]
rlabel metal2 36938 37009 36938 37009 0 chanx_left_in[8]
rlabel metal2 16790 1588 16790 1588 0 chanx_left_in[9]
rlabel metal3 1234 15708 1234 15708 0 chanx_left_out[0]
rlabel metal2 38226 34833 38226 34833 0 chanx_left_out[10]
rlabel metal1 15640 37094 15640 37094 0 chanx_left_out[11]
rlabel metal2 38226 8857 38226 8857 0 chanx_left_out[12]
rlabel metal2 38226 12461 38226 12461 0 chanx_left_out[13]
rlabel metal1 16928 37094 16928 37094 0 chanx_left_out[14]
rlabel metal1 10488 37094 10488 37094 0 chanx_left_out[15]
rlabel metal2 25806 1520 25806 1520 0 chanx_left_out[16]
rlabel metal2 9062 1520 9062 1520 0 chanx_left_out[17]
rlabel via2 38226 30005 38226 30005 0 chanx_left_out[18]
rlabel metal2 38042 1520 38042 1520 0 chanx_left_out[1]
rlabel metal2 38226 15793 38226 15793 0 chanx_left_out[2]
rlabel metal1 29486 37094 29486 37094 0 chanx_left_out[3]
rlabel metal1 12512 37094 12512 37094 0 chanx_left_out[4]
rlabel metal2 38226 2125 38226 2125 0 chanx_left_out[5]
rlabel metal2 38226 32113 38226 32113 0 chanx_left_out[6]
rlabel metal1 37260 37094 37260 37094 0 chanx_left_out[7]
rlabel metal1 21758 37094 21758 37094 0 chanx_left_out[8]
rlabel metal2 1794 18751 1794 18751 0 chanx_left_out[9]
rlabel metal2 38318 7701 38318 7701 0 chany_bottom_in[0]
rlabel metal3 1234 22508 1234 22508 0 chany_bottom_in[10]
rlabel metal2 4002 2941 4002 2941 0 chany_bottom_in[11]
rlabel metal1 25944 37230 25944 37230 0 chany_bottom_in[12]
rlabel metal3 1234 28628 1234 28628 0 chany_bottom_in[13]
rlabel metal2 30314 1588 30314 1588 0 chany_bottom_in[14]
rlabel metal1 33672 37230 33672 37230 0 chany_bottom_in[15]
rlabel metal1 1794 4080 1794 4080 0 chany_bottom_in[16]
rlabel metal2 2622 2166 2622 2166 0 chany_bottom_in[17]
rlabel metal2 11638 1588 11638 1588 0 chany_bottom_in[18]
rlabel metal2 36110 1588 36110 1588 0 chany_bottom_in[1]
rlabel metal2 38318 17119 38318 17119 0 chany_bottom_in[2]
rlabel metal2 38318 11033 38318 11033 0 chany_bottom_in[3]
rlabel metal2 3818 4607 3818 4607 0 chany_bottom_in[4]
rlabel metal3 1234 33388 1234 33388 0 chany_bottom_in[5]
rlabel metal2 38318 3145 38318 3145 0 chany_bottom_in[6]
rlabel metal1 4738 37230 4738 37230 0 chany_bottom_in[7]
rlabel via2 38318 14365 38318 14365 0 chany_bottom_in[8]
rlabel via2 38318 25245 38318 25245 0 chany_bottom_in[9]
rlabel metal2 31602 1520 31602 1520 0 chany_bottom_out[0]
rlabel via2 38226 27285 38226 27285 0 chany_bottom_out[10]
rlabel metal1 6302 37094 6302 37094 0 chany_bottom_out[11]
rlabel metal3 1234 23868 1234 23868 0 chany_bottom_out[12]
rlabel metal2 19366 1520 19366 1520 0 chany_bottom_out[13]
rlabel metal2 46 1792 46 1792 0 chany_bottom_out[14]
rlabel metal2 23874 1520 23874 1520 0 chany_bottom_out[15]
rlabel metal1 7912 37094 7912 37094 0 chany_bottom_out[16]
rlabel metal1 20148 37094 20148 37094 0 chany_bottom_out[17]
rlabel metal3 1234 4828 1234 4828 0 chany_bottom_out[18]
rlabel metal1 920 36890 920 36890 0 chany_bottom_out[1]
rlabel metal2 5842 1520 5842 1520 0 chany_bottom_out[2]
rlabel metal2 1334 1520 1334 1520 0 chany_bottom_out[3]
rlabel metal1 34960 37094 34960 37094 0 chany_bottom_out[4]
rlabel metal1 27876 37094 27876 37094 0 chany_bottom_out[5]
rlabel metal2 18078 1520 18078 1520 0 chany_bottom_out[6]
rlabel metal1 38778 36890 38778 36890 0 chany_bottom_out[7]
rlabel metal2 38226 4301 38226 4301 0 chany_bottom_out[8]
rlabel metal1 1564 37094 1564 37094 0 chany_bottom_out[9]
rlabel metal2 38318 21913 38318 21913 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 7130 1588 7130 1588 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 13570 1588 13570 1588 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1886 6766 1886 6766 0 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 38318 24021 38318 24021 0 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 21298 1588 21298 1588 0 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 32384 37230 32384 37230 0 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 30544 37230 30544 37230 0 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 3726 37230 3726 37230 0 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 9200 37230 9200 37230 0 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal3 2047 8228 2047 8228 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 4094 7514 4094 7514 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal2 2714 21726 2714 21726 0 mem_bottom_track_11.DFFR_0_.D
rlabel metal1 20056 21522 20056 21522 0 mem_bottom_track_11.DFFR_0_.Q
rlabel metal2 22218 22814 22218 22814 0 mem_bottom_track_11.DFFR_1_.Q
rlabel metal1 13202 15470 13202 15470 0 mem_bottom_track_13.DFFR_0_.Q
rlabel metal1 13938 11730 13938 11730 0 mem_bottom_track_13.DFFR_1_.Q
rlabel metal1 23414 24786 23414 24786 0 mem_bottom_track_15.DFFR_0_.Q
rlabel metal2 22126 20128 22126 20128 0 mem_bottom_track_15.DFFR_1_.Q
rlabel metal1 2070 9010 2070 9010 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 22862 11764 22862 11764 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal1 7038 21590 7038 21590 0 mem_bottom_track_19.DFFR_0_.Q
rlabel metal1 8004 21522 8004 21522 0 mem_bottom_track_19.DFFR_1_.Q
rlabel metal1 9522 17068 9522 17068 0 mem_bottom_track_21.DFFR_0_.Q
rlabel metal1 8372 16966 8372 16966 0 mem_bottom_track_21.DFFR_1_.Q
rlabel metal2 5750 16286 5750 16286 0 mem_bottom_track_23.DFFR_0_.Q
rlabel metal2 2714 14620 2714 14620 0 mem_bottom_track_23.DFFR_1_.Q
rlabel metal1 14398 16558 14398 16558 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal2 10534 17850 10534 17850 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal2 11408 19924 11408 19924 0 mem_bottom_track_27.DFFR_0_.Q
rlabel metal1 8648 14246 8648 14246 0 mem_bottom_track_27.DFFR_1_.Q
rlabel metal2 20654 11628 20654 11628 0 mem_bottom_track_29.DFFR_0_.Q
rlabel metal2 14490 8262 14490 8262 0 mem_bottom_track_29.DFFR_1_.Q
rlabel metal1 6256 12682 6256 12682 0 mem_bottom_track_3.DFFR_0_.Q
rlabel metal1 5842 14790 5842 14790 0 mem_bottom_track_3.DFFR_1_.Q
rlabel metal1 10028 13702 10028 13702 0 mem_bottom_track_31.DFFR_0_.Q
rlabel metal2 14674 10404 14674 10404 0 mem_bottom_track_31.DFFR_1_.Q
rlabel metal2 2622 20128 2622 20128 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 4508 16422 4508 16422 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal1 8740 17170 8740 17170 0 mem_bottom_track_35.DFFR_0_.Q
rlabel metal1 13386 23732 13386 23732 0 mem_bottom_track_35.DFFR_1_.Q
rlabel metal1 15916 20910 15916 20910 0 mem_bottom_track_37.DFFR_0_.Q
rlabel metal1 7130 21998 7130 21998 0 mem_bottom_track_37.DFFR_1_.Q
rlabel metal2 17986 9826 17986 9826 0 mem_bottom_track_5.DFFR_0_.Q
rlabel metal1 14306 8908 14306 8908 0 mem_bottom_track_5.DFFR_1_.Q
rlabel metal1 12466 6698 12466 6698 0 mem_bottom_track_7.DFFR_0_.Q
rlabel metal1 13478 7888 13478 7888 0 mem_bottom_track_7.DFFR_1_.Q
rlabel metal2 24794 23205 24794 23205 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal2 13386 8636 13386 8636 0 mem_left_track_1.DFFR_0_.Q
rlabel metal1 13018 9520 13018 9520 0 mem_left_track_1.DFFR_1_.Q
rlabel metal2 20746 20944 20746 20944 0 mem_left_track_11.DFFR_0_.D
rlabel metal2 13386 15266 13386 15266 0 mem_left_track_11.DFFR_0_.Q
rlabel metal3 5934 12988 5934 12988 0 mem_left_track_11.DFFR_1_.Q
rlabel metal2 16882 26078 16882 26078 0 mem_left_track_13.DFFR_0_.Q
rlabel metal1 1886 20536 1886 20536 0 mem_left_track_13.DFFR_1_.Q
rlabel metal1 22356 20434 22356 20434 0 mem_left_track_15.DFFR_0_.Q
rlabel metal1 23460 18258 23460 18258 0 mem_left_track_15.DFFR_1_.Q
rlabel metal1 13110 19312 13110 19312 0 mem_left_track_17.DFFR_0_.Q
rlabel metal2 15410 22916 15410 22916 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 13570 13345 13570 13345 0 mem_left_track_19.DFFR_0_.Q
rlabel metal1 8648 13226 8648 13226 0 mem_left_track_19.DFFR_1_.Q
rlabel metal1 21160 17646 21160 17646 0 mem_left_track_21.DFFR_0_.Q
rlabel metal2 22770 19822 22770 19822 0 mem_left_track_21.DFFR_1_.Q
rlabel metal1 11040 19278 11040 19278 0 mem_left_track_23.DFFR_0_.Q
rlabel metal1 12926 24140 12926 24140 0 mem_left_track_23.DFFR_1_.Q
rlabel metal2 13294 8772 13294 8772 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 18814 10642 18814 10642 0 mem_left_track_25.DFFR_1_.Q
rlabel metal1 24656 21522 24656 21522 0 mem_left_track_27.DFFR_0_.Q
rlabel metal1 24196 17170 24196 17170 0 mem_left_track_27.DFFR_1_.Q
rlabel metal1 9752 17238 9752 17238 0 mem_left_track_29.DFFR_0_.Q
rlabel metal1 12742 26350 12742 26350 0 mem_left_track_29.DFFR_1_.Q
rlabel metal1 2530 8568 2530 8568 0 mem_left_track_3.DFFR_0_.Q
rlabel metal2 25438 10404 25438 10404 0 mem_left_track_3.DFFR_1_.Q
rlabel metal1 10895 22202 10895 22202 0 mem_left_track_31.DFFR_0_.Q
rlabel metal2 10994 20638 10994 20638 0 mem_left_track_31.DFFR_1_.Q
rlabel metal1 12650 19278 12650 19278 0 mem_left_track_33.DFFR_0_.Q
rlabel metal1 22218 16014 22218 16014 0 mem_left_track_33.DFFR_1_.Q
rlabel metal1 10534 13158 10534 13158 0 mem_left_track_35.DFFR_0_.Q
rlabel metal2 10534 9724 10534 9724 0 mem_left_track_35.DFFR_1_.Q
rlabel metal2 15088 13124 15088 13124 0 mem_left_track_37.DFFR_0_.Q
rlabel metal1 25346 13294 25346 13294 0 mem_left_track_5.DFFR_0_.Q
rlabel metal1 25438 13736 25438 13736 0 mem_left_track_5.DFFR_1_.Q
rlabel metal1 24518 17646 24518 17646 0 mem_left_track_7.DFFR_0_.Q
rlabel metal1 25254 18768 25254 18768 0 mem_left_track_7.DFFR_1_.Q
rlabel metal1 24380 18734 24380 18734 0 mem_left_track_9.DFFR_0_.Q
rlabel metal1 18676 31858 18676 31858 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal2 30038 24480 30038 24480 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 21022 12818 21022 12818 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 18952 18054 18952 18054 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20838 14314 20838 14314 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 22218 14416 22218 14416 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 28198 3740 28198 3740 0 mux_bottom_track_1.out
rlabel metal2 29854 26928 29854 26928 0 mux_bottom_track_11.INVTX1_0_.out
rlabel metal1 22770 9146 22770 9146 0 mux_bottom_track_11.INVTX1_1_.out
rlabel metal1 21666 33830 21666 33830 0 mux_bottom_track_11.INVTX1_2_.out
rlabel metal2 20930 20128 20930 20128 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 20838 24480 20838 24480 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23184 35666 23184 35666 0 mux_bottom_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 25024 35802 25024 35802 0 mux_bottom_track_11.out
rlabel metal1 18124 18734 18124 18734 0 mux_bottom_track_13.INVTX1_1_.out
rlabel metal1 14766 33830 14766 33830 0 mux_bottom_track_13.INVTX1_2_.out
rlabel metal2 15226 17374 15226 17374 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 14858 19074 14858 19074 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15594 17102 15594 17102 0 mux_bottom_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 17894 6426 17894 6426 0 mux_bottom_track_13.out
rlabel metal2 19090 18972 19090 18972 0 mux_bottom_track_15.INVTX1_1_.out
rlabel metal1 22586 24140 22586 24140 0 mux_bottom_track_15.INVTX1_2_.out
rlabel metal2 19182 18462 19182 18462 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23276 23834 23276 23834 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23046 23018 23046 23018 0 mux_bottom_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 36202 36550 36202 36550 0 mux_bottom_track_15.out
rlabel metal2 25622 21216 25622 21216 0 mux_bottom_track_17.INVTX1_1_.out
rlabel metal1 18354 6426 18354 6426 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal2 20286 15776 20286 15776 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 19366 13430 19366 13430 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33810 10710 33810 10710 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 36386 8908 36386 8908 0 mux_bottom_track_17.out
rlabel metal3 11799 15300 11799 15300 0 mux_bottom_track_19.INVTX1_2_.out
rlabel metal1 15640 21318 15640 21318 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 11500 15878 11500 15878 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 8326 20077 8326 20077 0 mux_bottom_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6624 36754 6624 36754 0 mux_bottom_track_19.out
rlabel metal1 10718 17782 10718 17782 0 mux_bottom_track_21.INVTX1_1_.out
rlabel metal1 14398 19686 14398 19686 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 35558 22814 35558 22814 0 mux_bottom_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 36938 25330 36938 25330 0 mux_bottom_track_21.out
rlabel metal1 12512 17646 12512 17646 0 mux_bottom_track_23.INVTX1_0_.out
rlabel metal2 4922 23358 4922 23358 0 mux_bottom_track_23.INVTX1_1_.out
rlabel metal2 6624 22644 6624 22644 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 6900 19210 6900 19210 0 mux_bottom_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 5796 34578 5796 34578 0 mux_bottom_track_23.out
rlabel metal2 25346 12920 25346 12920 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal2 33442 20638 33442 20638 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal2 18170 17476 18170 17476 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 2346 21165 2346 21165 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 1978 23868 1978 23868 0 mux_bottom_track_25.out
rlabel metal1 12650 21862 12650 21862 0 mux_bottom_track_27.INVTX1_0_.out
rlabel metal1 15226 34102 15226 34102 0 mux_bottom_track_27.INVTX1_1_.out
rlabel metal1 13616 21862 13616 21862 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16606 15402 16606 15402 0 mux_bottom_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 18538 7786 18538 7786 0 mux_bottom_track_27.out
rlabel metal2 28014 10744 28014 10744 0 mux_bottom_track_29.INVTX1_1_.out
rlabel metal2 21390 14382 21390 14382 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 14628 12682 14628 12682 0 mux_bottom_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 4416 2414 4416 2414 0 mux_bottom_track_29.out
rlabel metal2 13386 12959 13386 12959 0 mux_bottom_track_3.INVTX1_2_.out
rlabel metal2 13110 17884 13110 17884 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 11914 13294 11914 13294 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8234 16456 8234 16456 0 mux_bottom_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 4002 36550 4002 36550 0 mux_bottom_track_3.out
rlabel metal1 6670 13838 6670 13838 0 mux_bottom_track_31.INVTX1_1_.out
rlabel metal2 12650 15011 12650 15011 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16836 13226 16836 13226 0 mux_bottom_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21206 7004 21206 7004 0 mux_bottom_track_31.out
rlabel metal1 4600 27846 4600 27846 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal2 6302 16082 6302 16082 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 6946 31790 6946 31790 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 6578 33286 6578 33286 0 mux_bottom_track_33.out
rlabel metal1 9844 22610 9844 22610 0 mux_bottom_track_35.INVTX1_1_.out
rlabel metal1 13846 18938 13846 18938 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 15594 21998 15594 21998 0 mux_bottom_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 17434 29818 17434 29818 0 mux_bottom_track_35.out
rlabel via3 5773 31756 5773 31756 0 mux_bottom_track_37.INVTX1_2_.out
rlabel metal1 16146 19958 16146 19958 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9936 22950 9936 22950 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8188 18122 8188 18122 0 mux_bottom_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6762 5236 6762 5236 0 mux_bottom_track_37.out
rlabel metal2 18446 8398 18446 8398 0 mux_bottom_track_5.INVTX1_2_.out
rlabel metal1 12650 12750 12650 12750 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 18538 11543 18538 11543 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 13386 12682 13386 12682 0 mux_bottom_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 10074 4318 10074 4318 0 mux_bottom_track_5.out
rlabel metal1 9982 6834 9982 6834 0 mux_bottom_track_7.INVTX1_2_.out
rlabel metal1 13386 14484 13386 14484 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 12282 10948 12282 10948 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12972 10506 12972 10506 0 mux_bottom_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 5474 2448 5474 2448 0 mux_bottom_track_7.out
rlabel metal2 24426 22372 24426 22372 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal2 22126 22780 22126 22780 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 25070 22848 25070 22848 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23276 22474 23276 22474 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 29854 36550 29854 36550 0 mux_bottom_track_9.out
rlabel metal1 10994 5882 10994 5882 0 mux_left_track_1.INVTX1_0_.out
rlabel metal1 14536 13362 14536 13362 0 mux_left_track_1.INVTX1_1_.out
rlabel metal1 21528 14450 21528 14450 0 mux_left_track_1.INVTX1_2_.out
rlabel metal1 11592 13838 11592 13838 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 11730 14790 11730 14790 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 11086 13974 11086 13974 0 mux_left_track_1.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 2622 23120 2622 23120 0 mux_left_track_1.out
rlabel metal1 12972 14382 12972 14382 0 mux_left_track_11.INVTX1_0_.out
rlabel metal1 17388 19346 17388 19346 0 mux_left_track_11.INVTX1_1_.out
rlabel metal2 16882 18428 16882 18428 0 mux_left_track_11.INVTX1_2_.out
rlabel metal2 17342 17102 17342 17102 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18216 17510 18216 17510 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 28566 10676 28566 10676 0 mux_left_track_11.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31418 10506 31418 10506 0 mux_left_track_11.out
rlabel metal1 9292 25330 9292 25330 0 mux_left_track_13.INVTX1_0_.out
rlabel metal1 19320 20366 19320 20366 0 mux_left_track_13.INVTX1_2_.out
rlabel metal1 13294 25126 13294 25126 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 16790 24718 16790 24718 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 32798 26588 32798 26588 0 mux_left_track_13.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 33350 28730 33350 28730 0 mux_left_track_13.out
rlabel metal2 22310 15164 22310 15164 0 mux_left_track_15.INVTX1_0_.out
rlabel metal2 23322 21012 23322 21012 0 mux_left_track_15.INVTX1_2_.out
rlabel metal1 23414 19278 23414 19278 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22954 19720 22954 19720 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 23966 19040 23966 19040 0 mux_left_track_15.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32476 36754 32476 36754 0 mux_left_track_15.out
rlabel metal1 10580 33830 10580 33830 0 mux_left_track_17.INVTX1_0_.out
rlabel metal1 14214 14926 14214 14926 0 mux_left_track_17.INVTX1_2_.out
rlabel metal1 13616 23222 13616 23222 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15502 19788 15502 19788 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 15594 21223 15594 21223 0 mux_left_track_17.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 18262 34510 18262 34510 0 mux_left_track_17.out
rlabel metal1 31878 14450 31878 14450 0 mux_left_track_19.INVTX1_0_.out
rlabel metal1 14536 14042 14536 14042 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 15502 15742 15502 15742 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8970 15674 8970 15674 0 mux_left_track_19.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6348 15878 6348 15878 0 mux_left_track_19.out
rlabel metal1 23690 19448 23690 19448 0 mux_left_track_21.INVTX1_0_.out
rlabel metal1 21528 19414 21528 19414 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 23552 19890 23552 19890 0 mux_left_track_21.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 29578 27098 29578 27098 0 mux_left_track_21.out
rlabel metal2 6440 21420 6440 21420 0 mux_left_track_23.INVTX1_0_.out
rlabel metal2 25714 14960 25714 14960 0 mux_left_track_23.INVTX1_1_.out
rlabel metal1 14306 19414 14306 19414 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 13938 23154 13938 23154 0 mux_left_track_23.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15272 34578 15272 34578 0 mux_left_track_23.out
rlabel metal1 8372 6630 8372 6630 0 mux_left_track_25.INVTX1_0_.out
rlabel metal1 22816 14450 22816 14450 0 mux_left_track_25.INVTX1_1_.out
rlabel metal1 18308 11050 18308 11050 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 28382 10540 28382 10540 0 mux_left_track_25.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33120 9554 33120 9554 0 mux_left_track_25.out
rlabel metal1 24380 21862 24380 21862 0 mux_left_track_27.INVTX1_0_.out
rlabel metal1 24748 20434 24748 20434 0 mux_left_track_27.INVTX1_1_.out
rlabel metal1 23322 21862 23322 21862 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 24656 16422 24656 16422 0 mux_left_track_27.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35558 15028 35558 15028 0 mux_left_track_27.out
rlabel metal2 8878 25772 8878 25772 0 mux_left_track_29.INVTX1_0_.out
rlabel metal2 13754 24548 13754 24548 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 14766 27540 14766 27540 0 mux_left_track_29.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 15272 35054 15272 35054 0 mux_left_track_29.out
rlabel metal1 22402 12308 22402 12308 0 mux_left_track_3.INVTX1_0_.out
rlabel metal2 23138 13566 23138 13566 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 22954 15232 22954 15232 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 23966 12988 23966 12988 0 mux_left_track_3.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31740 5202 31740 5202 0 mux_left_track_3.out
rlabel metal2 25438 7327 25438 7327 0 mux_left_track_31.INVTX1_0_.out
rlabel metal1 14214 17510 14214 17510 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12512 31790 12512 31790 0 mux_left_track_31.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 12006 31994 12006 31994 0 mux_left_track_31.out
rlabel metal2 28106 28526 28106 28526 0 mux_left_track_33.INVTX1_0_.out
rlabel metal2 18630 22848 18630 22848 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20884 16150 20884 16150 0 mux_left_track_33.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 23230 10438 23230 10438 0 mux_left_track_33.out
rlabel metal1 6164 10574 6164 10574 0 mux_left_track_35.INVTX1_0_.out
rlabel metal1 9522 12342 9522 12342 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 9016 12614 9016 12614 0 mux_left_track_35.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 9614 5270 9614 5270 0 mux_left_track_35.out
rlabel metal1 9752 5814 9752 5814 0 mux_left_track_37.INVTX1_0_.out
rlabel metal2 14766 13702 14766 13702 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 16882 15368 16882 15368 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 24886 14416 24886 14416 0 mux_left_track_37.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 29854 21114 29854 21114 0 mux_left_track_37.out
rlabel metal2 24702 9996 24702 9996 0 mux_left_track_5.INVTX1_0_.out
rlabel metal2 25346 14484 25346 14484 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 23874 14144 23874 14144 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25484 14790 25484 14790 0 mux_left_track_5.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 31832 14586 31832 14586 0 mux_left_track_5.out
rlabel metal1 23322 17068 23322 17068 0 mux_left_track_7.INVTX1_0_.out
rlabel metal1 23460 16966 23460 16966 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 25438 20672 25438 20672 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 25024 19958 25024 19958 0 mux_left_track_7.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 27278 31926 27278 31926 0 mux_left_track_7.out
rlabel metal1 23046 18190 23046 18190 0 mux_left_track_9.INVTX1_0_.out
rlabel metal2 24058 20536 24058 20536 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 18538 21862 18538 21862 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 18308 21930 18308 21930 0 mux_left_track_9.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 14812 34578 14812 34578 0 mux_left_track_9.out
rlabel metal2 38134 9316 38134 9316 0 net1
rlabel metal1 4554 4114 4554 4114 0 net10
rlabel metal2 20102 14484 20102 14484 0 net100
rlabel metal1 11362 17102 11362 17102 0 net101
rlabel metal2 18170 11424 18170 11424 0 net102
rlabel metal1 8050 10030 8050 10030 0 net103
rlabel metal1 24518 23154 24518 23154 0 net104
rlabel metal2 20378 24956 20378 24956 0 net105
rlabel metal1 14582 21590 14582 21590 0 net106
rlabel metal2 22678 24208 22678 24208 0 net107
rlabel metal1 19412 13294 19412 13294 0 net108
rlabel metal2 9614 15402 9614 15402 0 net109
rlabel metal1 1564 30566 1564 30566 0 net11
rlabel metal2 9430 22916 9430 22916 0 net110
rlabel metal1 11224 14926 11224 14926 0 net111
rlabel metal1 22862 14994 22862 14994 0 net112
rlabel metal2 24610 13634 24610 13634 0 net113
rlabel metal1 25990 20978 25990 20978 0 net114
rlabel metal1 18906 22066 18906 22066 0 net115
rlabel metal2 17710 18020 17710 18020 0 net116
rlabel metal2 15962 25568 15962 25568 0 net117
rlabel metal1 22356 18802 22356 18802 0 net118
rlabel metal1 13984 17714 13984 17714 0 net119
rlabel metal1 4324 37162 4324 37162 0 net12
rlabel metal1 16882 16116 16882 16116 0 net120
rlabel metal1 16744 12954 16744 12954 0 net121
rlabel metal1 17342 20570 17342 20570 0 net122
rlabel metal2 5198 15776 5198 15776 0 net123
rlabel metal1 11730 18190 11730 18190 0 net124
rlabel metal1 15088 12886 15088 12886 0 net125
rlabel metal1 14444 12750 14444 12750 0 net126
rlabel metal1 16606 13158 16606 13158 0 net127
rlabel metal2 6762 23596 6762 23596 0 net128
rlabel metal1 16054 23630 16054 23630 0 net129
rlabel metal1 5060 2618 5060 2618 0 net13
rlabel metal1 23644 21454 23644 21454 0 net130
rlabel metal2 13110 23392 13110 23392 0 net131
rlabel metal1 21850 11220 21850 11220 0 net132
rlabel metal2 24610 16864 24610 16864 0 net133
rlabel metal1 13938 25330 13938 25330 0 net134
rlabel metal1 11408 22678 11408 22678 0 net135
rlabel metal1 19504 14450 19504 14450 0 net136
rlabel metal1 7774 11186 7774 11186 0 net137
rlabel metal2 1978 19482 1978 19482 0 net14
rlabel metal2 3910 23460 3910 23460 0 net15
rlabel metal2 33350 26894 33350 26894 0 net16
rlabel metal1 18170 37128 18170 37128 0 net17
rlabel metal1 30774 7854 30774 7854 0 net18
rlabel metal1 5796 21522 5796 21522 0 net19
rlabel metal2 38134 30668 38134 30668 0 net2
rlabel metal1 2806 32198 2806 32198 0 net20
rlabel metal2 5750 25500 5750 25500 0 net21
rlabel metal2 22678 4454 22678 4454 0 net22
rlabel metal1 14398 6290 14398 6290 0 net23
rlabel metal2 35650 4726 35650 4726 0 net24
rlabel metal1 6624 3706 6624 3706 0 net25
rlabel metal2 38134 21318 38134 21318 0 net26
rlabel metal1 23828 37094 23828 37094 0 net27
rlabel metal2 14306 35530 14306 35530 0 net28
rlabel metal1 36317 37094 36317 37094 0 net29
rlabel metal1 21850 37162 21850 37162 0 net3
rlabel metal1 17618 2618 17618 2618 0 net30
rlabel metal1 37674 8058 37674 8058 0 net31
rlabel metal1 6578 22678 6578 22678 0 net32
rlabel metal1 6670 3162 6670 3162 0 net33
rlabel metal1 25484 37094 25484 37094 0 net34
rlabel metal2 6578 27982 6578 27982 0 net35
rlabel metal1 28980 2550 28980 2550 0 net36
rlabel metal1 30866 37162 30866 37162 0 net37
rlabel metal1 2162 3978 2162 3978 0 net38
rlabel metal2 5750 4658 5750 4658 0 net39
rlabel metal2 36754 33422 36754 33422 0 net4
rlabel metal1 11454 2618 11454 2618 0 net40
rlabel metal1 36041 2618 36041 2618 0 net41
rlabel metal1 37007 17306 37007 17306 0 net42
rlabel metal1 37674 11322 37674 11322 0 net43
rlabel metal1 4186 2890 4186 2890 0 net44
rlabel metal1 2760 33286 2760 33286 0 net45
rlabel metal1 36064 3706 36064 3706 0 net46
rlabel metal2 4646 35530 4646 35530 0 net47
rlabel metal1 37007 14246 37007 14246 0 net48
rlabel metal2 33994 24106 33994 24106 0 net49
rlabel metal1 1886 6426 1886 6426 0 net5
rlabel metal1 37007 21862 37007 21862 0 net50
rlabel metal1 7360 2618 7360 2618 0 net51
rlabel metal1 14490 2618 14490 2618 0 net52
rlabel metal1 1610 6664 1610 6664 0 net53
rlabel metal2 37030 23324 37030 23324 0 net54
rlabel metal1 21620 8466 21620 8466 0 net55
rlabel metal1 31510 37094 31510 37094 0 net56
rlabel metal1 30268 37094 30268 37094 0 net57
rlabel metal2 4002 36992 4002 36992 0 net58
rlabel metal1 11500 36822 11500 36822 0 net59
rlabel metal1 34914 2312 34914 2312 0 net6
rlabel metal1 16560 2516 16560 2516 0 net60
rlabel metal1 10626 2414 10626 2414 0 net61
rlabel metal1 1656 17170 1656 17170 0 net62
rlabel metal1 35144 30906 35144 30906 0 net63
rlabel metal1 15456 34714 15456 34714 0 net64
rlabel metal2 38042 9146 38042 9146 0 net65
rlabel metal2 38042 13804 38042 13804 0 net66
rlabel metal2 16882 36244 16882 36244 0 net67
rlabel metal2 11638 36788 11638 36788 0 net68
rlabel metal1 25346 2414 25346 2414 0 net69
rlabel metal2 2346 36890 2346 36890 0 net7
rlabel metal1 9292 4998 9292 4998 0 net70
rlabel metal2 33626 28118 33626 28118 0 net71
rlabel metal2 36938 3706 36938 3706 0 net72
rlabel metal2 36110 15606 36110 15606 0 net73
rlabel metal1 28842 37230 28842 37230 0 net74
rlabel metal1 13524 37162 13524 37162 0 net75
rlabel metal2 37030 4828 37030 4828 0 net76
rlabel metal1 35236 29818 35236 29818 0 net77
rlabel metal2 37490 36924 37490 36924 0 net78
rlabel metal1 21344 37230 21344 37230 0 net79
rlabel metal1 37720 36006 37720 36006 0 net8
rlabel metal1 4232 10438 4232 10438 0 net80
rlabel metal1 32338 2448 32338 2448 0 net81
rlabel metal1 37398 27438 37398 27438 0 net82
rlabel metal1 6072 34714 6072 34714 0 net83
rlabel metal1 1702 23834 1702 23834 0 net84
rlabel metal1 18906 5542 18906 5542 0 net85
rlabel metal1 3404 2618 3404 2618 0 net86
rlabel metal1 23966 2414 23966 2414 0 net87
rlabel metal1 7360 34714 7360 34714 0 net88
rlabel metal1 19320 37230 19320 37230 0 net89
rlabel metal1 29210 2618 29210 2618 0 net9
rlabel metal1 1610 5168 1610 5168 0 net90
rlabel metal1 2576 36754 2576 36754 0 net91
rlabel metal1 6808 2414 6808 2414 0 net92
rlabel metal1 1610 2448 1610 2448 0 net93
rlabel metal1 33212 36890 33212 36890 0 net94
rlabel metal2 27830 37060 27830 37060 0 net95
rlabel metal1 17940 5542 17940 5542 0 net96
rlabel metal1 38042 36788 38042 36788 0 net97
rlabel metal1 37122 7174 37122 7174 0 net98
rlabel metal1 3174 36618 3174 36618 0 net99
rlabel metal2 27094 1554 27094 1554 0 pReset
rlabel metal2 1610 20094 1610 20094 0 prog_clk
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
