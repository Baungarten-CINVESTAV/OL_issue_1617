magic
tech sky130A
magscale 1 2
timestamp 1674219698
<< viali >>
rect 2145 37417 2179 37451
rect 17049 37417 17083 37451
rect 33241 37417 33275 37451
rect 6837 37349 6871 37383
rect 10333 37281 10367 37315
rect 14933 37281 14967 37315
rect 20637 37281 20671 37315
rect 22661 37281 22695 37315
rect 30941 37281 30975 37315
rect 34897 37281 34931 37315
rect 2053 37213 2087 37247
rect 2697 37213 2731 37247
rect 4169 37213 4203 37247
rect 4629 37213 4663 37247
rect 6653 37213 6687 37247
rect 7481 37213 7515 37247
rect 9137 37213 9171 37247
rect 10609 37213 10643 37247
rect 11713 37213 11747 37247
rect 13001 37213 13035 37247
rect 14473 37213 14507 37247
rect 15209 37213 15243 37247
rect 18337 37213 18371 37247
rect 19901 37213 19935 37247
rect 20913 37213 20947 37247
rect 22937 37213 22971 37247
rect 24593 37213 24627 37247
rect 25329 37213 25363 37247
rect 27169 37213 27203 37247
rect 27905 37213 27939 37247
rect 28825 37213 28859 37247
rect 29745 37213 29779 37247
rect 31217 37213 31251 37247
rect 32321 37213 32355 37247
rect 33057 37213 33091 37247
rect 33793 37213 33827 37247
rect 35173 37213 35207 37247
rect 36185 37213 36219 37247
rect 37565 37213 37599 37247
rect 16957 37145 16991 37179
rect 2881 37077 2915 37111
rect 3985 37077 4019 37111
rect 4813 37077 4847 37111
rect 7297 37077 7331 37111
rect 9321 37077 9355 37111
rect 11897 37077 11931 37111
rect 13185 37077 13219 37111
rect 14289 37077 14323 37111
rect 18153 37077 18187 37111
rect 20085 37077 20119 37111
rect 24777 37077 24811 37111
rect 25513 37077 25547 37111
rect 27353 37077 27387 37111
rect 28089 37077 28123 37111
rect 28641 37077 28675 37111
rect 29929 37077 29963 37111
rect 32505 37077 32539 37111
rect 33977 37077 34011 37111
rect 36369 37077 36403 37111
rect 37657 37077 37691 37111
rect 1777 36873 1811 36907
rect 3249 36873 3283 36907
rect 11897 36873 11931 36907
rect 19625 36873 19659 36907
rect 22201 36873 22235 36907
rect 23489 36873 23523 36907
rect 36829 36873 36863 36907
rect 3157 36805 3191 36839
rect 4077 36805 4111 36839
rect 15669 36805 15703 36839
rect 38117 36805 38151 36839
rect 1593 36737 1627 36771
rect 2421 36737 2455 36771
rect 5457 36737 5491 36771
rect 6745 36737 6779 36771
rect 9137 36737 9171 36771
rect 11713 36737 11747 36771
rect 17877 36737 17911 36771
rect 18521 36737 18555 36771
rect 19441 36737 19475 36771
rect 22017 36737 22051 36771
rect 23305 36737 23339 36771
rect 25789 36737 25823 36771
rect 28089 36737 28123 36771
rect 29285 36737 29319 36771
rect 30941 36737 30975 36771
rect 35909 36737 35943 36771
rect 36645 36737 36679 36771
rect 9413 36669 9447 36703
rect 4261 36601 4295 36635
rect 15853 36601 15887 36635
rect 17693 36601 17727 36635
rect 25605 36601 25639 36635
rect 27905 36601 27939 36635
rect 30757 36601 30791 36635
rect 36093 36601 36127 36635
rect 2513 36533 2547 36567
rect 5457 36533 5491 36567
rect 6561 36533 6595 36567
rect 18337 36533 18371 36567
rect 29101 36533 29135 36567
rect 38209 36533 38243 36567
rect 1777 36329 1811 36363
rect 5365 36329 5399 36363
rect 9137 36329 9171 36363
rect 22385 36329 22419 36363
rect 37473 36329 37507 36363
rect 1593 36125 1627 36159
rect 2513 36125 2547 36159
rect 5549 36125 5583 36159
rect 9321 36125 9355 36159
rect 22569 36125 22603 36159
rect 36369 36125 36403 36159
rect 37289 36125 37323 36159
rect 38025 36125 38059 36159
rect 2329 35989 2363 36023
rect 36185 35989 36219 36023
rect 38209 35989 38243 36023
rect 11713 35785 11747 35819
rect 11897 35649 11931 35683
rect 36921 35649 36955 35683
rect 38025 35649 38059 35683
rect 1593 35581 1627 35615
rect 1869 35581 1903 35615
rect 36737 35445 36771 35479
rect 38209 35445 38243 35479
rect 38209 35241 38243 35275
rect 10701 35037 10735 35071
rect 38025 35037 38059 35071
rect 10793 34901 10827 34935
rect 1593 34697 1627 34731
rect 27629 34697 27663 34731
rect 35449 34697 35483 34731
rect 1777 34561 1811 34595
rect 6561 34561 6595 34595
rect 10793 34561 10827 34595
rect 27813 34561 27847 34595
rect 34713 34561 34747 34595
rect 34989 34561 35023 34595
rect 35633 34561 35667 34595
rect 6653 34493 6687 34527
rect 37473 34493 37507 34527
rect 37749 34493 37783 34527
rect 10885 34357 10919 34391
rect 10885 34153 10919 34187
rect 27537 34153 27571 34187
rect 10793 33949 10827 33983
rect 22661 33949 22695 33983
rect 24593 33949 24627 33983
rect 27721 33949 27755 33983
rect 24685 33881 24719 33915
rect 22753 33813 22787 33847
rect 23489 33609 23523 33643
rect 1777 33473 1811 33507
rect 2421 33473 2455 33507
rect 23673 33473 23707 33507
rect 30389 33473 30423 33507
rect 38117 33473 38151 33507
rect 1593 33337 1627 33371
rect 30481 33337 30515 33371
rect 38301 33337 38335 33371
rect 2237 33269 2271 33303
rect 2973 33065 3007 33099
rect 2329 32997 2363 33031
rect 1593 32861 1627 32895
rect 2513 32861 2547 32895
rect 3157 32861 3191 32895
rect 6929 32861 6963 32895
rect 29745 32861 29779 32895
rect 1777 32725 1811 32759
rect 2237 32725 2271 32759
rect 7021 32725 7055 32759
rect 29837 32725 29871 32759
rect 1593 32385 1627 32419
rect 3065 32385 3099 32419
rect 3709 32385 3743 32419
rect 28549 32385 28583 32419
rect 37749 32385 37783 32419
rect 37473 32317 37507 32351
rect 1777 32181 1811 32215
rect 2881 32181 2915 32215
rect 3525 32181 3559 32215
rect 28641 32181 28675 32215
rect 2973 31977 3007 32011
rect 35541 31977 35575 32011
rect 1685 31909 1719 31943
rect 2421 31841 2455 31875
rect 4077 31841 4111 31875
rect 1869 31773 1903 31807
rect 2329 31773 2363 31807
rect 3157 31773 3191 31807
rect 3985 31773 4019 31807
rect 17969 31773 18003 31807
rect 18061 31773 18095 31807
rect 35725 31773 35759 31807
rect 37473 31773 37507 31807
rect 37749 31773 37783 31807
rect 11805 31637 11839 31671
rect 4997 31433 5031 31467
rect 20453 31433 20487 31467
rect 4077 31365 4111 31399
rect 1869 31297 1903 31331
rect 3249 31297 3283 31331
rect 3985 31297 4019 31331
rect 5181 31297 5215 31331
rect 11713 31297 11747 31331
rect 18705 31297 18739 31331
rect 19349 31297 19383 31331
rect 20637 31297 20671 31331
rect 2513 31229 2547 31263
rect 12449 31229 12483 31263
rect 18797 31161 18831 31195
rect 1961 31093 1995 31127
rect 3341 31093 3375 31127
rect 11805 31093 11839 31127
rect 19441 31093 19475 31127
rect 6561 30889 6595 30923
rect 13369 30889 13403 30923
rect 7849 30821 7883 30855
rect 2697 30753 2731 30787
rect 11713 30753 11747 30787
rect 19901 30753 19935 30787
rect 23029 30753 23063 30787
rect 2605 30685 2639 30719
rect 3433 30685 3467 30719
rect 5089 30685 5123 30719
rect 5825 30685 5859 30719
rect 6469 30685 6503 30719
rect 7757 30685 7791 30719
rect 9137 30685 9171 30719
rect 9781 30685 9815 30719
rect 10977 30685 11011 30719
rect 13277 30685 13311 30719
rect 15025 30685 15059 30719
rect 1961 30617 1995 30651
rect 9229 30617 9263 30651
rect 11805 30617 11839 30651
rect 12725 30617 12759 30651
rect 19993 30617 20027 30651
rect 20913 30617 20947 30651
rect 22753 30617 22787 30651
rect 22845 30617 22879 30651
rect 38117 30617 38151 30651
rect 2053 30549 2087 30583
rect 3249 30549 3283 30583
rect 4445 30549 4479 30583
rect 5181 30549 5215 30583
rect 5917 30549 5951 30583
rect 7113 30549 7147 30583
rect 8401 30549 8435 30583
rect 9873 30549 9907 30583
rect 11069 30549 11103 30583
rect 15117 30549 15151 30583
rect 38209 30549 38243 30583
rect 16129 30345 16163 30379
rect 8861 30277 8895 30311
rect 8953 30277 8987 30311
rect 13369 30277 13403 30311
rect 13461 30277 13495 30311
rect 15577 30277 15611 30311
rect 19625 30277 19659 30311
rect 21373 30277 21407 30311
rect 22569 30277 22603 30311
rect 1593 30209 1627 30243
rect 2697 30209 2731 30243
rect 3341 30209 3375 30243
rect 3985 30209 4019 30243
rect 5273 30209 5307 30243
rect 7205 30209 7239 30243
rect 7665 30209 7699 30243
rect 10325 30215 10359 30249
rect 10425 30209 10459 30243
rect 10977 30209 11011 30243
rect 11897 30209 11931 30243
rect 12357 30209 12391 30243
rect 14841 30209 14875 30243
rect 15485 30209 15519 30243
rect 16313 30209 16347 30243
rect 21281 30209 21315 30243
rect 22385 30209 22419 30243
rect 3433 30141 3467 30175
rect 5733 30141 5767 30175
rect 9229 30141 9263 30175
rect 12449 30141 12483 30175
rect 14381 30141 14415 30175
rect 18797 30141 18831 30175
rect 19533 30141 19567 30175
rect 19809 30141 19843 30175
rect 1777 30073 1811 30107
rect 5089 30073 5123 30107
rect 2789 30005 2823 30039
rect 4077 30005 4111 30039
rect 7021 30005 7055 30039
rect 7757 30005 7791 30039
rect 11069 30005 11103 30039
rect 11713 30005 11747 30039
rect 14933 30005 14967 30039
rect 2697 29801 2731 29835
rect 16405 29801 16439 29835
rect 22109 29801 22143 29835
rect 26157 29801 26191 29835
rect 20085 29733 20119 29767
rect 10517 29665 10551 29699
rect 11069 29665 11103 29699
rect 12449 29665 12483 29699
rect 12909 29665 12943 29699
rect 20821 29665 20855 29699
rect 1593 29597 1627 29631
rect 2605 29597 2639 29631
rect 3249 29597 3283 29631
rect 4537 29597 4571 29631
rect 5181 29597 5215 29631
rect 5825 29597 5859 29631
rect 6469 29597 6503 29631
rect 7113 29597 7147 29631
rect 7757 29597 7791 29631
rect 8401 29597 8435 29631
rect 9137 29597 9171 29631
rect 9965 29593 9999 29627
rect 14565 29597 14599 29631
rect 15669 29597 15703 29631
rect 16313 29597 16347 29631
rect 18705 29597 18739 29631
rect 20729 29597 20763 29631
rect 22017 29597 22051 29631
rect 24593 29597 24627 29631
rect 26065 29597 26099 29631
rect 26709 29597 26743 29631
rect 38301 29597 38335 29631
rect 4629 29529 4663 29563
rect 6561 29529 6595 29563
rect 10618 29529 10652 29563
rect 12541 29529 12575 29563
rect 19533 29529 19567 29563
rect 19625 29529 19659 29563
rect 1777 29461 1811 29495
rect 3341 29461 3375 29495
rect 5273 29461 5307 29495
rect 5917 29461 5951 29495
rect 7205 29461 7239 29495
rect 7849 29461 7883 29495
rect 8493 29461 8527 29495
rect 9229 29461 9263 29495
rect 9781 29461 9815 29495
rect 14657 29461 14691 29495
rect 15761 29461 15795 29495
rect 18797 29461 18831 29495
rect 23765 29461 23799 29495
rect 24685 29461 24719 29495
rect 26801 29461 26835 29495
rect 38117 29461 38151 29495
rect 8401 29257 8435 29291
rect 9505 29257 9539 29291
rect 10241 29189 10275 29223
rect 12081 29189 12115 29223
rect 12817 29189 12851 29223
rect 14749 29189 14783 29223
rect 18981 29189 19015 29223
rect 20453 29189 20487 29223
rect 20545 29189 20579 29223
rect 23581 29189 23615 29223
rect 23673 29189 23707 29223
rect 25145 29189 25179 29223
rect 25237 29189 25271 29223
rect 1869 29121 1903 29155
rect 2513 29121 2547 29155
rect 3249 29121 3283 29155
rect 3985 29121 4019 29155
rect 4629 29121 4663 29155
rect 5733 29121 5767 29155
rect 7113 29121 7147 29155
rect 8309 29121 8343 29155
rect 9413 29121 9447 29155
rect 11989 29121 12023 29155
rect 15301 29121 15335 29155
rect 15761 29121 15795 29155
rect 15853 29121 15887 29155
rect 16865 29121 16899 29155
rect 18153 29121 18187 29155
rect 1961 29053 1995 29087
rect 5825 29053 5859 29087
rect 10149 29053 10183 29087
rect 10793 29053 10827 29087
rect 12725 29053 12759 29087
rect 13645 29053 13679 29087
rect 14657 29053 14691 29087
rect 18889 29053 18923 29087
rect 19349 29053 19383 29087
rect 21097 29053 21131 29087
rect 23949 29053 23983 29087
rect 25421 29053 25455 29087
rect 37473 29053 37507 29087
rect 37749 29053 37783 29087
rect 2605 28985 2639 29019
rect 3341 28985 3375 29019
rect 4077 28985 4111 29019
rect 4721 28985 4755 29019
rect 7205 28985 7239 29019
rect 16957 28985 16991 29019
rect 18245 28917 18279 28951
rect 18797 28713 18831 28747
rect 20177 28713 20211 28747
rect 24593 28713 24627 28747
rect 26893 28713 26927 28747
rect 17601 28645 17635 28679
rect 23489 28645 23523 28679
rect 7849 28577 7883 28611
rect 25329 28577 25363 28611
rect 25605 28577 25639 28611
rect 1961 28509 1995 28543
rect 2605 28509 2639 28543
rect 3249 28509 3283 28543
rect 3985 28509 4019 28543
rect 4629 28509 4663 28543
rect 5273 28509 5307 28543
rect 6101 28509 6135 28543
rect 6837 28509 6871 28543
rect 7757 28509 7791 28543
rect 8401 28509 8435 28543
rect 9229 28509 9263 28543
rect 10241 28509 10275 28543
rect 10793 28509 10827 28543
rect 11621 28509 11655 28543
rect 16221 28509 16255 28543
rect 16865 28509 16899 28543
rect 17509 28509 17543 28543
rect 18705 28509 18739 28543
rect 19441 28509 19475 28543
rect 20361 28509 20395 28543
rect 20821 28509 20855 28543
rect 21925 28509 21959 28543
rect 23305 28509 23339 28543
rect 24777 28509 24811 28543
rect 26801 28509 26835 28543
rect 27445 28509 27479 28543
rect 31953 28509 31987 28543
rect 7021 28441 7055 28475
rect 12357 28441 12391 28475
rect 12449 28441 12483 28475
rect 13369 28441 13403 28475
rect 14381 28441 14415 28475
rect 14473 28441 14507 28475
rect 15393 28441 15427 28475
rect 25421 28441 25455 28475
rect 2053 28373 2087 28407
rect 2697 28373 2731 28407
rect 3341 28373 3375 28407
rect 4077 28373 4111 28407
rect 4721 28373 4755 28407
rect 5365 28373 5399 28407
rect 6193 28373 6227 28407
rect 8493 28373 8527 28407
rect 9321 28373 9355 28407
rect 10057 28373 10091 28407
rect 10885 28373 10919 28407
rect 11713 28373 11747 28407
rect 16313 28373 16347 28407
rect 16957 28373 16991 28407
rect 19533 28373 19567 28407
rect 20913 28373 20947 28407
rect 22017 28373 22051 28407
rect 27537 28373 27571 28407
rect 32045 28373 32079 28407
rect 3433 28169 3467 28203
rect 11989 28169 12023 28203
rect 24317 28169 24351 28203
rect 24961 28169 24995 28203
rect 5457 28101 5491 28135
rect 6009 28101 6043 28135
rect 7113 28101 7147 28135
rect 8033 28101 8067 28135
rect 13277 28101 13311 28135
rect 13369 28101 13403 28135
rect 18613 28101 18647 28135
rect 20554 28101 20588 28135
rect 22109 28101 22143 28135
rect 22201 28101 22235 28135
rect 23673 28101 23707 28135
rect 25605 28101 25639 28135
rect 25697 28101 25731 28135
rect 27261 28101 27295 28135
rect 1593 28033 1627 28067
rect 2697 28033 2731 28067
rect 3341 28033 3375 28067
rect 3985 28033 4019 28067
rect 4629 28033 4663 28067
rect 8493 28033 8527 28067
rect 9321 28033 9355 28067
rect 9965 28033 9999 28067
rect 10609 28033 10643 28067
rect 11897 28033 11931 28067
rect 12541 28033 12575 28067
rect 12633 28033 12667 28067
rect 15209 28033 15243 28067
rect 16129 28033 16163 28067
rect 16865 28033 16899 28067
rect 17509 28033 17543 28067
rect 23581 28033 23615 28067
rect 24225 28033 24259 28067
rect 24869 28033 24903 28067
rect 27169 28033 27203 28067
rect 2789 27965 2823 27999
rect 5365 27965 5399 27999
rect 7021 27965 7055 27999
rect 9413 27965 9447 27999
rect 14105 27965 14139 27999
rect 15301 27965 15335 27999
rect 18521 27965 18555 27999
rect 19533 27965 19567 27999
rect 20453 27965 20487 27999
rect 20729 27965 20763 27999
rect 23121 27965 23155 27999
rect 26617 27965 26651 27999
rect 1777 27897 1811 27931
rect 4721 27897 4755 27931
rect 10057 27897 10091 27931
rect 17601 27897 17635 27931
rect 4077 27829 4111 27863
rect 8585 27829 8619 27863
rect 10701 27829 10735 27863
rect 16221 27829 16255 27863
rect 16957 27829 16991 27863
rect 20729 27557 20763 27591
rect 8493 27489 8527 27523
rect 9597 27489 9631 27523
rect 10793 27489 10827 27523
rect 12357 27489 12391 27523
rect 13001 27489 13035 27523
rect 20177 27489 20211 27523
rect 21373 27489 21407 27523
rect 22569 27489 22603 27523
rect 23581 27489 23615 27523
rect 25697 27489 25731 27523
rect 26617 27489 26651 27523
rect 27629 27489 27663 27523
rect 37749 27489 37783 27523
rect 1593 27421 1627 27455
rect 2605 27421 2639 27455
rect 3249 27421 3283 27455
rect 4261 27421 4295 27455
rect 4905 27421 4939 27455
rect 7481 27421 7515 27455
rect 8401 27421 8435 27455
rect 12265 27421 12299 27455
rect 12909 27421 12943 27455
rect 13553 27421 13587 27455
rect 17601 27421 17635 27455
rect 18705 27421 18739 27455
rect 19441 27421 19475 27455
rect 28365 27421 28399 27455
rect 37473 27421 37507 27455
rect 5641 27353 5675 27387
rect 5733 27353 5767 27387
rect 6653 27353 6687 27387
rect 7573 27353 7607 27387
rect 9229 27353 9263 27387
rect 9321 27353 9355 27387
rect 10885 27353 10919 27387
rect 11805 27353 11839 27387
rect 14933 27353 14967 27387
rect 15025 27353 15059 27387
rect 15577 27353 15611 27387
rect 16129 27353 16163 27387
rect 16221 27353 16255 27387
rect 17141 27353 17175 27387
rect 18797 27353 18831 27387
rect 20269 27353 20303 27387
rect 21465 27353 21499 27387
rect 22017 27353 22051 27387
rect 22661 27353 22695 27387
rect 25789 27353 25823 27387
rect 27261 27353 27295 27387
rect 27353 27353 27387 27387
rect 1777 27285 1811 27319
rect 2697 27285 2731 27319
rect 3341 27285 3375 27319
rect 4353 27285 4387 27319
rect 4997 27285 5031 27319
rect 13645 27285 13679 27319
rect 17693 27285 17727 27319
rect 19533 27285 19567 27319
rect 28457 27285 28491 27319
rect 21373 27081 21407 27115
rect 25881 27081 25915 27115
rect 30757 27081 30791 27115
rect 8309 27013 8343 27047
rect 8861 27013 8895 27047
rect 9505 27013 9539 27047
rect 11897 27013 11931 27047
rect 19073 27013 19107 27047
rect 19165 27013 19199 27047
rect 22753 27013 22787 27047
rect 27721 27013 27755 27047
rect 29285 27013 29319 27047
rect 1961 26945 1995 26979
rect 2605 26945 2639 26979
rect 3249 26945 3283 26979
rect 3893 26945 3927 26979
rect 4537 26945 4571 26979
rect 5181 26945 5215 26979
rect 5825 26945 5859 26979
rect 6653 26945 6687 26979
rect 7297 26945 7331 26979
rect 10977 26945 11011 26979
rect 13553 26945 13587 26979
rect 14197 26945 14231 26979
rect 14841 26945 14875 26979
rect 15669 26945 15703 26979
rect 16865 26945 16899 26979
rect 17509 26945 17543 26979
rect 18153 26945 18187 26979
rect 20545 26945 20579 26979
rect 21281 26945 21315 26979
rect 25789 26945 25823 26979
rect 30665 26945 30699 26979
rect 38301 26945 38335 26979
rect 3985 26877 4019 26911
rect 8217 26877 8251 26911
rect 9413 26877 9447 26911
rect 9689 26877 9723 26911
rect 11805 26877 11839 26911
rect 12817 26877 12851 26911
rect 14289 26877 14323 26911
rect 20085 26877 20119 26911
rect 22661 26877 22695 26911
rect 22937 26877 22971 26911
rect 27629 26877 27663 26911
rect 28641 26877 28675 26911
rect 29193 26877 29227 26911
rect 3341 26809 3375 26843
rect 5273 26809 5307 26843
rect 6745 26809 6779 26843
rect 29745 26809 29779 26843
rect 38117 26809 38151 26843
rect 2053 26741 2087 26775
rect 2697 26741 2731 26775
rect 4629 26741 4663 26775
rect 5917 26741 5951 26775
rect 7389 26741 7423 26775
rect 11069 26741 11103 26775
rect 13645 26741 13679 26775
rect 14933 26741 14967 26775
rect 15761 26741 15795 26775
rect 16957 26741 16991 26775
rect 17601 26741 17635 26775
rect 18245 26741 18279 26775
rect 20637 26741 20671 26775
rect 18797 26537 18831 26571
rect 22385 26537 22419 26571
rect 26525 26537 26559 26571
rect 28825 26537 28859 26571
rect 23029 26469 23063 26503
rect 36369 26469 36403 26503
rect 38209 26469 38243 26503
rect 4077 26401 4111 26435
rect 5273 26401 5307 26435
rect 10977 26401 11011 26435
rect 11989 26401 12023 26435
rect 13093 26401 13127 26435
rect 13369 26401 13403 26435
rect 14657 26401 14691 26435
rect 15669 26401 15703 26435
rect 16221 26401 16255 26435
rect 19625 26401 19659 26435
rect 20637 26401 20671 26435
rect 21189 26401 21223 26435
rect 27721 26401 27755 26435
rect 1593 26333 1627 26367
rect 5181 26333 5215 26367
rect 5825 26333 5859 26367
rect 6653 26333 6687 26367
rect 9873 26333 9907 26367
rect 17141 26333 17175 26367
rect 18061 26333 18095 26367
rect 18705 26333 18739 26367
rect 22293 26333 22327 26367
rect 22937 26333 22971 26367
rect 25329 26333 25363 26367
rect 26433 26333 26467 26367
rect 27077 26333 27111 26367
rect 28733 26333 28767 26367
rect 36553 26333 36587 26367
rect 38025 26333 38059 26367
rect 2697 26265 2731 26299
rect 2789 26265 2823 26299
rect 3341 26265 3375 26299
rect 4169 26265 4203 26299
rect 4721 26265 4755 26299
rect 5917 26265 5951 26299
rect 7481 26265 7515 26299
rect 7573 26265 7607 26299
rect 8493 26265 8527 26299
rect 9229 26265 9263 26299
rect 9321 26265 9355 26299
rect 11069 26265 11103 26299
rect 13185 26265 13219 26299
rect 14381 26265 14415 26299
rect 14473 26265 14507 26299
rect 15761 26265 15795 26299
rect 18153 26265 18187 26299
rect 19717 26265 19751 26299
rect 21281 26265 21315 26299
rect 21833 26265 21867 26299
rect 1777 26197 1811 26231
rect 6745 26197 6779 26231
rect 17233 26197 17267 26231
rect 25421 26197 25455 26231
rect 27169 26197 27203 26231
rect 6745 25993 6779 26027
rect 22753 25993 22787 26027
rect 23397 25993 23431 26027
rect 30665 25993 30699 26027
rect 2329 25925 2363 25959
rect 4169 25925 4203 25959
rect 5365 25925 5399 25959
rect 8033 25925 8067 25959
rect 8125 25925 8159 25959
rect 10149 25925 10183 25959
rect 11805 25925 11839 25959
rect 11897 25925 11931 25959
rect 17785 25925 17819 25959
rect 19533 25925 19567 25959
rect 20453 25925 20487 25959
rect 25605 25925 25639 25959
rect 27353 25925 27387 25959
rect 27905 25925 27939 25959
rect 6653 25857 6687 25891
rect 7297 25857 7331 25891
rect 13277 25857 13311 25891
rect 13921 25857 13955 25891
rect 14565 25857 14599 25891
rect 15209 25857 15243 25891
rect 15853 25857 15887 25891
rect 16865 25857 16899 25891
rect 17693 25857 17727 25891
rect 18337 25857 18371 25891
rect 20913 25857 20947 25891
rect 22017 25857 22051 25891
rect 22661 25857 22695 25891
rect 23305 25857 23339 25891
rect 30573 25857 30607 25891
rect 2237 25789 2271 25823
rect 3249 25789 3283 25823
rect 4077 25789 4111 25823
rect 4353 25789 4387 25823
rect 5273 25789 5307 25823
rect 5917 25789 5951 25823
rect 8401 25789 8435 25823
rect 10057 25789 10091 25823
rect 10333 25789 10367 25823
rect 12817 25789 12851 25823
rect 15301 25789 15335 25823
rect 16957 25789 16991 25823
rect 19441 25789 19475 25823
rect 25513 25789 25547 25823
rect 26341 25789 26375 25823
rect 27261 25789 27295 25823
rect 14657 25721 14691 25755
rect 7389 25653 7423 25687
rect 13369 25653 13403 25687
rect 14013 25653 14047 25687
rect 15945 25653 15979 25687
rect 18429 25653 18463 25687
rect 21005 25653 21039 25687
rect 22109 25653 22143 25687
rect 1777 25449 1811 25483
rect 15577 25449 15611 25483
rect 29929 25449 29963 25483
rect 21097 25381 21131 25415
rect 4905 25313 4939 25347
rect 5917 25313 5951 25347
rect 9690 25313 9724 25347
rect 14933 25313 14967 25347
rect 19533 25313 19567 25347
rect 19809 25313 19843 25347
rect 22109 25313 22143 25347
rect 22385 25313 22419 25347
rect 26249 25313 26283 25347
rect 1961 25245 1995 25279
rect 4169 25245 4203 25279
rect 4261 25245 4295 25279
rect 6377 25245 6411 25279
rect 11345 25245 11379 25279
rect 13553 25245 13587 25279
rect 14833 25245 14867 25279
rect 15485 25245 15519 25279
rect 18061 25245 18095 25279
rect 18705 25245 18739 25279
rect 21005 25245 21039 25279
rect 23765 25245 23799 25279
rect 28549 25245 28583 25279
rect 30113 25245 30147 25279
rect 38025 25245 38059 25279
rect 2513 25177 2547 25211
rect 3249 25177 3283 25211
rect 4997 25177 5031 25211
rect 6653 25177 6687 25211
rect 9774 25177 9808 25211
rect 10701 25177 10735 25211
rect 11621 25177 11655 25211
rect 16221 25177 16255 25211
rect 16313 25177 16347 25211
rect 17233 25177 17267 25211
rect 19625 25177 19659 25211
rect 22201 25177 22235 25211
rect 26341 25177 26375 25211
rect 26893 25177 26927 25211
rect 37657 25177 37691 25211
rect 8125 25109 8159 25143
rect 13093 25109 13127 25143
rect 13645 25109 13679 25143
rect 18153 25109 18187 25143
rect 18797 25109 18831 25143
rect 23857 25109 23891 25143
rect 28641 25109 28675 25143
rect 38209 25109 38243 25143
rect 22753 24905 22787 24939
rect 26433 24905 26467 24939
rect 1869 24837 1903 24871
rect 4261 24837 4295 24871
rect 5181 24837 5215 24871
rect 6745 24837 6779 24871
rect 8677 24837 8711 24871
rect 11989 24837 12023 24871
rect 14105 24837 14139 24871
rect 15761 24837 15795 24871
rect 17049 24837 17083 24871
rect 17969 24837 18003 24871
rect 19349 24837 19383 24871
rect 20821 24837 20855 24871
rect 20913 24837 20947 24871
rect 23489 24837 23523 24871
rect 24409 24837 24443 24871
rect 25053 24837 25087 24871
rect 28273 24837 28307 24871
rect 28825 24837 28859 24871
rect 3249 24769 3283 24803
rect 7757 24769 7791 24803
rect 10977 24769 11011 24803
rect 18521 24769 18555 24803
rect 22017 24769 22051 24803
rect 22661 24769 22695 24803
rect 25605 24769 25639 24803
rect 26341 24769 26375 24803
rect 37565 24769 37599 24803
rect 1777 24701 1811 24735
rect 2789 24701 2823 24735
rect 4169 24701 4203 24735
rect 5825 24701 5859 24735
rect 6653 24701 6687 24735
rect 8401 24701 8435 24735
rect 11713 24701 11747 24735
rect 14013 24701 14047 24735
rect 15025 24701 15059 24735
rect 15669 24701 15703 24735
rect 16313 24701 16347 24735
rect 16957 24701 16991 24735
rect 19257 24701 19291 24735
rect 19533 24701 19567 24735
rect 23397 24701 23431 24735
rect 24961 24701 24995 24735
rect 28181 24701 28215 24735
rect 7205 24633 7239 24667
rect 10149 24633 10183 24667
rect 11069 24633 11103 24667
rect 13461 24633 13495 24667
rect 21373 24633 21407 24667
rect 3433 24565 3467 24599
rect 7849 24565 7883 24599
rect 18613 24565 18647 24599
rect 22109 24565 22143 24599
rect 37657 24565 37691 24599
rect 4077 24361 4111 24395
rect 8585 24361 8619 24395
rect 9768 24361 9802 24395
rect 14657 24361 14691 24395
rect 16129 24361 16163 24395
rect 28181 24361 28215 24395
rect 19717 24293 19751 24327
rect 23765 24293 23799 24327
rect 1593 24225 1627 24259
rect 6377 24225 6411 24259
rect 9505 24225 9539 24259
rect 11713 24225 11747 24259
rect 15485 24225 15519 24259
rect 20269 24225 20303 24259
rect 20729 24225 20763 24259
rect 24685 24225 24719 24259
rect 25329 24225 25363 24259
rect 3985 24157 4019 24191
rect 4629 24157 4663 24191
rect 6837 24157 6871 24191
rect 15393 24157 15427 24191
rect 16037 24157 16071 24191
rect 18705 24157 18739 24191
rect 18797 24157 18831 24191
rect 21833 24157 21867 24191
rect 22477 24157 22511 24191
rect 26433 24157 26467 24191
rect 28089 24157 28123 24191
rect 30021 24157 30055 24191
rect 37473 24157 37507 24191
rect 37749 24157 37783 24191
rect 1869 24089 1903 24123
rect 4905 24089 4939 24123
rect 7113 24089 7147 24123
rect 11989 24089 12023 24123
rect 13737 24089 13771 24123
rect 14565 24089 14599 24123
rect 16773 24089 16807 24123
rect 16865 24089 16899 24123
rect 17785 24089 17819 24123
rect 19533 24089 19567 24123
rect 20361 24089 20395 24123
rect 23213 24089 23247 24123
rect 23305 24089 23339 24123
rect 24777 24089 24811 24123
rect 3341 24021 3375 24055
rect 11253 24021 11287 24055
rect 21925 24021 21959 24055
rect 22569 24021 22603 24055
rect 26525 24021 26559 24055
rect 30113 24021 30147 24055
rect 30665 24021 30699 24055
rect 3617 23817 3651 23851
rect 23673 23817 23707 23851
rect 24961 23817 24995 23851
rect 7297 23749 7331 23783
rect 8033 23749 8067 23783
rect 14473 23749 14507 23783
rect 16221 23749 16255 23783
rect 17325 23749 17359 23783
rect 18797 23749 18831 23783
rect 18889 23749 18923 23783
rect 19809 23749 19843 23783
rect 20453 23749 20487 23783
rect 20545 23749 20579 23783
rect 22201 23749 22235 23783
rect 23121 23749 23155 23783
rect 27353 23749 27387 23783
rect 28641 23749 28675 23783
rect 30573 23749 30607 23783
rect 30665 23749 30699 23783
rect 4261 23681 4295 23715
rect 6561 23681 6595 23715
rect 7941 23681 7975 23715
rect 10609 23681 10643 23715
rect 16129 23681 16163 23715
rect 23581 23681 23615 23715
rect 24225 23681 24259 23715
rect 24869 23681 24903 23715
rect 25513 23681 25547 23715
rect 26157 23681 26191 23715
rect 29837 23681 29871 23715
rect 1869 23613 1903 23647
rect 2145 23613 2179 23647
rect 4537 23613 4571 23647
rect 8585 23613 8619 23647
rect 8861 23613 8895 23647
rect 11805 23613 11839 23647
rect 12081 23613 12115 23647
rect 13829 23613 13863 23647
rect 14381 23613 14415 23647
rect 14657 23613 14691 23647
rect 17233 23613 17267 23647
rect 17509 23613 17543 23647
rect 21097 23613 21131 23647
rect 22109 23613 22143 23647
rect 27261 23613 27295 23647
rect 27905 23613 27939 23647
rect 28549 23613 28583 23647
rect 29193 23613 29227 23647
rect 30849 23613 30883 23647
rect 6009 23545 6043 23579
rect 24317 23477 24351 23511
rect 25605 23477 25639 23511
rect 26249 23477 26283 23511
rect 29653 23477 29687 23511
rect 5733 23273 5767 23307
rect 23489 23273 23523 23307
rect 15945 23205 15979 23239
rect 1593 23137 1627 23171
rect 3985 23137 4019 23171
rect 6837 23137 6871 23171
rect 9597 23137 9631 23171
rect 13737 23137 13771 23171
rect 17417 23137 17451 23171
rect 18245 23137 18279 23171
rect 19901 23137 19935 23171
rect 24685 23137 24719 23171
rect 24961 23137 24995 23171
rect 26801 23137 26835 23171
rect 28641 23137 28675 23171
rect 6561 23069 6595 23103
rect 9321 23069 9355 23103
rect 11713 23069 11747 23103
rect 15853 23069 15887 23103
rect 23397 23069 23431 23103
rect 29745 23069 29779 23103
rect 1869 23001 1903 23035
rect 4261 23001 4295 23035
rect 8585 23001 8619 23035
rect 11989 23001 12023 23035
rect 14381 23001 14415 23035
rect 14473 23001 14507 23035
rect 15393 23001 15427 23035
rect 16589 23001 16623 23035
rect 16681 23001 16715 23035
rect 18337 23001 18371 23035
rect 18889 23001 18923 23035
rect 19993 23001 20027 23035
rect 20913 23001 20947 23035
rect 21925 23001 21959 23035
rect 22017 23001 22051 23035
rect 22937 23001 22971 23035
rect 24777 23001 24811 23035
rect 26893 23001 26927 23035
rect 27813 23001 27847 23035
rect 28365 23001 28399 23035
rect 28457 23001 28491 23035
rect 3341 22933 3375 22967
rect 11069 22933 11103 22967
rect 29837 22933 29871 22967
rect 5917 22729 5951 22763
rect 27261 22729 27295 22763
rect 28089 22729 28123 22763
rect 4445 22661 4479 22695
rect 6745 22661 6779 22695
rect 12173 22661 12207 22695
rect 14289 22661 14323 22695
rect 16221 22661 16255 22695
rect 17049 22661 17083 22695
rect 18521 22661 18555 22695
rect 18613 22661 18647 22695
rect 22385 22661 22419 22695
rect 23949 22661 23983 22695
rect 25973 22661 26007 22695
rect 26065 22661 26099 22695
rect 29377 22661 29411 22695
rect 4169 22593 4203 22627
rect 7297 22593 7331 22627
rect 7757 22593 7791 22627
rect 10241 22593 10275 22627
rect 16129 22593 16163 22627
rect 20453 22593 20487 22627
rect 21097 22593 21131 22627
rect 27169 22593 27203 22627
rect 27997 22593 28031 22627
rect 30757 22593 30791 22627
rect 38025 22593 38059 22627
rect 1869 22525 1903 22559
rect 2145 22525 2179 22559
rect 6653 22525 6687 22559
rect 8033 22525 8067 22559
rect 9781 22525 9815 22559
rect 10977 22525 11011 22559
rect 11897 22525 11931 22559
rect 13645 22525 13679 22559
rect 14197 22525 14231 22559
rect 14565 22525 14599 22559
rect 16957 22525 16991 22559
rect 17233 22525 17267 22559
rect 18797 22525 18831 22559
rect 22293 22525 22327 22559
rect 22569 22525 22603 22559
rect 23857 22525 23891 22559
rect 24869 22525 24903 22559
rect 29285 22525 29319 22559
rect 29561 22525 29595 22559
rect 3617 22457 3651 22491
rect 26525 22457 26559 22491
rect 30849 22457 30883 22491
rect 38209 22457 38243 22491
rect 20545 22389 20579 22423
rect 21189 22389 21223 22423
rect 4334 22185 4368 22219
rect 6548 22185 6582 22219
rect 18153 22185 18187 22219
rect 20085 22185 20119 22219
rect 24685 22185 24719 22219
rect 28917 22117 28951 22151
rect 1685 22049 1719 22083
rect 1961 22049 1995 22083
rect 3433 22049 3467 22083
rect 6285 22049 6319 22083
rect 9229 22049 9263 22083
rect 10057 22049 10091 22083
rect 10609 22049 10643 22083
rect 11621 22049 11655 22083
rect 13369 22049 13403 22083
rect 14657 22049 14691 22083
rect 15301 22049 15335 22083
rect 20729 22049 20763 22083
rect 21373 22049 21407 22083
rect 22293 22049 22327 22083
rect 24041 22049 24075 22083
rect 26985 22049 27019 22083
rect 4077 21981 4111 22015
rect 10517 21981 10551 22015
rect 11345 21981 11379 22015
rect 14565 21981 14599 22015
rect 17141 21981 17175 22015
rect 18061 21981 18095 22015
rect 18705 21981 18739 22015
rect 19993 21981 20027 22015
rect 22201 21981 22235 22015
rect 24593 21981 24627 22015
rect 26893 21981 26927 22015
rect 34161 21981 34195 22015
rect 38301 21981 38335 22015
rect 9321 21913 9355 21947
rect 11069 21913 11103 21947
rect 15370 21913 15404 21947
rect 15945 21913 15979 21947
rect 16497 21913 16531 21947
rect 16589 21913 16623 21947
rect 20821 21913 20855 21947
rect 23397 21913 23431 21947
rect 23489 21913 23523 21947
rect 28365 21913 28399 21947
rect 28457 21913 28491 21947
rect 5825 21845 5859 21879
rect 8033 21845 8067 21879
rect 18797 21845 18831 21879
rect 33977 21845 34011 21879
rect 38117 21845 38151 21879
rect 4629 21641 4663 21675
rect 11345 21641 11379 21675
rect 21281 21641 21315 21675
rect 23581 21641 23615 21675
rect 24225 21641 24259 21675
rect 38209 21641 38243 21675
rect 3157 21573 3191 21607
rect 5457 21573 5491 21607
rect 7849 21573 7883 21607
rect 9597 21573 9631 21607
rect 10793 21573 10827 21607
rect 11897 21573 11931 21607
rect 13737 21573 13771 21607
rect 14289 21573 14323 21607
rect 15761 21573 15795 21607
rect 18521 21573 18555 21607
rect 18613 21573 18647 21607
rect 19809 21573 19843 21607
rect 26525 21573 26559 21607
rect 27353 21573 27387 21607
rect 28917 21573 28951 21607
rect 1593 21505 1627 21539
rect 2881 21505 2915 21539
rect 6929 21505 6963 21539
rect 7573 21505 7607 21539
rect 10057 21505 10091 21539
rect 14933 21505 14967 21539
rect 16313 21505 16347 21539
rect 17141 21505 17175 21539
rect 17785 21505 17819 21539
rect 21189 21505 21223 21539
rect 22017 21505 22051 21539
rect 22845 21505 22879 21539
rect 23489 21505 23523 21539
rect 24133 21505 24167 21539
rect 24777 21505 24811 21539
rect 25421 21505 25455 21539
rect 26433 21505 26467 21539
rect 29929 21505 29963 21539
rect 38117 21505 38151 21539
rect 1869 21437 1903 21471
rect 5365 21437 5399 21471
rect 11805 21437 11839 21471
rect 12817 21437 12851 21471
rect 13645 21437 13679 21471
rect 15669 21437 15703 21471
rect 17877 21437 17911 21471
rect 19717 21437 19751 21471
rect 20269 21437 20303 21471
rect 25513 21437 25547 21471
rect 27261 21437 27295 21471
rect 27537 21437 27571 21471
rect 28825 21437 28859 21471
rect 30021 21437 30055 21471
rect 5917 21369 5951 21403
rect 17233 21369 17267 21403
rect 19073 21369 19107 21403
rect 29377 21369 29411 21403
rect 7021 21301 7055 21335
rect 15025 21301 15059 21335
rect 22109 21301 22143 21335
rect 22937 21301 22971 21335
rect 24869 21301 24903 21335
rect 12725 21097 12759 21131
rect 16405 21097 16439 21131
rect 29837 21097 29871 21131
rect 3341 21029 3375 21063
rect 18797 21029 18831 21063
rect 25789 21029 25823 21063
rect 1593 20961 1627 20995
rect 4905 20961 4939 20995
rect 7573 20961 7607 20995
rect 10241 20961 10275 20995
rect 11253 20961 11287 20995
rect 19533 20961 19567 20995
rect 20545 20961 20579 20995
rect 22293 20961 22327 20995
rect 25237 20961 25271 20995
rect 28549 20961 28583 20995
rect 3985 20893 4019 20927
rect 10977 20893 11011 20927
rect 13553 20893 13587 20927
rect 16313 20893 16347 20927
rect 18705 20893 18739 20927
rect 21557 20893 21591 20927
rect 22201 20893 22235 20927
rect 22845 20893 22879 20927
rect 23489 20893 23523 20927
rect 26341 20893 26375 20927
rect 27813 20893 27847 20927
rect 29745 20893 29779 20927
rect 1869 20825 1903 20859
rect 5181 20825 5215 20859
rect 6929 20825 6963 20859
rect 7665 20825 7699 20859
rect 8585 20825 8619 20859
rect 9229 20825 9263 20859
rect 9321 20825 9355 20859
rect 14381 20825 14415 20859
rect 14473 20825 14507 20859
rect 15393 20825 15427 20859
rect 17049 20825 17083 20859
rect 17141 20825 17175 20859
rect 18061 20825 18095 20859
rect 19625 20825 19659 20859
rect 25329 20825 25363 20859
rect 26433 20825 26467 20859
rect 28641 20825 28675 20859
rect 29193 20825 29227 20859
rect 4169 20757 4203 20791
rect 13645 20757 13679 20791
rect 21649 20757 21683 20791
rect 22937 20757 22971 20791
rect 23581 20757 23615 20791
rect 27905 20757 27939 20791
rect 14657 20553 14691 20587
rect 17417 20553 17451 20587
rect 25053 20553 25087 20587
rect 26249 20553 26283 20587
rect 28457 20553 28491 20587
rect 4997 20485 5031 20519
rect 5089 20485 5123 20519
rect 6653 20485 6687 20519
rect 7665 20485 7699 20519
rect 9965 20485 9999 20519
rect 10885 20485 10919 20519
rect 13737 20485 13771 20519
rect 15393 20485 15427 20519
rect 18797 20485 18831 20519
rect 19717 20485 19751 20519
rect 20269 20485 20303 20519
rect 22385 20485 22419 20519
rect 1869 20417 1903 20451
rect 7389 20417 7423 20451
rect 9505 20417 9539 20451
rect 14565 20417 14599 20451
rect 17325 20417 17359 20451
rect 17969 20417 18003 20451
rect 20913 20417 20947 20451
rect 23397 20417 23431 20451
rect 24317 20417 24351 20451
rect 24961 20417 24995 20451
rect 25605 20417 25639 20451
rect 26433 20417 26467 20451
rect 27169 20417 27203 20451
rect 28365 20417 28399 20451
rect 29009 20417 29043 20451
rect 29653 20417 29687 20451
rect 2145 20349 2179 20383
rect 3893 20349 3927 20383
rect 6009 20349 6043 20383
rect 9137 20349 9171 20383
rect 9873 20349 9907 20383
rect 11713 20349 11747 20383
rect 11976 20349 12010 20383
rect 15301 20349 15335 20383
rect 16129 20349 16163 20383
rect 18705 20349 18739 20383
rect 22293 20349 22327 20383
rect 25697 20349 25731 20383
rect 22845 20281 22879 20315
rect 27261 20281 27295 20315
rect 6745 20213 6779 20247
rect 18061 20213 18095 20247
rect 20361 20213 20395 20247
rect 21005 20213 21039 20247
rect 23489 20213 23523 20247
rect 24409 20213 24443 20247
rect 29101 20213 29135 20247
rect 29745 20213 29779 20247
rect 1856 20009 1890 20043
rect 3341 20009 3375 20043
rect 8493 20009 8527 20043
rect 13645 20009 13679 20043
rect 21097 20009 21131 20043
rect 23673 20009 23707 20043
rect 18153 19941 18187 19975
rect 27721 19941 27755 19975
rect 1593 19873 1627 19907
rect 4077 19873 4111 19907
rect 5917 19873 5951 19907
rect 10241 19873 10275 19907
rect 10885 19873 10919 19907
rect 17049 19873 17083 19907
rect 19533 19873 19567 19907
rect 19809 19873 19843 19907
rect 8401 19805 8435 19839
rect 13553 19805 13587 19839
rect 18705 19805 18739 19839
rect 21005 19805 21039 19839
rect 21649 19805 21683 19839
rect 23581 19805 23615 19839
rect 24593 19805 24627 19839
rect 26341 19805 26375 19839
rect 26985 19805 27019 19839
rect 27629 19805 27663 19839
rect 28273 19805 28307 19839
rect 28917 19805 28951 19839
rect 31033 19805 31067 19839
rect 38301 19805 38335 19839
rect 4169 19737 4203 19771
rect 5089 19737 5123 19771
rect 6193 19737 6227 19771
rect 9218 19737 9252 19771
rect 9321 19737 9355 19771
rect 11161 19737 11195 19771
rect 12909 19737 12943 19771
rect 14381 19737 14415 19771
rect 14473 19737 14507 19771
rect 15393 19737 15427 19771
rect 16037 19737 16071 19771
rect 16129 19737 16163 19771
rect 17601 19737 17635 19771
rect 17693 19737 17727 19771
rect 19634 19737 19668 19771
rect 22477 19737 22511 19771
rect 22569 19737 22603 19771
rect 23121 19737 23155 19771
rect 25697 19737 25731 19771
rect 29929 19737 29963 19771
rect 30021 19737 30055 19771
rect 30573 19737 30607 19771
rect 7665 19669 7699 19703
rect 18797 19669 18831 19703
rect 21741 19669 21775 19703
rect 24685 19669 24719 19703
rect 25789 19669 25823 19703
rect 26433 19669 26467 19703
rect 27077 19669 27111 19703
rect 28365 19669 28399 19703
rect 29009 19669 29043 19703
rect 31125 19669 31159 19703
rect 38117 19669 38151 19703
rect 3525 19465 3559 19499
rect 20177 19465 20211 19499
rect 31585 19465 31619 19499
rect 37657 19465 37691 19499
rect 6009 19397 6043 19431
rect 9505 19397 9539 19431
rect 10149 19397 10183 19431
rect 12173 19397 12207 19431
rect 12265 19397 12299 19431
rect 13737 19397 13771 19431
rect 13829 19397 13863 19431
rect 14749 19397 14783 19431
rect 15301 19397 15335 19431
rect 15393 19397 15427 19431
rect 16313 19397 16347 19431
rect 16957 19397 16991 19431
rect 17049 19397 17083 19431
rect 18705 19397 18739 19431
rect 20821 19397 20855 19431
rect 20913 19397 20947 19431
rect 22477 19397 22511 19431
rect 22569 19397 22603 19431
rect 24041 19397 24075 19431
rect 24133 19397 24167 19431
rect 25605 19397 25639 19431
rect 25697 19397 25731 19431
rect 26617 19397 26651 19431
rect 27353 19397 27387 19431
rect 28273 19397 28307 19431
rect 28825 19397 28859 19431
rect 28917 19397 28951 19431
rect 29837 19397 29871 19431
rect 30389 19397 30423 19431
rect 30481 19397 30515 19431
rect 1777 19329 1811 19363
rect 6837 19329 6871 19363
rect 7481 19329 7515 19363
rect 20085 19329 20119 19363
rect 31493 19329 31527 19363
rect 37841 19329 37875 19363
rect 2053 19261 2087 19295
rect 3985 19261 4019 19295
rect 4261 19261 4295 19295
rect 7757 19261 7791 19295
rect 10057 19261 10091 19295
rect 10885 19261 10919 19295
rect 13185 19261 13219 19295
rect 17601 19261 17635 19295
rect 18613 19261 18647 19295
rect 18889 19261 18923 19295
rect 21097 19261 21131 19295
rect 23397 19261 23431 19295
rect 27261 19261 27295 19295
rect 30665 19261 30699 19295
rect 24593 19193 24627 19227
rect 6929 19125 6963 19159
rect 3341 18921 3375 18955
rect 9321 18921 9355 18955
rect 26893 18921 26927 18955
rect 11621 18853 11655 18887
rect 1593 18785 1627 18819
rect 3985 18785 4019 18819
rect 4261 18785 4295 18819
rect 6009 18785 6043 18819
rect 12357 18785 12391 18819
rect 18889 18785 18923 18819
rect 19901 18785 19935 18819
rect 20545 18785 20579 18819
rect 21097 18785 21131 18819
rect 22293 18785 22327 18819
rect 22937 18785 22971 18819
rect 25697 18785 25731 18819
rect 29837 18785 29871 18819
rect 30113 18785 30147 18819
rect 31217 18785 31251 18819
rect 31493 18785 31527 18819
rect 6561 18717 6595 18751
rect 9229 18717 9263 18751
rect 9873 18717 9907 18751
rect 15853 18717 15887 18751
rect 17693 18717 17727 18751
rect 23765 18717 23799 18751
rect 26157 18717 26191 18751
rect 26801 18717 26835 18751
rect 28641 18717 28675 18751
rect 32689 18717 32723 18751
rect 38301 18717 38335 18751
rect 1869 18649 1903 18683
rect 6837 18649 6871 18683
rect 8585 18649 8619 18683
rect 10149 18649 10183 18683
rect 12449 18649 12483 18683
rect 13369 18649 13403 18683
rect 14381 18649 14415 18683
rect 14473 18649 14507 18683
rect 15393 18649 15427 18683
rect 16129 18649 16163 18683
rect 17038 18649 17072 18683
rect 17134 18649 17168 18683
rect 18245 18649 18279 18683
rect 18337 18649 18371 18683
rect 19986 18649 20020 18683
rect 21189 18649 21223 18683
rect 21741 18649 21775 18683
rect 22385 18649 22419 18683
rect 25053 18649 25087 18683
rect 25145 18649 25179 18683
rect 27537 18649 27571 18683
rect 27629 18649 27663 18683
rect 28181 18649 28215 18683
rect 29929 18649 29963 18683
rect 31309 18649 31343 18683
rect 23857 18581 23891 18615
rect 26249 18581 26283 18615
rect 28733 18581 28767 18615
rect 32781 18581 32815 18615
rect 38117 18581 38151 18615
rect 18981 18377 19015 18411
rect 30849 18377 30883 18411
rect 2237 18309 2271 18343
rect 3157 18309 3191 18343
rect 5641 18309 5675 18343
rect 12449 18309 12483 18343
rect 13369 18309 13403 18343
rect 14197 18309 14231 18343
rect 15393 18309 15427 18343
rect 16957 18309 16991 18343
rect 17049 18309 17083 18343
rect 19625 18309 19659 18343
rect 19717 18309 19751 18343
rect 20913 18309 20947 18343
rect 23213 18309 23247 18343
rect 23305 18309 23339 18343
rect 24869 18309 24903 18343
rect 25973 18309 26007 18343
rect 26065 18309 26099 18343
rect 28733 18309 28767 18343
rect 9328 18241 9362 18275
rect 18889 18241 18923 18275
rect 20269 18241 20303 18275
rect 22017 18241 22051 18275
rect 25421 18241 25455 18275
rect 27169 18241 27203 18275
rect 27813 18241 27847 18275
rect 30113 18241 30147 18275
rect 30757 18241 30791 18275
rect 31401 18241 31435 18275
rect 2145 18173 2179 18207
rect 3617 18173 3651 18207
rect 3893 18173 3927 18207
rect 6837 18173 6871 18207
rect 7113 18173 7147 18207
rect 8861 18173 8895 18207
rect 12357 18173 12391 18207
rect 14105 18173 14139 18207
rect 14381 18173 14415 18207
rect 15301 18173 15335 18207
rect 16313 18173 16347 18207
rect 17969 18173 18003 18207
rect 20821 18173 20855 18207
rect 24225 18173 24259 18207
rect 24777 18173 24811 18207
rect 26341 18173 26375 18207
rect 28641 18173 28675 18207
rect 29653 18173 29687 18207
rect 21373 18105 21407 18139
rect 27261 18105 27295 18139
rect 9578 18037 9612 18071
rect 11069 18037 11103 18071
rect 22109 18037 22143 18071
rect 27905 18037 27939 18071
rect 30205 18037 30239 18071
rect 31493 18037 31527 18071
rect 1948 17833 1982 17867
rect 22017 17833 22051 17867
rect 25881 17833 25915 17867
rect 3433 17765 3467 17799
rect 21373 17765 21407 17799
rect 31677 17765 31711 17799
rect 1685 17697 1719 17731
rect 3985 17697 4019 17731
rect 6009 17697 6043 17731
rect 6469 17697 6503 17731
rect 9873 17697 9907 17731
rect 13369 17697 13403 17731
rect 15393 17697 15427 17731
rect 16129 17697 16163 17731
rect 17049 17697 17083 17731
rect 17693 17697 17727 17731
rect 20821 17697 20855 17731
rect 26525 17697 26559 17731
rect 27537 17697 27571 17731
rect 8493 17629 8527 17663
rect 10609 17629 10643 17663
rect 12633 17629 12667 17663
rect 13093 17629 13127 17663
rect 18337 17629 18371 17663
rect 21925 17629 21959 17663
rect 22569 17629 22603 17663
rect 23213 17629 23247 17663
rect 23857 17629 23891 17663
rect 25789 17629 25823 17663
rect 26433 17629 26467 17663
rect 28733 17629 28767 17663
rect 31125 17629 31159 17663
rect 31585 17629 31619 17663
rect 4261 17561 4295 17595
rect 6745 17561 6779 17595
rect 9154 17561 9188 17595
rect 10885 17561 10919 17595
rect 14381 17561 14415 17595
rect 14473 17561 14507 17595
rect 16221 17561 16255 17595
rect 17778 17561 17812 17595
rect 19533 17561 19567 17595
rect 19625 17561 19659 17595
rect 20177 17561 20211 17595
rect 20922 17561 20956 17595
rect 24685 17561 24719 17595
rect 24777 17561 24811 17595
rect 25329 17561 25363 17595
rect 27261 17561 27295 17595
rect 27353 17561 27387 17595
rect 29837 17561 29871 17595
rect 29929 17561 29963 17595
rect 30481 17561 30515 17595
rect 22661 17493 22695 17527
rect 23305 17493 23339 17527
rect 23949 17493 23983 17527
rect 28825 17493 28859 17527
rect 30941 17493 30975 17527
rect 1777 17289 1811 17323
rect 24041 17289 24075 17323
rect 28457 17289 28491 17323
rect 4353 17221 4387 17255
rect 4905 17221 4939 17255
rect 4997 17221 5031 17255
rect 6929 17221 6963 17255
rect 9137 17221 9171 17255
rect 11989 17221 12023 17255
rect 14105 17221 14139 17255
rect 15393 17221 15427 17255
rect 16313 17221 16347 17255
rect 17049 17221 17083 17255
rect 18797 17221 18831 17255
rect 19717 17221 19751 17255
rect 20545 17221 20579 17255
rect 22201 17221 22235 17255
rect 22293 17221 22327 17255
rect 23397 17221 23431 17255
rect 24869 17221 24903 17255
rect 25421 17221 25455 17255
rect 27353 17221 27387 17255
rect 29469 17221 29503 17255
rect 1593 17153 1627 17187
rect 2329 17153 2363 17187
rect 6653 17153 6687 17187
rect 8861 17153 8895 17187
rect 11713 17153 11747 17187
rect 22845 17153 22879 17187
rect 23305 17153 23339 17187
rect 23949 17153 23983 17187
rect 25881 17153 25915 17187
rect 28365 17153 28399 17187
rect 30481 17153 30515 17187
rect 37749 17153 37783 17187
rect 2605 17085 2639 17119
rect 5181 17085 5215 17119
rect 10885 17085 10919 17119
rect 13461 17085 13495 17119
rect 14013 17085 14047 17119
rect 15301 17085 15335 17119
rect 16957 17085 16991 17119
rect 17969 17085 18003 17119
rect 18705 17085 18739 17119
rect 20453 17085 20487 17119
rect 21465 17085 21499 17119
rect 24777 17085 24811 17119
rect 27261 17085 27295 17119
rect 27537 17085 27571 17119
rect 29377 17085 29411 17119
rect 37473 17085 37507 17119
rect 8401 17017 8435 17051
rect 14565 17017 14599 17051
rect 29929 17017 29963 17051
rect 2237 16949 2271 16983
rect 25973 16949 26007 16983
rect 30573 16949 30607 16983
rect 4077 16745 4111 16779
rect 23029 16745 23063 16779
rect 23673 16745 23707 16779
rect 38209 16745 38243 16779
rect 1685 16609 1719 16643
rect 4353 16609 4387 16643
rect 6561 16609 6595 16643
rect 6837 16609 6871 16643
rect 9873 16609 9907 16643
rect 10609 16609 10643 16643
rect 15485 16609 15519 16643
rect 17325 16609 17359 16643
rect 20729 16609 20763 16643
rect 21465 16609 21499 16643
rect 22477 16609 22511 16643
rect 8585 16541 8619 16575
rect 13093 16541 13127 16575
rect 14473 16541 14507 16575
rect 20637 16541 20671 16575
rect 22937 16541 22971 16575
rect 23581 16541 23615 16575
rect 27721 16541 27755 16575
rect 28365 16541 28399 16575
rect 28457 16541 28491 16575
rect 29009 16541 29043 16575
rect 29101 16541 29135 16575
rect 29745 16541 29779 16575
rect 30389 16541 30423 16575
rect 31033 16541 31067 16575
rect 1961 16473 1995 16507
rect 4629 16473 4663 16507
rect 9137 16473 9171 16507
rect 10885 16473 10919 16507
rect 12633 16473 12667 16507
rect 13369 16473 13403 16507
rect 14565 16473 14599 16507
rect 15209 16473 15243 16507
rect 15301 16473 15335 16507
rect 17417 16473 17451 16507
rect 18337 16473 18371 16507
rect 19533 16473 19567 16507
rect 19625 16473 19659 16507
rect 20177 16473 20211 16507
rect 21557 16473 21591 16507
rect 24685 16473 24719 16507
rect 24777 16473 24811 16507
rect 25697 16473 25731 16507
rect 26249 16473 26283 16507
rect 26341 16473 26375 16507
rect 27261 16473 27295 16507
rect 29837 16473 29871 16507
rect 38117 16473 38151 16507
rect 3433 16405 3467 16439
rect 6101 16405 6135 16439
rect 27813 16405 27847 16439
rect 30481 16405 30515 16439
rect 31125 16405 31159 16439
rect 5411 16201 5445 16235
rect 7113 16201 7147 16235
rect 26249 16201 26283 16235
rect 27261 16201 27295 16235
rect 31585 16201 31619 16235
rect 35909 16201 35943 16235
rect 7941 16133 7975 16167
rect 10977 16133 11011 16167
rect 15393 16133 15427 16167
rect 16313 16133 16347 16167
rect 17042 16133 17076 16167
rect 18797 16133 18831 16167
rect 18889 16133 18923 16167
rect 20637 16133 20671 16167
rect 21281 16133 21315 16167
rect 22109 16133 22143 16167
rect 22201 16133 22235 16167
rect 24317 16133 24351 16167
rect 28273 16133 28307 16167
rect 29193 16133 29227 16167
rect 29745 16133 29779 16167
rect 29837 16133 29871 16167
rect 1685 16065 1719 16099
rect 2697 16065 2731 16099
rect 5181 16065 5215 16099
rect 7021 16065 7055 16099
rect 10241 16065 10275 16099
rect 11713 16065 11747 16099
rect 14197 16065 14231 16099
rect 19901 16065 19935 16099
rect 20545 16065 20579 16099
rect 21197 16055 21231 16089
rect 23581 16065 23615 16099
rect 24225 16065 24259 16099
rect 24869 16065 24903 16099
rect 25513 16065 25547 16099
rect 26157 16065 26191 16099
rect 27169 16065 27203 16099
rect 30849 16065 30883 16099
rect 31493 16065 31527 16099
rect 36093 16065 36127 16099
rect 2973 15997 3007 16031
rect 4721 15997 4755 16031
rect 7665 15997 7699 16031
rect 9689 15997 9723 16031
rect 11989 15997 12023 16031
rect 13737 15997 13771 16031
rect 14381 15997 14415 16031
rect 15301 15997 15335 16031
rect 16957 15997 16991 16031
rect 17969 15997 18003 16031
rect 23121 15997 23155 16031
rect 28181 15997 28215 16031
rect 30021 15997 30055 16031
rect 19349 15929 19383 15963
rect 25605 15929 25639 15963
rect 1777 15861 1811 15895
rect 19993 15861 20027 15895
rect 23673 15861 23707 15895
rect 24961 15861 24995 15895
rect 30941 15861 30975 15895
rect 3341 15657 3375 15691
rect 4077 15657 4111 15691
rect 11069 15657 11103 15691
rect 26525 15657 26559 15691
rect 27169 15657 27203 15691
rect 16037 15589 16071 15623
rect 28917 15589 28951 15623
rect 1593 15521 1627 15555
rect 4905 15521 4939 15555
rect 5641 15521 5675 15555
rect 7389 15521 7423 15555
rect 9321 15521 9355 15555
rect 11529 15521 11563 15555
rect 14289 15521 14323 15555
rect 17877 15521 17911 15555
rect 18889 15521 18923 15555
rect 23949 15521 23983 15555
rect 25329 15521 25363 15555
rect 28365 15521 28399 15555
rect 5365 15453 5399 15487
rect 8585 15453 8619 15487
rect 17233 15453 17267 15487
rect 19441 15453 19475 15487
rect 24593 15453 24627 15487
rect 25973 15453 26007 15487
rect 26433 15453 26467 15487
rect 27077 15453 27111 15487
rect 29745 15453 29779 15487
rect 30389 15453 30423 15487
rect 31033 15453 31067 15487
rect 38025 15453 38059 15487
rect 1869 15385 1903 15419
rect 4169 15385 4203 15419
rect 7941 15385 7975 15419
rect 8033 15385 8067 15419
rect 9597 15385 9631 15419
rect 11805 15385 11839 15419
rect 14565 15385 14599 15419
rect 16589 15385 16623 15419
rect 16681 15385 16715 15419
rect 17969 15385 18003 15419
rect 20637 15385 20671 15419
rect 21373 15385 21407 15419
rect 21465 15385 21499 15419
rect 22385 15385 22419 15419
rect 22937 15385 22971 15419
rect 23029 15385 23063 15419
rect 25421 15385 25455 15419
rect 28457 15385 28491 15419
rect 31125 15385 31159 15419
rect 13277 15317 13311 15351
rect 19533 15317 19567 15351
rect 20729 15317 20763 15351
rect 24685 15317 24719 15351
rect 29837 15317 29871 15351
rect 30481 15317 30515 15351
rect 38209 15317 38243 15351
rect 17141 15113 17175 15147
rect 25237 15113 25271 15147
rect 27813 15113 27847 15147
rect 29929 15113 29963 15147
rect 1869 15045 1903 15079
rect 7665 15045 7699 15079
rect 10241 15045 10275 15079
rect 11161 15045 11195 15079
rect 11989 15045 12023 15079
rect 13737 15045 13771 15079
rect 15393 15045 15427 15079
rect 17877 15045 17911 15079
rect 19533 15045 19567 15079
rect 20821 15045 20855 15079
rect 22201 15045 22235 15079
rect 23121 15045 23155 15079
rect 23673 15045 23707 15079
rect 23765 15045 23799 15079
rect 28733 15045 28767 15079
rect 28825 15045 28859 15079
rect 30573 15045 30607 15079
rect 1593 14977 1627 15011
rect 4261 14977 4295 15011
rect 6561 14967 6595 15001
rect 7389 14977 7423 15011
rect 9413 14977 9447 15011
rect 11713 14977 11747 15011
rect 14197 14977 14231 15011
rect 17049 14977 17083 15011
rect 21373 14977 21407 15011
rect 25145 14977 25179 15011
rect 25789 14977 25823 15011
rect 26433 14977 26467 15011
rect 27169 14977 27203 15011
rect 29837 14977 29871 15011
rect 30481 14977 30515 15011
rect 31125 14977 31159 15011
rect 38025 14977 38059 15011
rect 3617 14909 3651 14943
rect 4537 14909 4571 14943
rect 10149 14909 10183 14943
rect 14381 14909 14415 14943
rect 15301 14909 15335 14943
rect 15577 14909 15611 14943
rect 17785 14909 17819 14943
rect 18061 14909 18095 14943
rect 19441 14909 19475 14943
rect 19901 14909 19935 14943
rect 20729 14909 20763 14943
rect 22109 14909 22143 14943
rect 24593 14909 24627 14943
rect 29193 14909 29227 14943
rect 27261 14841 27295 14875
rect 3893 14773 3927 14807
rect 6009 14773 6043 14807
rect 6653 14773 6687 14807
rect 25881 14773 25915 14807
rect 26525 14773 26559 14807
rect 31217 14773 31251 14807
rect 37841 14773 37875 14807
rect 10964 14569 10998 14603
rect 22109 14569 22143 14603
rect 23765 14569 23799 14603
rect 27077 14569 27111 14603
rect 27721 14569 27755 14603
rect 37381 14569 37415 14603
rect 1685 14433 1719 14467
rect 1961 14433 1995 14467
rect 3985 14433 4019 14467
rect 6009 14433 6043 14467
rect 6561 14433 6595 14467
rect 9505 14433 9539 14467
rect 10701 14433 10735 14467
rect 12725 14433 12759 14467
rect 13369 14433 13403 14467
rect 16497 14433 16531 14467
rect 17877 14433 17911 14467
rect 20545 14433 20579 14467
rect 24685 14433 24719 14467
rect 28365 14433 28399 14467
rect 31125 14433 31159 14467
rect 31401 14433 31435 14467
rect 13185 14365 13219 14399
rect 19441 14365 19475 14399
rect 22017 14365 22051 14399
rect 23673 14365 23707 14399
rect 25329 14365 25363 14399
rect 26993 14367 27027 14401
rect 27629 14367 27663 14401
rect 28273 14365 28307 14399
rect 28917 14365 28951 14399
rect 30389 14365 30423 14399
rect 37565 14365 37599 14399
rect 38025 14365 38059 14399
rect 4261 14297 4295 14331
rect 6837 14297 6871 14331
rect 8585 14297 8619 14331
rect 9597 14297 9631 14331
rect 10149 14297 10183 14331
rect 14289 14297 14323 14331
rect 17601 14297 17635 14331
rect 17693 14297 17727 14331
rect 20646 14297 20680 14331
rect 21557 14297 21591 14331
rect 23029 14297 23063 14331
rect 24777 14297 24811 14331
rect 25881 14297 25915 14331
rect 25973 14297 26007 14331
rect 26525 14297 26559 14331
rect 29009 14297 29043 14331
rect 31217 14297 31251 14331
rect 3433 14229 3467 14263
rect 15577 14229 15611 14263
rect 19533 14229 19567 14263
rect 23121 14229 23155 14263
rect 29745 14229 29779 14263
rect 30481 14229 30515 14263
rect 38209 14229 38243 14263
rect 21189 14025 21223 14059
rect 26525 14025 26559 14059
rect 30757 14025 30791 14059
rect 38117 14025 38151 14059
rect 4537 13957 4571 13991
rect 5457 13957 5491 13991
rect 10609 13957 10643 13991
rect 11161 13957 11195 13991
rect 11989 13957 12023 13991
rect 14473 13957 14507 13991
rect 16957 13957 16991 13991
rect 17049 13957 17083 13991
rect 19533 13957 19567 13991
rect 19625 13957 19659 13991
rect 20545 13957 20579 13991
rect 22201 13957 22235 13991
rect 23397 13957 23431 13991
rect 25053 13957 25087 13991
rect 27905 13957 27939 13991
rect 29009 13957 29043 13991
rect 29101 13957 29135 13991
rect 1593 13889 1627 13923
rect 6009 13889 6043 13923
rect 6561 13889 6595 13923
rect 15853 13889 15887 13923
rect 18061 13889 18095 13923
rect 18153 13889 18187 13923
rect 18705 13889 18739 13923
rect 21097 13889 21131 13923
rect 26433 13889 26467 13923
rect 27169 13889 27203 13923
rect 27813 13889 27847 13923
rect 30665 13889 30699 13923
rect 38301 13889 38335 13923
rect 2513 13821 2547 13855
rect 2789 13821 2823 13855
rect 5365 13821 5399 13855
rect 7389 13821 7423 13855
rect 7665 13821 7699 13855
rect 9413 13821 9447 13855
rect 10517 13821 10551 13855
rect 11713 13821 11747 13855
rect 13737 13821 13771 13855
rect 14381 13821 14415 13855
rect 15209 13821 15243 13855
rect 16129 13821 16163 13855
rect 18797 13821 18831 13855
rect 22109 13821 22143 13855
rect 22477 13821 22511 13855
rect 23305 13821 23339 13855
rect 24961 13821 24995 13855
rect 25881 13821 25915 13855
rect 29377 13821 29411 13855
rect 17509 13753 17543 13787
rect 23857 13753 23891 13787
rect 1777 13685 1811 13719
rect 6745 13685 6779 13719
rect 27261 13685 27295 13719
rect 3433 13481 3467 13515
rect 21005 13481 21039 13515
rect 23213 13481 23247 13515
rect 23857 13481 23891 13515
rect 26433 13413 26467 13447
rect 27629 13413 27663 13447
rect 1685 13345 1719 13379
rect 4077 13345 4111 13379
rect 4353 13345 4387 13379
rect 8585 13345 8619 13379
rect 11989 13345 12023 13379
rect 13737 13345 13771 13379
rect 15393 13345 15427 13379
rect 16313 13345 16347 13379
rect 16681 13345 16715 13379
rect 21649 13345 21683 13379
rect 28273 13345 28307 13379
rect 6561 13277 6595 13311
rect 9229 13277 9263 13311
rect 11713 13277 11747 13311
rect 17417 13277 17451 13311
rect 17509 13277 17543 13311
rect 18889 13277 18923 13311
rect 20177 13277 20211 13311
rect 20913 13277 20947 13311
rect 23121 13277 23155 13311
rect 23765 13277 23799 13311
rect 24593 13277 24627 13311
rect 28181 13277 28215 13311
rect 28825 13277 28859 13311
rect 29745 13277 29779 13311
rect 1961 13209 1995 13243
rect 6101 13209 6135 13243
rect 6837 13209 6871 13243
rect 9505 13209 9539 13243
rect 11253 13209 11287 13243
rect 14381 13209 14415 13243
rect 14473 13209 14507 13243
rect 16405 13209 16439 13243
rect 18245 13209 18279 13243
rect 18337 13209 18371 13243
rect 19533 13209 19567 13243
rect 19625 13209 19659 13243
rect 21741 13209 21775 13243
rect 22661 13209 22695 13243
rect 24685 13209 24719 13243
rect 25881 13209 25915 13243
rect 25973 13209 26007 13243
rect 27077 13209 27111 13243
rect 27169 13209 27203 13243
rect 29837 13209 29871 13243
rect 28917 13141 28951 13175
rect 23305 12937 23339 12971
rect 23949 12937 23983 12971
rect 25237 12937 25271 12971
rect 32413 12937 32447 12971
rect 2421 12869 2455 12903
rect 4169 12869 4203 12903
rect 4813 12869 4847 12903
rect 6929 12869 6963 12903
rect 9413 12869 9447 12903
rect 14473 12869 14507 12903
rect 15393 12869 15427 12903
rect 17049 12869 17083 12903
rect 17141 12869 17175 12903
rect 18337 12869 18371 12903
rect 20177 12869 20211 12903
rect 21097 12869 21131 12903
rect 22109 12869 22143 12903
rect 22201 12869 22235 12903
rect 26065 12869 26099 12903
rect 27261 12869 27295 12903
rect 27997 12869 28031 12903
rect 30849 12869 30883 12903
rect 2145 12801 2179 12835
rect 8677 12801 8711 12835
rect 9137 12801 9171 12835
rect 15853 12801 15887 12835
rect 23213 12801 23247 12835
rect 23857 12801 23891 12835
rect 24501 12801 24535 12835
rect 25145 12801 25179 12835
rect 27169 12801 27203 12835
rect 32321 12801 32355 12835
rect 38025 12801 38059 12835
rect 4721 12733 4755 12767
rect 5733 12733 5767 12767
rect 6653 12733 6687 12767
rect 11161 12733 11195 12767
rect 11805 12733 11839 12767
rect 12081 12733 12115 12767
rect 13829 12733 13863 12767
rect 14381 12733 14415 12767
rect 16129 12733 16163 12767
rect 17509 12733 17543 12767
rect 18245 12733 18279 12767
rect 19073 12733 19107 12767
rect 20085 12733 20119 12767
rect 22753 12733 22787 12767
rect 25973 12733 26007 12767
rect 26617 12733 26651 12767
rect 27905 12733 27939 12767
rect 28181 12733 28215 12767
rect 30757 12733 30791 12767
rect 31677 12733 31711 12767
rect 24593 12665 24627 12699
rect 38209 12597 38243 12631
rect 1948 12393 1982 12427
rect 27445 12393 27479 12427
rect 34897 12393 34931 12427
rect 20637 12325 20671 12359
rect 21281 12325 21315 12359
rect 24685 12325 24719 12359
rect 28641 12325 28675 12359
rect 1685 12257 1719 12291
rect 5089 12257 5123 12291
rect 5733 12257 5767 12291
rect 9873 12257 9907 12291
rect 11253 12257 11287 12291
rect 11529 12257 11563 12291
rect 16865 12257 16899 12291
rect 20085 12257 20119 12291
rect 25881 12257 25915 12291
rect 26157 12257 26191 12291
rect 30941 12257 30975 12291
rect 7757 12189 7791 12223
rect 8585 12189 8619 12223
rect 10517 12189 10551 12223
rect 15669 12189 15703 12223
rect 17509 12189 17543 12223
rect 21189 12189 21223 12223
rect 23673 12189 23707 12223
rect 24593 12189 24627 12223
rect 27353 12189 27387 12223
rect 35081 12189 35115 12223
rect 4077 12121 4111 12155
rect 4169 12121 4203 12155
rect 6009 12121 6043 12155
rect 8401 12121 8435 12155
rect 9137 12121 9171 12155
rect 13277 12121 13311 12155
rect 14289 12121 14323 12155
rect 15025 12121 15059 12155
rect 16957 12121 16991 12155
rect 18061 12121 18095 12155
rect 18153 12121 18187 12155
rect 18705 12121 18739 12155
rect 20177 12121 20211 12155
rect 22201 12121 22235 12155
rect 22293 12121 22327 12155
rect 23213 12121 23247 12155
rect 25973 12121 26007 12155
rect 28457 12121 28491 12155
rect 3433 12053 3467 12087
rect 10609 12053 10643 12087
rect 15761 12053 15795 12087
rect 23765 12053 23799 12087
rect 3341 11849 3375 11883
rect 8493 11849 8527 11883
rect 8861 11849 8895 11883
rect 20361 11849 20395 11883
rect 21005 11849 21039 11883
rect 28825 11849 28859 11883
rect 34069 11849 34103 11883
rect 6009 11781 6043 11815
rect 9413 11781 9447 11815
rect 14565 11781 14599 11815
rect 15117 11781 15151 11815
rect 15761 11781 15795 11815
rect 16957 11781 16991 11815
rect 17049 11781 17083 11815
rect 18521 11781 18555 11815
rect 18613 11781 18647 11815
rect 19717 11781 19751 11815
rect 22109 11781 22143 11815
rect 22937 11781 22971 11815
rect 24317 11781 24351 11815
rect 24409 11781 24443 11815
rect 25881 11781 25915 11815
rect 25973 11781 26007 11815
rect 1593 11713 1627 11747
rect 6745 11713 6779 11747
rect 11161 11713 11195 11747
rect 11897 11713 11931 11747
rect 19625 11713 19659 11747
rect 20269 11713 20303 11747
rect 20913 11713 20947 11747
rect 22017 11713 22051 11747
rect 27169 11713 27203 11747
rect 27813 11713 27847 11747
rect 28733 11713 28767 11747
rect 33977 11713 34011 11747
rect 1869 11645 1903 11679
rect 3985 11645 4019 11679
rect 4261 11645 4295 11679
rect 7021 11645 7055 11679
rect 9137 11645 9171 11679
rect 12173 11645 12207 11679
rect 13921 11645 13955 11679
rect 14473 11645 14507 11679
rect 15669 11645 15703 11679
rect 17601 11645 17635 11679
rect 18797 11645 18831 11679
rect 22845 11645 22879 11679
rect 23121 11645 23155 11679
rect 24593 11645 24627 11679
rect 26249 11645 26283 11679
rect 37473 11645 37507 11679
rect 37749 11645 37783 11679
rect 16221 11577 16255 11611
rect 27261 11577 27295 11611
rect 27905 11509 27939 11543
rect 19533 11305 19567 11339
rect 21741 11305 21775 11339
rect 22385 11305 22419 11339
rect 25329 11305 25363 11339
rect 25973 11305 26007 11339
rect 26617 11305 26651 11339
rect 27261 11305 27295 11339
rect 3433 11237 3467 11271
rect 4077 11237 4111 11271
rect 13645 11237 13679 11271
rect 1685 11169 1719 11203
rect 1961 11169 1995 11203
rect 5549 11169 5583 11203
rect 9873 11169 9907 11203
rect 10885 11169 10919 11203
rect 14289 11169 14323 11203
rect 16037 11169 16071 11203
rect 16865 11169 16899 11203
rect 17141 11169 17175 11203
rect 21189 11169 21223 11203
rect 23397 11169 23431 11203
rect 23673 11169 23707 11203
rect 4905 11101 4939 11135
rect 8125 11101 8159 11135
rect 12909 11101 12943 11135
rect 13553 11101 13587 11135
rect 18705 11101 18739 11135
rect 19441 11101 19475 11135
rect 21649 11101 21683 11135
rect 22293 11101 22327 11135
rect 24777 11101 24811 11135
rect 25237 11101 25271 11135
rect 25881 11101 25915 11135
rect 26525 11101 26559 11135
rect 27169 11101 27203 11135
rect 27813 11101 27847 11135
rect 4169 11033 4203 11067
rect 5825 11033 5859 11067
rect 7573 11033 7607 11067
rect 8401 11033 8435 11067
rect 9137 11033 9171 11067
rect 11161 11033 11195 11067
rect 14565 11033 14599 11067
rect 16957 11033 16991 11067
rect 18061 11033 18095 11067
rect 18153 11033 18187 11067
rect 20177 11033 20211 11067
rect 20269 11033 20303 11067
rect 23489 11033 23523 11067
rect 24593 10965 24627 10999
rect 27905 10965 27939 10999
rect 22109 10761 22143 10795
rect 23397 10761 23431 10795
rect 24041 10761 24075 10795
rect 26157 10761 26191 10795
rect 1869 10693 1903 10727
rect 6009 10693 6043 10727
rect 6929 10693 6963 10727
rect 9413 10693 9447 10727
rect 12173 10693 12207 10727
rect 13921 10693 13955 10727
rect 14473 10693 14507 10727
rect 14565 10693 14599 10727
rect 15117 10693 15151 10727
rect 15669 10693 15703 10727
rect 15761 10693 15795 10727
rect 16313 10693 16347 10727
rect 16957 10693 16991 10727
rect 17049 10693 17083 10727
rect 19165 10693 19199 10727
rect 20913 10693 20947 10727
rect 25053 10693 25087 10727
rect 38301 10693 38335 10727
rect 1593 10625 1627 10659
rect 3985 10625 4019 10659
rect 8677 10625 8711 10659
rect 11897 10625 11931 10659
rect 20361 10625 20395 10659
rect 20813 10625 20847 10659
rect 22017 10625 22051 10659
rect 22661 10625 22695 10659
rect 23305 10625 23339 10659
rect 23949 10625 23983 10659
rect 26065 10625 26099 10659
rect 27169 10625 27203 10659
rect 38117 10625 38151 10659
rect 4261 10557 4295 10591
rect 6653 10557 6687 10591
rect 9137 10557 9171 10591
rect 11161 10557 11195 10591
rect 17233 10557 17267 10591
rect 19073 10557 19107 10591
rect 19717 10557 19751 10591
rect 22753 10557 22787 10591
rect 24961 10557 24995 10591
rect 25237 10557 25271 10591
rect 3341 10421 3375 10455
rect 3709 10421 3743 10455
rect 20177 10421 20211 10455
rect 27261 10421 27295 10455
rect 3433 10217 3467 10251
rect 4537 10217 4571 10251
rect 20821 10217 20855 10251
rect 21465 10217 21499 10251
rect 22753 10217 22787 10251
rect 24685 10217 24719 10251
rect 25329 10217 25363 10251
rect 32873 10217 32907 10251
rect 8493 10149 8527 10183
rect 23949 10149 23983 10183
rect 1685 10081 1719 10115
rect 1961 10081 1995 10115
rect 4077 10081 4111 10115
rect 5089 10081 5123 10115
rect 7113 10081 7147 10115
rect 9137 10081 9171 10115
rect 9413 10081 9447 10115
rect 15485 10081 15519 10115
rect 16957 10081 16991 10115
rect 22109 10081 22143 10115
rect 27077 10081 27111 10115
rect 27905 10081 27939 10115
rect 4353 10013 4387 10047
rect 11713 10013 11747 10047
rect 14473 10013 14507 10047
rect 18889 10013 18923 10047
rect 19533 10013 19567 10047
rect 20729 10013 20763 10047
rect 21373 10013 21407 10047
rect 22017 10013 22051 10047
rect 22661 10013 22695 10047
rect 24593 10013 24627 10047
rect 25237 10013 25271 10047
rect 25881 10013 25915 10047
rect 32781 10013 32815 10047
rect 37473 10013 37507 10047
rect 37749 10013 37783 10047
rect 5365 9945 5399 9979
rect 7941 9945 7975 9979
rect 8033 9945 8067 9979
rect 11161 9945 11195 9979
rect 11989 9945 12023 9979
rect 13737 9945 13771 9979
rect 14749 9945 14783 9979
rect 15577 9945 15611 9979
rect 16129 9945 16163 9979
rect 16681 9945 16715 9979
rect 16773 9945 16807 9979
rect 18245 9945 18279 9979
rect 18337 9945 18371 9979
rect 19717 9945 19751 9979
rect 23397 9945 23431 9979
rect 23489 9945 23523 9979
rect 27169 9945 27203 9979
rect 25973 9877 26007 9911
rect 26065 9673 26099 9707
rect 1869 9605 1903 9639
rect 8861 9605 8895 9639
rect 9689 9605 9723 9639
rect 13921 9605 13955 9639
rect 14565 9605 14599 9639
rect 15669 9605 15703 9639
rect 15761 9605 15795 9639
rect 16313 9605 16347 9639
rect 17406 9605 17440 9639
rect 17502 9605 17536 9639
rect 21373 9605 21407 9639
rect 22201 9605 22235 9639
rect 22753 9605 22787 9639
rect 23857 9605 23891 9639
rect 27905 9605 27939 9639
rect 1593 9537 1627 9571
rect 4077 9537 4111 9571
rect 8769 9537 8803 9571
rect 9413 9537 9447 9571
rect 15117 9537 15151 9571
rect 18521 9537 18555 9571
rect 19441 9537 19475 9571
rect 20637 9537 20671 9571
rect 20729 9537 20763 9571
rect 21281 9537 21315 9571
rect 24869 9537 24903 9571
rect 25973 9537 26007 9571
rect 27169 9537 27203 9571
rect 27813 9537 27847 9571
rect 3617 9469 3651 9503
rect 5825 9469 5859 9503
rect 6561 9469 6595 9503
rect 6837 9469 6871 9503
rect 11897 9469 11931 9503
rect 14473 9469 14507 9503
rect 17693 9469 17727 9503
rect 18705 9469 18739 9503
rect 19717 9469 19751 9503
rect 22109 9469 22143 9503
rect 23765 9469 23799 9503
rect 24317 9401 24351 9435
rect 4340 9333 4374 9367
rect 8309 9333 8343 9367
rect 11161 9333 11195 9367
rect 12160 9333 12194 9367
rect 24961 9333 24995 9367
rect 27261 9333 27295 9367
rect 10701 9129 10735 9163
rect 19533 9129 19567 9163
rect 21373 9129 21407 9163
rect 3341 9061 3375 9095
rect 8585 9061 8619 9095
rect 24685 9061 24719 9095
rect 3985 8993 4019 9027
rect 9229 8993 9263 9027
rect 9873 8993 9907 9027
rect 11253 8993 11287 9027
rect 13277 8993 13311 9027
rect 16313 8993 16347 9027
rect 17325 8993 17359 9027
rect 18797 8993 18831 9027
rect 22845 8993 22879 9027
rect 27537 8993 27571 9027
rect 1593 8925 1627 8959
rect 6837 8925 6871 8959
rect 10609 8925 10643 8959
rect 19441 8925 19475 8959
rect 21281 8925 21315 8959
rect 23673 8925 23707 8959
rect 24593 8925 24627 8959
rect 25513 8925 25547 8959
rect 38025 8925 38059 8959
rect 1869 8857 1903 8891
rect 4261 8857 4295 8891
rect 6009 8857 6043 8891
rect 7113 8857 7147 8891
rect 9321 8857 9355 8891
rect 11529 8857 11563 8891
rect 14277 8857 14311 8891
rect 15117 8857 15151 8891
rect 16405 8857 16439 8891
rect 17877 8857 17911 8891
rect 17969 8857 18003 8891
rect 20177 8857 20211 8891
rect 20269 8857 20303 8891
rect 20821 8857 20855 8891
rect 22569 8857 22603 8891
rect 22661 8857 22695 8891
rect 27261 8857 27295 8891
rect 27353 8857 27387 8891
rect 23765 8789 23799 8823
rect 25605 8789 25639 8823
rect 38209 8789 38243 8823
rect 6009 8585 6043 8619
rect 20085 8585 20119 8619
rect 21097 8585 21131 8619
rect 25145 8585 25179 8619
rect 29009 8585 29043 8619
rect 9413 8517 9447 8551
rect 15393 8517 15427 8551
rect 16946 8517 16980 8551
rect 17049 8517 17083 8551
rect 18245 8517 18279 8551
rect 18337 8517 18371 8551
rect 22486 8517 22520 8551
rect 23949 8517 23983 8551
rect 4261 8449 4295 8483
rect 9137 8449 9171 8483
rect 14381 8449 14415 8483
rect 19993 8449 20027 8483
rect 21005 8449 21039 8483
rect 23857 8449 23891 8483
rect 24501 8449 24535 8483
rect 25053 8449 25087 8483
rect 25513 8449 25547 8483
rect 26065 8449 26099 8483
rect 28917 8449 28951 8483
rect 1593 8381 1627 8415
rect 1869 8381 1903 8415
rect 3617 8381 3651 8415
rect 4537 8381 4571 8415
rect 6929 8381 6963 8415
rect 7205 8381 7239 8415
rect 11161 8381 11195 8415
rect 11713 8381 11747 8415
rect 11989 8381 12023 8415
rect 13737 8381 13771 8415
rect 15301 8381 15335 8415
rect 16313 8381 16347 8415
rect 19257 8381 19291 8415
rect 22385 8381 22419 8415
rect 23397 8381 23431 8415
rect 8677 8313 8711 8347
rect 17509 8313 17543 8347
rect 24593 8313 24627 8347
rect 25881 8313 25915 8347
rect 14657 8245 14691 8279
rect 3341 8041 3375 8075
rect 8493 8041 8527 8075
rect 11884 8041 11918 8075
rect 16037 8041 16071 8075
rect 21465 8041 21499 8075
rect 23397 8041 23431 8075
rect 26249 8041 26283 8075
rect 38117 8041 38151 8075
rect 11161 7973 11195 8007
rect 1869 7905 1903 7939
rect 4721 7905 4755 7939
rect 5825 7905 5859 7939
rect 7573 7905 7607 7939
rect 16589 7905 16623 7939
rect 17601 7905 17635 7939
rect 18429 7905 18463 7939
rect 19533 7905 19567 7939
rect 20453 7905 20487 7939
rect 22753 7905 22787 7939
rect 24961 7905 24995 7939
rect 1593 7837 1627 7871
rect 3985 7837 4019 7871
rect 5549 7837 5583 7871
rect 8401 7837 8435 7871
rect 9413 7837 9447 7871
rect 11621 7837 11655 7871
rect 14289 7837 14323 7871
rect 19441 7837 19475 7871
rect 20361 7837 20395 7871
rect 21373 7837 21407 7871
rect 22017 7837 22051 7871
rect 22661 7837 22695 7871
rect 23305 7837 23339 7871
rect 26157 7837 26191 7871
rect 38301 7837 38335 7871
rect 9689 7769 9723 7803
rect 13645 7769 13679 7803
rect 14565 7769 14599 7803
rect 16681 7769 16715 7803
rect 18153 7769 18187 7803
rect 18245 7769 18279 7803
rect 24685 7769 24719 7803
rect 24777 7769 24811 7803
rect 22109 7701 22143 7735
rect 1777 7497 1811 7531
rect 5089 7497 5123 7531
rect 16221 7497 16255 7531
rect 22109 7497 22143 7531
rect 23397 7497 23431 7531
rect 24501 7497 24535 7531
rect 24869 7497 24903 7531
rect 25237 7497 25271 7531
rect 38209 7497 38243 7531
rect 4997 7429 5031 7463
rect 5917 7429 5951 7463
rect 6837 7429 6871 7463
rect 7941 7429 7975 7463
rect 10149 7429 10183 7463
rect 17049 7429 17083 7463
rect 19533 7429 19567 7463
rect 20913 7429 20947 7463
rect 24041 7429 24075 7463
rect 1593 7361 1627 7395
rect 5825 7361 5859 7395
rect 6745 7361 6779 7395
rect 9689 7361 9723 7395
rect 13921 7361 13955 7395
rect 16129 7361 16163 7395
rect 18797 7361 18831 7395
rect 19441 7361 19475 7395
rect 20085 7361 20119 7395
rect 22017 7361 22051 7395
rect 22661 7361 22695 7395
rect 23305 7361 23339 7395
rect 23949 7361 23983 7395
rect 24409 7361 24443 7395
rect 38117 7361 38151 7395
rect 2421 7293 2455 7327
rect 2697 7293 2731 7327
rect 4445 7293 4479 7327
rect 7665 7293 7699 7327
rect 10885 7293 10919 7327
rect 11713 7293 11747 7327
rect 11989 7293 12023 7327
rect 14197 7293 14231 7327
rect 16957 7293 16991 7327
rect 17969 7293 18003 7327
rect 18889 7293 18923 7327
rect 20821 7293 20855 7327
rect 13461 7225 13495 7259
rect 20177 7225 20211 7259
rect 21373 7225 21407 7259
rect 15669 7157 15703 7191
rect 22753 7157 22787 7191
rect 1948 6953 1982 6987
rect 18797 6953 18831 6987
rect 6285 6885 6319 6919
rect 1685 6817 1719 6851
rect 3433 6817 3467 6851
rect 4537 6817 4571 6851
rect 17509 6817 17543 6851
rect 20177 6817 20211 6851
rect 20821 6817 20855 6851
rect 21465 6817 21499 6851
rect 23397 6817 23431 6851
rect 24685 6817 24719 6851
rect 27905 6817 27939 6851
rect 33057 6817 33091 6851
rect 6745 6749 6779 6783
rect 9597 6749 9631 6783
rect 9689 6749 9723 6783
rect 10425 6749 10459 6783
rect 12449 6749 12483 6783
rect 13277 6749 13311 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 15117 6749 15151 6783
rect 18705 6749 18739 6783
rect 19441 6749 19475 6783
rect 20085 6749 20119 6783
rect 20729 6749 20763 6783
rect 21373 6749 21407 6783
rect 22017 6749 22051 6783
rect 22661 6749 22695 6783
rect 23305 6749 23339 6783
rect 24593 6749 24627 6783
rect 25881 6749 25915 6783
rect 27813 6749 27847 6783
rect 32965 6749 32999 6783
rect 4813 6681 4847 6715
rect 7021 6681 7055 6715
rect 10701 6681 10735 6715
rect 13553 6681 13587 6715
rect 15393 6681 15427 6715
rect 16681 6681 16715 6715
rect 16773 6681 16807 6715
rect 8493 6613 8527 6647
rect 19533 6613 19567 6647
rect 22109 6613 22143 6647
rect 22753 6613 22787 6647
rect 25973 6613 26007 6647
rect 5917 6409 5951 6443
rect 9873 6409 9907 6443
rect 10701 6409 10735 6443
rect 22293 6409 22327 6443
rect 23581 6409 23615 6443
rect 23949 6409 23983 6443
rect 2329 6341 2363 6375
rect 4077 6341 4111 6375
rect 6561 6341 6595 6375
rect 7297 6341 7331 6375
rect 11989 6341 12023 6375
rect 14197 6341 14231 6375
rect 15117 6341 15151 6375
rect 17049 6341 17083 6375
rect 20085 6341 20119 6375
rect 21925 6341 21959 6375
rect 2053 6273 2087 6307
rect 4537 6273 4571 6307
rect 5825 6273 5859 6307
rect 8125 6273 8159 6307
rect 10609 6273 10643 6307
rect 11713 6273 11747 6307
rect 15669 6273 15703 6307
rect 17601 6273 17635 6307
rect 18429 6273 18463 6307
rect 19349 6273 19383 6307
rect 19441 6273 19475 6307
rect 19993 6273 20027 6307
rect 20637 6273 20671 6307
rect 21281 6273 21315 6307
rect 21833 6273 21867 6307
rect 22845 6273 22879 6307
rect 23305 6273 23339 6307
rect 24133 6273 24167 6307
rect 32321 6273 32355 6307
rect 8401 6205 8435 6239
rect 14105 6205 14139 6239
rect 15853 6205 15887 6239
rect 16957 6205 16991 6239
rect 20729 6205 20763 6239
rect 4721 6137 4755 6171
rect 13461 6137 13495 6171
rect 21373 6137 21407 6171
rect 18521 6069 18555 6103
rect 22661 6069 22695 6103
rect 23121 6069 23155 6103
rect 32413 6069 32447 6103
rect 1856 5865 1890 5899
rect 3341 5865 3375 5899
rect 9229 5865 9263 5899
rect 10057 5865 10091 5899
rect 16957 5865 16991 5899
rect 18153 5865 18187 5899
rect 18797 5865 18831 5899
rect 20085 5865 20119 5899
rect 21465 5865 21499 5899
rect 37657 5865 37691 5899
rect 5733 5797 5767 5831
rect 8033 5797 8067 5831
rect 12357 5797 12391 5831
rect 14381 5797 14415 5831
rect 1593 5729 1627 5763
rect 4261 5729 4295 5763
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 13093 5729 13127 5763
rect 3985 5661 4019 5695
rect 9137 5661 9171 5695
rect 9965 5661 9999 5695
rect 10977 5661 11011 5695
rect 11069 5661 11103 5695
rect 11621 5661 11655 5695
rect 12265 5661 12299 5695
rect 12909 5661 12943 5695
rect 14289 5661 14323 5695
rect 16865 5661 16899 5695
rect 18061 5661 18095 5695
rect 18705 5661 18739 5695
rect 19993 5661 20027 5695
rect 20721 5661 20755 5695
rect 20821 5661 20855 5695
rect 21373 5661 21407 5695
rect 22201 5661 22235 5695
rect 22661 5661 22695 5695
rect 23305 5661 23339 5695
rect 37381 5661 37415 5695
rect 38025 5661 38059 5695
rect 15025 5593 15059 5627
rect 15117 5593 15151 5627
rect 16037 5593 16071 5627
rect 22753 5593 22787 5627
rect 11713 5525 11747 5559
rect 22017 5525 22051 5559
rect 23397 5525 23431 5559
rect 37197 5525 37231 5559
rect 38209 5525 38243 5559
rect 6009 5321 6043 5355
rect 8861 5321 8895 5355
rect 9505 5321 9539 5355
rect 11069 5321 11103 5355
rect 13001 5321 13035 5355
rect 14289 5321 14323 5355
rect 14933 5321 14967 5355
rect 16221 5321 16255 5355
rect 19441 5321 19475 5355
rect 2329 5253 2363 5287
rect 6837 5253 6871 5287
rect 12357 5253 12391 5287
rect 13645 5253 13679 5287
rect 18797 5253 18831 5287
rect 21925 5253 21959 5287
rect 2053 5185 2087 5219
rect 8769 5185 8803 5219
rect 9405 5183 9439 5217
rect 10333 5185 10367 5219
rect 10977 5185 11011 5219
rect 12265 5185 12299 5219
rect 12909 5185 12943 5219
rect 13553 5185 13587 5219
rect 14197 5185 14231 5219
rect 14841 5185 14875 5219
rect 15485 5185 15519 5219
rect 16129 5185 16163 5219
rect 17417 5185 17451 5219
rect 18061 5185 18095 5219
rect 18153 5185 18187 5219
rect 18705 5185 18739 5219
rect 19349 5185 19383 5219
rect 20085 5185 20119 5219
rect 20729 5185 20763 5219
rect 21833 5185 21867 5219
rect 22845 5185 22879 5219
rect 23305 5185 23339 5219
rect 38025 5185 38059 5219
rect 4261 5117 4295 5151
rect 4537 5117 4571 5151
rect 6561 5117 6595 5151
rect 17509 5117 17543 5151
rect 23397 5117 23431 5151
rect 15577 5049 15611 5083
rect 20177 5049 20211 5083
rect 22661 5049 22695 5083
rect 3801 4981 3835 5015
rect 8309 4981 8343 5015
rect 10425 4981 10459 5015
rect 20821 4981 20855 5015
rect 22293 4981 22327 5015
rect 38209 4981 38243 5015
rect 7849 4777 7883 4811
rect 8493 4777 8527 4811
rect 9229 4777 9263 4811
rect 10425 4777 10459 4811
rect 11713 4777 11747 4811
rect 13001 4777 13035 4811
rect 14657 4777 14691 4811
rect 17877 4777 17911 4811
rect 20821 4777 20855 4811
rect 22109 4777 22143 4811
rect 3433 4709 3467 4743
rect 4905 4709 4939 4743
rect 7297 4709 7331 4743
rect 11069 4709 11103 4743
rect 13645 4709 13679 4743
rect 16589 4709 16623 4743
rect 17233 4709 17267 4743
rect 18521 4709 18555 4743
rect 1685 4641 1719 4675
rect 1961 4641 1995 4675
rect 15301 4641 15335 4675
rect 21373 4641 21407 4675
rect 3801 4573 3835 4607
rect 4721 4573 4755 4607
rect 5273 4573 5307 4607
rect 5549 4573 5583 4607
rect 7757 4573 7791 4607
rect 8401 4573 8435 4607
rect 9137 4573 9171 4607
rect 10333 4573 10367 4607
rect 10977 4573 11011 4607
rect 11621 4573 11655 4607
rect 12265 4573 12299 4607
rect 12909 4573 12943 4607
rect 13553 4573 13587 4607
rect 14565 4573 14599 4607
rect 15209 4573 15243 4607
rect 15853 4573 15887 4607
rect 16497 4573 16531 4607
rect 17141 4573 17175 4607
rect 17785 4573 17819 4607
rect 18429 4573 18463 4607
rect 19441 4573 19475 4607
rect 20085 4573 20119 4607
rect 20729 4573 20763 4607
rect 22017 4573 22051 4607
rect 22661 4573 22695 4607
rect 23305 4573 23339 4607
rect 31309 4573 31343 4607
rect 38025 4573 38059 4607
rect 5825 4505 5859 4539
rect 12357 4505 12391 4539
rect 15945 4505 15979 4539
rect 19533 4505 19567 4539
rect 20177 4505 20211 4539
rect 3985 4437 4019 4471
rect 4445 4437 4479 4471
rect 22753 4437 22787 4471
rect 23397 4437 23431 4471
rect 31125 4437 31159 4471
rect 38209 4437 38243 4471
rect 2421 4233 2455 4267
rect 9137 4233 9171 4267
rect 1685 4165 1719 4199
rect 3065 4165 3099 4199
rect 3985 4165 4019 4199
rect 23397 4165 23431 4199
rect 1869 4097 1903 4131
rect 2329 4097 2363 4131
rect 6561 4097 6595 4131
rect 7757 4097 7791 4131
rect 8401 4097 8435 4131
rect 9045 4097 9079 4131
rect 9689 4097 9723 4131
rect 10333 4097 10367 4131
rect 10977 4097 11011 4131
rect 11069 4097 11103 4131
rect 12265 4097 12299 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 13553 4097 13587 4131
rect 14197 4097 14231 4131
rect 14289 4097 14323 4131
rect 14841 4097 14875 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 16129 4097 16163 4131
rect 16865 4097 16899 4131
rect 17509 4097 17543 4131
rect 18153 4097 18187 4131
rect 18797 4097 18831 4131
rect 19441 4097 19475 4131
rect 19533 4097 19567 4131
rect 20269 4097 20303 4131
rect 20913 4097 20947 4131
rect 22017 4097 22051 4131
rect 22661 4097 22695 4131
rect 23305 4097 23339 4131
rect 24133 4097 24167 4131
rect 38025 4097 38059 4131
rect 3709 4029 3743 4063
rect 22109 4029 22143 4063
rect 3249 3961 3283 3995
rect 6745 3961 6779 3995
rect 8493 3961 8527 3995
rect 10425 3961 10459 3995
rect 12357 3961 12391 3995
rect 16221 3961 16255 3995
rect 17601 3961 17635 3995
rect 18889 3961 18923 3995
rect 20085 3961 20119 3995
rect 5457 3893 5491 3927
rect 7849 3893 7883 3927
rect 9781 3893 9815 3927
rect 13645 3893 13679 3927
rect 14933 3893 14967 3927
rect 16957 3893 16991 3927
rect 18245 3893 18279 3927
rect 20729 3893 20763 3927
rect 22753 3893 22787 3927
rect 23949 3893 23983 3927
rect 38209 3893 38243 3927
rect 6745 3689 6779 3723
rect 8493 3689 8527 3723
rect 10425 3689 10459 3723
rect 11713 3689 11747 3723
rect 12357 3689 12391 3723
rect 13645 3689 13679 3723
rect 16129 3689 16163 3723
rect 18061 3689 18095 3723
rect 18797 3689 18831 3723
rect 20821 3689 20855 3723
rect 24593 3689 24627 3723
rect 36737 3689 36771 3723
rect 9781 3621 9815 3655
rect 11069 3621 11103 3655
rect 20085 3621 20119 3655
rect 37381 3621 37415 3655
rect 1685 3553 1719 3587
rect 1961 3553 1995 3587
rect 4353 3553 4387 3587
rect 17325 3553 17359 3587
rect 38301 3553 38335 3587
rect 6561 3485 6595 3519
rect 7297 3485 7331 3519
rect 8401 3485 8435 3519
rect 9689 3485 9723 3519
rect 10333 3485 10367 3519
rect 10977 3485 11011 3519
rect 11621 3485 11655 3519
rect 12257 3485 12291 3519
rect 12909 3485 12943 3519
rect 13553 3485 13587 3519
rect 14749 3485 14783 3519
rect 14841 3485 14875 3519
rect 15393 3485 15427 3519
rect 16037 3485 16071 3519
rect 16681 3485 16715 3519
rect 17969 3485 18003 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 20729 3485 20763 3519
rect 21373 3485 21407 3519
rect 22017 3485 22051 3519
rect 22845 3485 22879 3519
rect 24041 3485 24075 3519
rect 24777 3485 24811 3519
rect 36921 3485 36955 3519
rect 37565 3485 37599 3519
rect 4629 3417 4663 3451
rect 16773 3417 16807 3451
rect 38117 3417 38151 3451
rect 3433 3349 3467 3383
rect 6101 3349 6135 3383
rect 7481 3349 7515 3383
rect 13001 3349 13035 3383
rect 15485 3349 15519 3383
rect 19533 3349 19567 3383
rect 21465 3349 21499 3383
rect 21833 3349 21867 3383
rect 22293 3349 22327 3383
rect 22661 3349 22695 3383
rect 23857 3349 23891 3383
rect 3341 3145 3375 3179
rect 6745 3145 6779 3179
rect 9873 3145 9907 3179
rect 12909 3145 12943 3179
rect 13553 3145 13587 3179
rect 15485 3145 15519 3179
rect 18153 3145 18187 3179
rect 19625 3145 19659 3179
rect 22017 3145 22051 3179
rect 25789 3145 25823 3179
rect 27813 3145 27847 3179
rect 32965 3145 32999 3179
rect 36737 3145 36771 3179
rect 1869 3077 1903 3111
rect 9229 3077 9263 3111
rect 10701 3077 10735 3111
rect 24961 3077 24995 3111
rect 1593 3009 1627 3043
rect 3801 3009 3835 3043
rect 6561 3009 6595 3043
rect 7297 3009 7331 3043
rect 8033 3009 8067 3043
rect 9137 3009 9171 3043
rect 9781 3009 9815 3043
rect 10517 3009 10551 3043
rect 11713 3009 11747 3043
rect 12817 3009 12851 3043
rect 13461 3009 13495 3043
rect 14105 3009 14139 3043
rect 14749 3009 14783 3043
rect 15393 3009 15427 3043
rect 16129 3009 16163 3043
rect 16313 3009 16347 3043
rect 16865 3009 16899 3043
rect 18337 3009 18371 3043
rect 18981 3009 19015 3043
rect 19441 3009 19475 3043
rect 20361 3009 20395 3043
rect 21005 3009 21039 3043
rect 22201 3009 22235 3043
rect 22845 3009 22879 3043
rect 23489 3009 23523 3043
rect 23949 3009 23983 3043
rect 25421 3009 25455 3043
rect 25973 3009 26007 3043
rect 26617 3009 26651 3043
rect 27997 3009 28031 3043
rect 33149 3009 33183 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 4077 2941 4111 2975
rect 7481 2873 7515 2907
rect 14841 2873 14875 2907
rect 18797 2873 18831 2907
rect 20177 2873 20211 2907
rect 20821 2873 20855 2907
rect 26433 2873 26467 2907
rect 5549 2805 5583 2839
rect 8217 2805 8251 2839
rect 11897 2805 11931 2839
rect 14197 2805 14231 2839
rect 17049 2805 17083 2839
rect 22661 2805 22695 2839
rect 23305 2805 23339 2839
rect 24133 2805 24167 2839
rect 25053 2805 25087 2839
rect 38209 2805 38243 2839
rect 3341 2601 3375 2635
rect 16865 2601 16899 2635
rect 19441 2601 19475 2635
rect 25881 2601 25915 2635
rect 35081 2601 35115 2635
rect 4629 2533 4663 2567
rect 5273 2533 5307 2567
rect 22293 2533 22327 2567
rect 27445 2533 27479 2567
rect 30757 2533 30791 2567
rect 35909 2533 35943 2567
rect 1593 2465 1627 2499
rect 1869 2465 1903 2499
rect 17785 2465 17819 2499
rect 20361 2465 20395 2499
rect 3985 2397 4019 2431
rect 5733 2397 5767 2431
rect 7205 2397 7239 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 9229 2397 9263 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 11713 2397 11747 2431
rect 12357 2397 12391 2431
rect 13553 2397 13587 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 15209 2397 15243 2431
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 23305 2397 23339 2431
rect 24593 2397 24627 2431
rect 24869 2397 24903 2431
rect 26065 2397 26099 2431
rect 28457 2397 28491 2431
rect 29929 2397 29963 2431
rect 30297 2397 30331 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 37749 2397 37783 2431
rect 5089 2329 5123 2363
rect 11805 2329 11839 2363
rect 22109 2329 22143 2363
rect 27261 2329 27295 2363
rect 34989 2329 35023 2363
rect 35725 2329 35759 2363
rect 4169 2261 4203 2295
rect 5917 2261 5951 2295
rect 6561 2261 6595 2295
rect 7389 2261 7423 2295
rect 8125 2261 8159 2295
rect 12541 2261 12575 2295
rect 13645 2261 13679 2295
rect 14381 2261 14415 2295
rect 23489 2261 23523 2295
rect 28641 2261 28675 2295
rect 29745 2261 29779 2295
rect 30389 2261 30423 2295
rect 31309 2261 31343 2295
rect 32505 2261 32539 2295
rect 33793 2261 33827 2295
rect 36829 2261 36863 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 2133 37451 2191 37457
rect 2133 37417 2145 37451
rect 2179 37448 2191 37451
rect 16758 37448 16764 37460
rect 2179 37420 16764 37448
rect 2179 37417 2191 37420
rect 2133 37411 2191 37417
rect 16758 37408 16764 37420
rect 16816 37408 16822 37460
rect 17037 37451 17095 37457
rect 17037 37417 17049 37451
rect 17083 37448 17095 37451
rect 22738 37448 22744 37460
rect 17083 37420 22744 37448
rect 17083 37417 17095 37420
rect 17037 37411 17095 37417
rect 22738 37408 22744 37420
rect 22796 37408 22802 37460
rect 32214 37408 32220 37460
rect 32272 37448 32278 37460
rect 33229 37451 33287 37457
rect 33229 37448 33241 37451
rect 32272 37420 33241 37448
rect 32272 37408 32278 37420
rect 33229 37417 33241 37420
rect 33275 37417 33287 37451
rect 33229 37411 33287 37417
rect 6825 37383 6883 37389
rect 6825 37349 6837 37383
rect 6871 37380 6883 37383
rect 20162 37380 20168 37392
rect 6871 37352 20168 37380
rect 6871 37349 6883 37352
rect 6825 37343 6883 37349
rect 20162 37340 20168 37352
rect 20220 37340 20226 37392
rect 2866 37272 2872 37324
rect 2924 37312 2930 37324
rect 10318 37312 10324 37324
rect 2924 37284 4200 37312
rect 10279 37284 10324 37312
rect 2924 37272 2930 37284
rect 1946 37204 1952 37256
rect 2004 37244 2010 37256
rect 2041 37247 2099 37253
rect 2041 37244 2053 37247
rect 2004 37216 2053 37244
rect 2004 37204 2010 37216
rect 2041 37213 2053 37216
rect 2087 37213 2099 37247
rect 2041 37207 2099 37213
rect 2685 37247 2743 37253
rect 2685 37213 2697 37247
rect 2731 37244 2743 37247
rect 2958 37244 2964 37256
rect 2731 37216 2964 37244
rect 2731 37213 2743 37216
rect 2685 37207 2743 37213
rect 2958 37204 2964 37216
rect 3016 37204 3022 37256
rect 4172 37253 4200 37284
rect 10318 37272 10324 37284
rect 10376 37272 10382 37324
rect 14826 37272 14832 37324
rect 14884 37312 14890 37324
rect 14921 37315 14979 37321
rect 14921 37312 14933 37315
rect 14884 37284 14933 37312
rect 14884 37272 14890 37284
rect 14921 37281 14933 37284
rect 14967 37281 14979 37315
rect 20622 37312 20628 37324
rect 20583 37284 20628 37312
rect 14921 37275 14979 37281
rect 20622 37272 20628 37284
rect 20680 37272 20686 37324
rect 22554 37272 22560 37324
rect 22612 37312 22618 37324
rect 22649 37315 22707 37321
rect 22649 37312 22661 37315
rect 22612 37284 22661 37312
rect 22612 37272 22618 37284
rect 22649 37281 22661 37284
rect 22695 37281 22707 37315
rect 30926 37312 30932 37324
rect 30887 37284 30932 37312
rect 22649 37275 22707 37281
rect 30926 37272 30932 37284
rect 30984 37272 30990 37324
rect 34146 37272 34152 37324
rect 34204 37312 34210 37324
rect 34885 37315 34943 37321
rect 34885 37312 34897 37315
rect 34204 37284 34897 37312
rect 34204 37272 34210 37284
rect 34885 37281 34897 37284
rect 34931 37281 34943 37315
rect 34885 37275 34943 37281
rect 4157 37247 4215 37253
rect 4157 37213 4169 37247
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4617 37247 4675 37253
rect 4617 37213 4629 37247
rect 4663 37244 4675 37247
rect 5718 37244 5724 37256
rect 4663 37216 5724 37244
rect 4663 37213 4675 37216
rect 4617 37207 4675 37213
rect 5718 37204 5724 37216
rect 5776 37204 5782 37256
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 6641 37247 6699 37253
rect 6641 37244 6653 37247
rect 5868 37216 6653 37244
rect 5868 37204 5874 37216
rect 6641 37213 6653 37216
rect 6687 37213 6699 37247
rect 6641 37207 6699 37213
rect 7098 37204 7104 37256
rect 7156 37244 7162 37256
rect 7469 37247 7527 37253
rect 7469 37244 7481 37247
rect 7156 37216 7481 37244
rect 7156 37204 7162 37216
rect 7469 37213 7481 37216
rect 7515 37213 7527 37247
rect 9122 37244 9128 37256
rect 9083 37216 9128 37244
rect 7469 37207 7527 37213
rect 9122 37204 9128 37216
rect 9180 37204 9186 37256
rect 10594 37244 10600 37256
rect 10555 37216 10600 37244
rect 10594 37204 10600 37216
rect 10652 37204 10658 37256
rect 11701 37247 11759 37253
rect 11701 37213 11713 37247
rect 11747 37213 11759 37247
rect 12986 37244 12992 37256
rect 12947 37216 12992 37244
rect 11701 37207 11759 37213
rect 6822 37176 6828 37188
rect 3988 37148 6828 37176
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 3988 37117 4016 37148
rect 6822 37136 6828 37148
rect 6880 37136 6886 37188
rect 10778 37176 10784 37188
rect 7300 37148 10784 37176
rect 2869 37111 2927 37117
rect 2869 37108 2881 37111
rect 2832 37080 2881 37108
rect 2832 37068 2838 37080
rect 2869 37077 2881 37080
rect 2915 37077 2927 37111
rect 2869 37071 2927 37077
rect 3973 37111 4031 37117
rect 3973 37077 3985 37111
rect 4019 37077 4031 37111
rect 3973 37071 4031 37077
rect 4614 37068 4620 37120
rect 4672 37108 4678 37120
rect 7300 37117 7328 37148
rect 10778 37136 10784 37148
rect 10836 37136 10842 37188
rect 11716 37176 11744 37207
rect 12986 37204 12992 37216
rect 13044 37204 13050 37256
rect 13538 37204 13544 37256
rect 13596 37244 13602 37256
rect 14461 37247 14519 37253
rect 14461 37244 14473 37247
rect 13596 37216 14473 37244
rect 13596 37204 13602 37216
rect 14461 37213 14473 37216
rect 14507 37213 14519 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 14461 37207 14519 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 18046 37204 18052 37256
rect 18104 37244 18110 37256
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18104 37216 18337 37244
rect 18104 37204 18110 37216
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 19889 37247 19947 37253
rect 19889 37213 19901 37247
rect 19935 37244 19947 37247
rect 20070 37244 20076 37256
rect 19935 37216 20076 37244
rect 19935 37213 19947 37216
rect 19889 37207 19947 37213
rect 20070 37204 20076 37216
rect 20128 37204 20134 37256
rect 20898 37244 20904 37256
rect 20859 37216 20904 37244
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 22925 37247 22983 37253
rect 22925 37213 22937 37247
rect 22971 37213 22983 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 22925 37207 22983 37213
rect 16114 37176 16120 37188
rect 11716 37148 16120 37176
rect 16114 37136 16120 37148
rect 16172 37136 16178 37188
rect 16574 37136 16580 37188
rect 16632 37176 16638 37188
rect 16945 37179 17003 37185
rect 16945 37176 16957 37179
rect 16632 37148 16957 37176
rect 16632 37136 16638 37148
rect 16945 37145 16957 37148
rect 16991 37145 17003 37179
rect 22940 37176 22968 37207
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 25314 37244 25320 37256
rect 25275 37216 25320 37244
rect 25314 37204 25320 37216
rect 25372 37204 25378 37256
rect 26234 37204 26240 37256
rect 26292 37244 26298 37256
rect 27157 37247 27215 37253
rect 27157 37244 27169 37247
rect 26292 37216 27169 37244
rect 26292 37204 26298 37216
rect 27157 37213 27169 37216
rect 27203 37213 27215 37247
rect 27157 37207 27215 37213
rect 27522 37204 27528 37256
rect 27580 37244 27586 37256
rect 27893 37247 27951 37253
rect 27893 37244 27905 37247
rect 27580 37216 27905 37244
rect 27580 37204 27586 37216
rect 27893 37213 27905 37216
rect 27939 37213 27951 37247
rect 27893 37207 27951 37213
rect 28813 37247 28871 37253
rect 28813 37213 28825 37247
rect 28859 37213 28871 37247
rect 29730 37244 29736 37256
rect 29691 37216 29736 37244
rect 28813 37207 28871 37213
rect 26970 37176 26976 37188
rect 22940 37148 26976 37176
rect 16945 37139 17003 37145
rect 26970 37136 26976 37148
rect 27028 37136 27034 37188
rect 27062 37136 27068 37188
rect 27120 37176 27126 37188
rect 27120 37148 27660 37176
rect 27120 37136 27126 37148
rect 4801 37111 4859 37117
rect 4801 37108 4813 37111
rect 4672 37080 4813 37108
rect 4672 37068 4678 37080
rect 4801 37077 4813 37080
rect 4847 37077 4859 37111
rect 4801 37071 4859 37077
rect 7285 37111 7343 37117
rect 7285 37077 7297 37111
rect 7331 37077 7343 37111
rect 7285 37071 7343 37077
rect 8386 37068 8392 37120
rect 8444 37108 8450 37120
rect 9309 37111 9367 37117
rect 9309 37108 9321 37111
rect 8444 37080 9321 37108
rect 8444 37068 8450 37080
rect 9309 37077 9321 37080
rect 9355 37077 9367 37111
rect 9309 37071 9367 37077
rect 11606 37068 11612 37120
rect 11664 37108 11670 37120
rect 11885 37111 11943 37117
rect 11885 37108 11897 37111
rect 11664 37080 11897 37108
rect 11664 37068 11670 37080
rect 11885 37077 11897 37080
rect 11931 37077 11943 37111
rect 11885 37071 11943 37077
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 13173 37111 13231 37117
rect 13173 37108 13185 37111
rect 12952 37080 13185 37108
rect 12952 37068 12958 37080
rect 13173 37077 13185 37080
rect 13219 37077 13231 37111
rect 13173 37071 13231 37077
rect 14277 37111 14335 37117
rect 14277 37077 14289 37111
rect 14323 37108 14335 37111
rect 15010 37108 15016 37120
rect 14323 37080 15016 37108
rect 14323 37077 14335 37080
rect 14277 37071 14335 37077
rect 15010 37068 15016 37080
rect 15068 37068 15074 37120
rect 17954 37068 17960 37120
rect 18012 37108 18018 37120
rect 18141 37111 18199 37117
rect 18141 37108 18153 37111
rect 18012 37080 18153 37108
rect 18012 37068 18018 37080
rect 18141 37077 18153 37080
rect 18187 37077 18199 37111
rect 18141 37071 18199 37077
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20073 37111 20131 37117
rect 20073 37108 20085 37111
rect 20036 37080 20085 37108
rect 20036 37068 20042 37080
rect 20073 37077 20085 37080
rect 20119 37077 20131 37111
rect 20073 37071 20131 37077
rect 24486 37068 24492 37120
rect 24544 37108 24550 37120
rect 24765 37111 24823 37117
rect 24765 37108 24777 37111
rect 24544 37080 24777 37108
rect 24544 37068 24550 37080
rect 24765 37077 24777 37080
rect 24811 37077 24823 37111
rect 24765 37071 24823 37077
rect 25130 37068 25136 37120
rect 25188 37108 25194 37120
rect 25501 37111 25559 37117
rect 25501 37108 25513 37111
rect 25188 37080 25513 37108
rect 25188 37068 25194 37080
rect 25501 37077 25513 37080
rect 25547 37077 25559 37111
rect 25501 37071 25559 37077
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 26476 37080 27353 37108
rect 26476 37068 26482 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27632 37108 27660 37148
rect 27706 37136 27712 37188
rect 27764 37176 27770 37188
rect 28828 37176 28856 37207
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 31202 37244 31208 37256
rect 31163 37216 31208 37244
rect 31202 37204 31208 37216
rect 31260 37204 31266 37256
rect 32309 37247 32367 37253
rect 32309 37213 32321 37247
rect 32355 37213 32367 37247
rect 33042 37244 33048 37256
rect 33003 37216 33048 37244
rect 32309 37207 32367 37213
rect 32324 37176 32352 37207
rect 33042 37204 33048 37216
rect 33100 37204 33106 37256
rect 33778 37244 33784 37256
rect 33739 37216 33784 37244
rect 33778 37204 33784 37216
rect 33836 37204 33842 37256
rect 35161 37247 35219 37253
rect 35161 37213 35173 37247
rect 35207 37244 35219 37247
rect 35207 37216 35894 37244
rect 35207 37213 35219 37216
rect 35161 37207 35219 37213
rect 27764 37148 28856 37176
rect 28920 37148 32352 37176
rect 35866 37176 35894 37216
rect 36078 37204 36084 37256
rect 36136 37244 36142 37256
rect 36173 37247 36231 37253
rect 36173 37244 36185 37247
rect 36136 37216 36185 37244
rect 36136 37204 36142 37216
rect 36173 37213 36185 37216
rect 36219 37213 36231 37247
rect 36173 37207 36231 37213
rect 36722 37204 36728 37256
rect 36780 37244 36786 37256
rect 37553 37247 37611 37253
rect 37553 37244 37565 37247
rect 36780 37216 37565 37244
rect 36780 37204 36786 37216
rect 37553 37213 37565 37216
rect 37599 37213 37611 37247
rect 37553 37207 37611 37213
rect 36538 37176 36544 37188
rect 35866 37148 36544 37176
rect 27764 37136 27770 37148
rect 28077 37111 28135 37117
rect 28077 37108 28089 37111
rect 27632 37080 28089 37108
rect 27341 37071 27399 37077
rect 28077 37077 28089 37080
rect 28123 37077 28135 37111
rect 28626 37108 28632 37120
rect 28587 37080 28632 37108
rect 28077 37071 28135 37077
rect 28626 37068 28632 37080
rect 28684 37068 28690 37120
rect 28718 37068 28724 37120
rect 28776 37108 28782 37120
rect 28920 37108 28948 37148
rect 36538 37136 36544 37148
rect 36596 37136 36602 37188
rect 28776 37080 28948 37108
rect 28776 37068 28782 37080
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 29917 37111 29975 37117
rect 29917 37108 29929 37111
rect 29696 37080 29929 37108
rect 29696 37068 29702 37080
rect 29917 37077 29929 37080
rect 29963 37077 29975 37111
rect 29917 37071 29975 37077
rect 31754 37068 31760 37120
rect 31812 37108 31818 37120
rect 32493 37111 32551 37117
rect 32493 37108 32505 37111
rect 31812 37080 32505 37108
rect 31812 37068 31818 37080
rect 32493 37077 32505 37080
rect 32539 37077 32551 37111
rect 32493 37071 32551 37077
rect 33502 37068 33508 37120
rect 33560 37108 33566 37120
rect 33965 37111 34023 37117
rect 33965 37108 33977 37111
rect 33560 37080 33977 37108
rect 33560 37068 33566 37080
rect 33965 37077 33977 37080
rect 34011 37077 34023 37111
rect 33965 37071 34023 37077
rect 35894 37068 35900 37120
rect 35952 37108 35958 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 35952 37080 36369 37108
rect 35952 37068 35958 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 37642 37108 37648 37120
rect 37603 37080 37648 37108
rect 36357 37071 36415 37077
rect 37642 37068 37648 37080
rect 37700 37068 37706 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1302 36864 1308 36916
rect 1360 36904 1366 36916
rect 1765 36907 1823 36913
rect 1765 36904 1777 36907
rect 1360 36876 1777 36904
rect 1360 36864 1366 36876
rect 1765 36873 1777 36876
rect 1811 36873 1823 36907
rect 1765 36867 1823 36873
rect 3237 36907 3295 36913
rect 3237 36873 3249 36907
rect 3283 36904 3295 36907
rect 8754 36904 8760 36916
rect 3283 36876 8760 36904
rect 3283 36873 3295 36876
rect 3237 36867 3295 36873
rect 8754 36864 8760 36876
rect 8812 36864 8818 36916
rect 11054 36864 11060 36916
rect 11112 36904 11118 36916
rect 11885 36907 11943 36913
rect 11885 36904 11897 36907
rect 11112 36876 11897 36904
rect 11112 36864 11118 36876
rect 11885 36873 11897 36876
rect 11931 36873 11943 36907
rect 11885 36867 11943 36873
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 15252 36876 19288 36904
rect 15252 36864 15258 36876
rect 3142 36836 3148 36848
rect 3103 36808 3148 36836
rect 3142 36796 3148 36808
rect 3200 36796 3206 36848
rect 3878 36796 3884 36848
rect 3936 36836 3942 36848
rect 4065 36839 4123 36845
rect 4065 36836 4077 36839
rect 3936 36808 4077 36836
rect 3936 36796 3942 36808
rect 4065 36805 4077 36808
rect 4111 36805 4123 36839
rect 4065 36799 4123 36805
rect 15470 36796 15476 36848
rect 15528 36836 15534 36848
rect 15657 36839 15715 36845
rect 15657 36836 15669 36839
rect 15528 36808 15669 36836
rect 15528 36796 15534 36808
rect 15657 36805 15669 36808
rect 15703 36805 15715 36839
rect 15657 36799 15715 36805
rect 17402 36796 17408 36848
rect 17460 36836 17466 36848
rect 19260 36836 19288 36876
rect 19334 36864 19340 36916
rect 19392 36904 19398 36916
rect 19613 36907 19671 36913
rect 19613 36904 19625 36907
rect 19392 36876 19625 36904
rect 19392 36864 19398 36876
rect 19613 36873 19625 36876
rect 19659 36873 19671 36907
rect 19613 36867 19671 36873
rect 22094 36864 22100 36916
rect 22152 36904 22158 36916
rect 22189 36907 22247 36913
rect 22189 36904 22201 36907
rect 22152 36876 22201 36904
rect 22152 36864 22158 36876
rect 22189 36873 22201 36876
rect 22235 36873 22247 36907
rect 23474 36904 23480 36916
rect 23435 36876 23480 36904
rect 22189 36867 22247 36873
rect 23474 36864 23480 36876
rect 23532 36864 23538 36916
rect 24762 36864 24768 36916
rect 24820 36904 24826 36916
rect 28626 36904 28632 36916
rect 24820 36876 28632 36904
rect 24820 36864 24826 36876
rect 28626 36864 28632 36876
rect 28684 36864 28690 36916
rect 36814 36904 36820 36916
rect 36775 36876 36820 36904
rect 36814 36864 36820 36876
rect 36872 36864 36878 36916
rect 17460 36808 18552 36836
rect 19260 36808 19564 36836
rect 17460 36796 17466 36808
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 2314 36768 2320 36780
rect 1627 36740 2320 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 2314 36728 2320 36740
rect 2372 36728 2378 36780
rect 2409 36771 2467 36777
rect 2409 36737 2421 36771
rect 2455 36768 2467 36771
rect 3050 36768 3056 36780
rect 2455 36740 3056 36768
rect 2455 36737 2467 36740
rect 2409 36731 2467 36737
rect 3050 36728 3056 36740
rect 3108 36728 3114 36780
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36737 5503 36771
rect 5445 36731 5503 36737
rect 5460 36700 5488 36731
rect 6454 36728 6460 36780
rect 6512 36768 6518 36780
rect 6733 36771 6791 36777
rect 6733 36768 6745 36771
rect 6512 36740 6745 36768
rect 6512 36728 6518 36740
rect 6733 36737 6745 36740
rect 6779 36737 6791 36771
rect 6733 36731 6791 36737
rect 9030 36728 9036 36780
rect 9088 36768 9094 36780
rect 9125 36771 9183 36777
rect 9125 36768 9137 36771
rect 9088 36740 9137 36768
rect 9088 36728 9094 36740
rect 9125 36737 9137 36740
rect 9171 36737 9183 36771
rect 11698 36768 11704 36780
rect 11659 36740 11704 36768
rect 9125 36731 9183 36737
rect 11698 36728 11704 36740
rect 11756 36728 11762 36780
rect 18524 36777 18552 36808
rect 17865 36771 17923 36777
rect 17865 36768 17877 36771
rect 16546 36740 17877 36768
rect 9214 36700 9220 36712
rect 5460 36672 9220 36700
rect 9214 36660 9220 36672
rect 9272 36660 9278 36712
rect 9398 36700 9404 36712
rect 9359 36672 9404 36700
rect 9398 36660 9404 36672
rect 9456 36660 9462 36712
rect 10962 36660 10968 36712
rect 11020 36700 11026 36712
rect 16546 36700 16574 36740
rect 17865 36737 17877 36740
rect 17911 36737 17923 36771
rect 17865 36731 17923 36737
rect 18509 36771 18567 36777
rect 18509 36737 18521 36771
rect 18555 36737 18567 36771
rect 19426 36768 19432 36780
rect 19387 36740 19432 36768
rect 18509 36731 18567 36737
rect 19426 36728 19432 36740
rect 19484 36728 19490 36780
rect 19536 36768 19564 36808
rect 20898 36796 20904 36848
rect 20956 36836 20962 36848
rect 20956 36808 30972 36836
rect 20956 36796 20962 36808
rect 21266 36768 21272 36780
rect 19536 36740 21272 36768
rect 21266 36728 21272 36740
rect 21324 36728 21330 36780
rect 22005 36771 22063 36777
rect 22005 36737 22017 36771
rect 22051 36768 22063 36771
rect 22370 36768 22376 36780
rect 22051 36740 22376 36768
rect 22051 36737 22063 36740
rect 22005 36731 22063 36737
rect 22370 36728 22376 36740
rect 22428 36728 22434 36780
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 23382 36768 23388 36780
rect 23339 36740 23388 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 23382 36728 23388 36740
rect 23440 36728 23446 36780
rect 25777 36771 25835 36777
rect 25777 36768 25789 36771
rect 23492 36740 25789 36768
rect 11020 36672 16574 36700
rect 11020 36660 11026 36672
rect 4249 36635 4307 36641
rect 4249 36601 4261 36635
rect 4295 36632 4307 36635
rect 5350 36632 5356 36644
rect 4295 36604 5356 36632
rect 4295 36601 4307 36604
rect 4249 36595 4307 36601
rect 5350 36592 5356 36604
rect 5408 36592 5414 36644
rect 10318 36592 10324 36644
rect 10376 36632 10382 36644
rect 15838 36632 15844 36644
rect 10376 36604 15844 36632
rect 10376 36592 10382 36604
rect 15838 36592 15844 36604
rect 15896 36592 15902 36644
rect 17681 36635 17739 36641
rect 17681 36601 17693 36635
rect 17727 36632 17739 36635
rect 17727 36604 21220 36632
rect 17727 36601 17739 36604
rect 17681 36595 17739 36601
rect 2501 36567 2559 36573
rect 2501 36533 2513 36567
rect 2547 36564 2559 36567
rect 3142 36564 3148 36576
rect 2547 36536 3148 36564
rect 2547 36533 2559 36536
rect 2501 36527 2559 36533
rect 3142 36524 3148 36536
rect 3200 36524 3206 36576
rect 5445 36567 5503 36573
rect 5445 36533 5457 36567
rect 5491 36564 5503 36567
rect 5534 36564 5540 36576
rect 5491 36536 5540 36564
rect 5491 36533 5503 36536
rect 5445 36527 5503 36533
rect 5534 36524 5540 36536
rect 5592 36524 5598 36576
rect 6549 36567 6607 36573
rect 6549 36533 6561 36567
rect 6595 36564 6607 36567
rect 10686 36564 10692 36576
rect 6595 36536 10692 36564
rect 6595 36533 6607 36536
rect 6549 36527 6607 36533
rect 10686 36524 10692 36536
rect 10744 36524 10750 36576
rect 18325 36567 18383 36573
rect 18325 36533 18337 36567
rect 18371 36564 18383 36567
rect 18690 36564 18696 36576
rect 18371 36536 18696 36564
rect 18371 36533 18383 36536
rect 18325 36527 18383 36533
rect 18690 36524 18696 36536
rect 18748 36524 18754 36576
rect 21192 36564 21220 36604
rect 21266 36592 21272 36644
rect 21324 36632 21330 36644
rect 23492 36632 23520 36740
rect 25777 36737 25789 36740
rect 25823 36737 25835 36771
rect 25777 36731 25835 36737
rect 26970 36728 26976 36780
rect 27028 36768 27034 36780
rect 28077 36771 28135 36777
rect 28077 36768 28089 36771
rect 27028 36740 28089 36768
rect 27028 36728 27034 36740
rect 28077 36737 28089 36740
rect 28123 36737 28135 36771
rect 28077 36731 28135 36737
rect 28994 36728 29000 36780
rect 29052 36768 29058 36780
rect 30944 36777 30972 36808
rect 38010 36796 38016 36848
rect 38068 36836 38074 36848
rect 38105 36839 38163 36845
rect 38105 36836 38117 36839
rect 38068 36808 38117 36836
rect 38068 36796 38074 36808
rect 38105 36805 38117 36808
rect 38151 36805 38163 36839
rect 38105 36799 38163 36805
rect 29273 36771 29331 36777
rect 29273 36768 29285 36771
rect 29052 36740 29285 36768
rect 29052 36728 29058 36740
rect 29273 36737 29285 36740
rect 29319 36737 29331 36771
rect 29273 36731 29331 36737
rect 30929 36771 30987 36777
rect 30929 36737 30941 36771
rect 30975 36737 30987 36771
rect 30929 36731 30987 36737
rect 35894 36728 35900 36780
rect 35952 36768 35958 36780
rect 36633 36771 36691 36777
rect 35952 36740 35997 36768
rect 35952 36728 35958 36740
rect 36633 36737 36645 36771
rect 36679 36737 36691 36771
rect 36633 36731 36691 36737
rect 28718 36700 28724 36712
rect 21324 36604 23520 36632
rect 23584 36672 28724 36700
rect 21324 36592 21330 36604
rect 23584 36564 23612 36672
rect 28718 36660 28724 36672
rect 28776 36660 28782 36712
rect 33042 36700 33048 36712
rect 30484 36672 33048 36700
rect 25593 36635 25651 36641
rect 25593 36601 25605 36635
rect 25639 36632 25651 36635
rect 27893 36635 27951 36641
rect 25639 36604 26234 36632
rect 25639 36601 25651 36604
rect 25593 36595 25651 36601
rect 21192 36536 23612 36564
rect 26206 36564 26234 36604
rect 27893 36601 27905 36635
rect 27939 36632 27951 36635
rect 30484 36632 30512 36672
rect 33042 36660 33048 36672
rect 33100 36660 33106 36712
rect 36648 36700 36676 36731
rect 35866 36672 36676 36700
rect 27939 36604 30512 36632
rect 30745 36635 30803 36641
rect 27939 36601 27951 36604
rect 27893 36595 27951 36601
rect 30745 36601 30757 36635
rect 30791 36632 30803 36635
rect 35866 36632 35894 36672
rect 30791 36604 35894 36632
rect 36081 36635 36139 36641
rect 30791 36601 30803 36604
rect 30745 36595 30803 36601
rect 36081 36601 36093 36635
rect 36127 36632 36139 36635
rect 38654 36632 38660 36644
rect 36127 36604 38660 36632
rect 36127 36601 36139 36604
rect 36081 36595 36139 36601
rect 38654 36592 38660 36604
rect 38712 36592 38718 36644
rect 28442 36564 28448 36576
rect 26206 36536 28448 36564
rect 28442 36524 28448 36536
rect 28500 36524 28506 36576
rect 28534 36524 28540 36576
rect 28592 36564 28598 36576
rect 29089 36567 29147 36573
rect 29089 36564 29101 36567
rect 28592 36536 29101 36564
rect 28592 36524 28598 36536
rect 29089 36533 29101 36536
rect 29135 36533 29147 36567
rect 29089 36527 29147 36533
rect 37826 36524 37832 36576
rect 37884 36564 37890 36576
rect 38197 36567 38255 36573
rect 38197 36564 38209 36567
rect 37884 36536 38209 36564
rect 37884 36524 37890 36536
rect 38197 36533 38209 36536
rect 38243 36533 38255 36567
rect 38197 36527 38255 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1762 36360 1768 36372
rect 1723 36332 1768 36360
rect 1762 36320 1768 36332
rect 1820 36320 1826 36372
rect 2314 36320 2320 36372
rect 2372 36360 2378 36372
rect 5353 36363 5411 36369
rect 5353 36360 5365 36363
rect 2372 36332 5365 36360
rect 2372 36320 2378 36332
rect 5353 36329 5365 36332
rect 5399 36329 5411 36363
rect 5353 36323 5411 36329
rect 5718 36320 5724 36372
rect 5776 36360 5782 36372
rect 9125 36363 9183 36369
rect 9125 36360 9137 36363
rect 5776 36332 9137 36360
rect 5776 36320 5782 36332
rect 9125 36329 9137 36332
rect 9171 36329 9183 36363
rect 9125 36323 9183 36329
rect 15838 36320 15844 36372
rect 15896 36360 15902 36372
rect 21910 36360 21916 36372
rect 15896 36332 21916 36360
rect 15896 36320 15902 36332
rect 21910 36320 21916 36332
rect 21968 36320 21974 36372
rect 22370 36360 22376 36372
rect 22331 36332 22376 36360
rect 22370 36320 22376 36332
rect 22428 36320 22434 36372
rect 24486 36320 24492 36372
rect 24544 36360 24550 36372
rect 31202 36360 31208 36372
rect 24544 36332 31208 36360
rect 24544 36320 24550 36332
rect 31202 36320 31208 36332
rect 31260 36320 31266 36372
rect 37458 36360 37464 36372
rect 37419 36332 37464 36360
rect 37458 36320 37464 36332
rect 37516 36320 37522 36372
rect 14 36184 20 36236
rect 72 36224 78 36236
rect 72 36196 2544 36224
rect 72 36184 78 36196
rect 2516 36165 2544 36196
rect 3142 36184 3148 36236
rect 3200 36224 3206 36236
rect 10962 36224 10968 36236
rect 3200 36196 10968 36224
rect 3200 36184 3206 36196
rect 10962 36184 10968 36196
rect 11020 36184 11026 36236
rect 28718 36184 28724 36236
rect 28776 36224 28782 36236
rect 28776 36196 38056 36224
rect 28776 36184 28782 36196
rect 1581 36159 1639 36165
rect 1581 36125 1593 36159
rect 1627 36125 1639 36159
rect 1581 36119 1639 36125
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36125 2559 36159
rect 5534 36156 5540 36168
rect 5495 36128 5540 36156
rect 2501 36119 2559 36125
rect 1596 36088 1624 36119
rect 5534 36116 5540 36128
rect 5592 36116 5598 36168
rect 9309 36159 9367 36165
rect 9309 36125 9321 36159
rect 9355 36156 9367 36159
rect 12250 36156 12256 36168
rect 9355 36128 12256 36156
rect 9355 36125 9367 36128
rect 9309 36119 9367 36125
rect 12250 36116 12256 36128
rect 12308 36116 12314 36168
rect 22557 36159 22615 36165
rect 22557 36125 22569 36159
rect 22603 36156 22615 36159
rect 24486 36156 24492 36168
rect 22603 36128 24492 36156
rect 22603 36125 22615 36128
rect 22557 36119 22615 36125
rect 24486 36116 24492 36128
rect 24544 36116 24550 36168
rect 33778 36156 33784 36168
rect 26206 36128 33784 36156
rect 2866 36088 2872 36100
rect 1596 36060 2872 36088
rect 2866 36048 2872 36060
rect 2924 36048 2930 36100
rect 21542 36048 21548 36100
rect 21600 36088 21606 36100
rect 26206 36088 26234 36128
rect 33778 36116 33784 36128
rect 33836 36116 33842 36168
rect 36170 36116 36176 36168
rect 36228 36156 36234 36168
rect 38028 36165 38056 36196
rect 36357 36159 36415 36165
rect 36357 36156 36369 36159
rect 36228 36128 36369 36156
rect 36228 36116 36234 36128
rect 36357 36125 36369 36128
rect 36403 36125 36415 36159
rect 36357 36119 36415 36125
rect 37277 36159 37335 36165
rect 37277 36125 37289 36159
rect 37323 36125 37335 36159
rect 37277 36119 37335 36125
rect 38013 36159 38071 36165
rect 38013 36125 38025 36159
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 21600 36060 26234 36088
rect 21600 36048 21606 36060
rect 29914 36048 29920 36100
rect 29972 36088 29978 36100
rect 37292 36088 37320 36119
rect 29972 36060 37320 36088
rect 29972 36048 29978 36060
rect 2317 36023 2375 36029
rect 2317 35989 2329 36023
rect 2363 36020 2375 36023
rect 4062 36020 4068 36032
rect 2363 35992 4068 36020
rect 2363 35989 2375 35992
rect 2317 35983 2375 35989
rect 4062 35980 4068 35992
rect 4120 35980 4126 36032
rect 36170 36020 36176 36032
rect 36131 35992 36176 36020
rect 36170 35980 36176 35992
rect 36228 35980 36234 36032
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 11701 35819 11759 35825
rect 11701 35785 11713 35819
rect 11747 35816 11759 35819
rect 12986 35816 12992 35828
rect 11747 35788 12992 35816
rect 11747 35785 11759 35788
rect 11701 35779 11759 35785
rect 12986 35776 12992 35788
rect 13044 35776 13050 35828
rect 39298 35748 39304 35760
rect 36924 35720 39304 35748
rect 11882 35680 11888 35692
rect 11843 35652 11888 35680
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 36924 35689 36952 35720
rect 39298 35708 39304 35720
rect 39356 35708 39362 35760
rect 36909 35683 36967 35689
rect 36909 35649 36921 35683
rect 36955 35649 36967 35683
rect 36909 35643 36967 35649
rect 38013 35683 38071 35689
rect 38013 35649 38025 35683
rect 38059 35649 38071 35683
rect 38013 35643 38071 35649
rect 1578 35612 1584 35624
rect 1539 35584 1584 35612
rect 1578 35572 1584 35584
rect 1636 35572 1642 35624
rect 1857 35615 1915 35621
rect 1857 35581 1869 35615
rect 1903 35612 1915 35615
rect 2130 35612 2136 35624
rect 1903 35584 2136 35612
rect 1903 35581 1915 35584
rect 1857 35575 1915 35581
rect 2130 35572 2136 35584
rect 2188 35572 2194 35624
rect 35526 35572 35532 35624
rect 35584 35612 35590 35624
rect 38028 35612 38056 35643
rect 35584 35584 38056 35612
rect 35584 35572 35590 35584
rect 34514 35436 34520 35488
rect 34572 35476 34578 35488
rect 36725 35479 36783 35485
rect 36725 35476 36737 35479
rect 34572 35448 36737 35476
rect 34572 35436 34578 35448
rect 36725 35445 36737 35448
rect 36771 35445 36783 35479
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 36725 35439 36783 35445
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 38197 35275 38255 35281
rect 38197 35241 38209 35275
rect 38243 35272 38255 35275
rect 38286 35272 38292 35284
rect 38243 35244 38292 35272
rect 38243 35241 38255 35244
rect 38197 35235 38255 35241
rect 38286 35232 38292 35244
rect 38344 35232 38350 35284
rect 11698 35164 11704 35216
rect 11756 35204 11762 35216
rect 28074 35204 28080 35216
rect 11756 35176 28080 35204
rect 11756 35164 11762 35176
rect 28074 35164 28080 35176
rect 28132 35164 28138 35216
rect 10686 35068 10692 35080
rect 10647 35040 10692 35068
rect 10686 35028 10692 35040
rect 10744 35028 10750 35080
rect 37274 35028 37280 35080
rect 37332 35068 37338 35080
rect 38013 35071 38071 35077
rect 38013 35068 38025 35071
rect 37332 35040 38025 35068
rect 37332 35028 37338 35040
rect 38013 35037 38025 35040
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 10781 34935 10839 34941
rect 10781 34901 10793 34935
rect 10827 34932 10839 34935
rect 13354 34932 13360 34944
rect 10827 34904 13360 34932
rect 10827 34901 10839 34904
rect 10781 34895 10839 34901
rect 13354 34892 13360 34904
rect 13412 34892 13418 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 5810 34728 5816 34740
rect 1627 34700 5816 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 5810 34688 5816 34700
rect 5868 34688 5874 34740
rect 27617 34731 27675 34737
rect 27617 34697 27629 34731
rect 27663 34728 27675 34731
rect 29730 34728 29736 34740
rect 27663 34700 29736 34728
rect 27663 34697 27675 34700
rect 27617 34691 27675 34697
rect 29730 34688 29736 34700
rect 29788 34688 29794 34740
rect 35437 34731 35495 34737
rect 35437 34697 35449 34731
rect 35483 34728 35495 34731
rect 35894 34728 35900 34740
rect 35483 34700 35900 34728
rect 35483 34697 35495 34700
rect 35437 34691 35495 34697
rect 35894 34688 35900 34700
rect 35952 34688 35958 34740
rect 11146 34660 11152 34672
rect 6886 34632 11152 34660
rect 1762 34592 1768 34604
rect 1723 34564 1768 34592
rect 1762 34552 1768 34564
rect 1820 34552 1826 34604
rect 4062 34552 4068 34604
rect 4120 34592 4126 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 4120 34564 6561 34592
rect 4120 34552 4126 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6549 34555 6607 34561
rect 6641 34527 6699 34533
rect 6641 34493 6653 34527
rect 6687 34524 6699 34527
rect 6886 34524 6914 34632
rect 11146 34620 11152 34632
rect 11204 34620 11210 34672
rect 10778 34592 10784 34604
rect 10739 34564 10784 34592
rect 10778 34552 10784 34564
rect 10836 34552 10842 34604
rect 27798 34592 27804 34604
rect 27759 34564 27804 34592
rect 27798 34552 27804 34564
rect 27856 34552 27862 34604
rect 28994 34552 29000 34604
rect 29052 34592 29058 34604
rect 34701 34595 34759 34601
rect 34701 34592 34713 34595
rect 29052 34564 34713 34592
rect 29052 34552 29058 34564
rect 34701 34561 34713 34564
rect 34747 34561 34759 34595
rect 34701 34555 34759 34561
rect 34977 34595 35035 34601
rect 34977 34561 34989 34595
rect 35023 34592 35035 34595
rect 35621 34595 35679 34601
rect 35621 34592 35633 34595
rect 35023 34564 35633 34592
rect 35023 34561 35035 34564
rect 34977 34555 35035 34561
rect 35621 34561 35633 34564
rect 35667 34561 35679 34595
rect 35621 34555 35679 34561
rect 6687 34496 6914 34524
rect 6687 34493 6699 34496
rect 6641 34487 6699 34493
rect 37182 34484 37188 34536
rect 37240 34524 37246 34536
rect 37461 34527 37519 34533
rect 37461 34524 37473 34527
rect 37240 34496 37473 34524
rect 37240 34484 37246 34496
rect 37461 34493 37473 34496
rect 37507 34493 37519 34527
rect 37734 34524 37740 34536
rect 37695 34496 37740 34524
rect 37461 34487 37519 34493
rect 37734 34484 37740 34496
rect 37792 34484 37798 34536
rect 10502 34348 10508 34400
rect 10560 34388 10566 34400
rect 10873 34391 10931 34397
rect 10873 34388 10885 34391
rect 10560 34360 10885 34388
rect 10560 34348 10566 34360
rect 10873 34357 10885 34360
rect 10919 34357 10931 34391
rect 10873 34351 10931 34357
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 10873 34187 10931 34193
rect 10873 34153 10885 34187
rect 10919 34184 10931 34187
rect 11882 34184 11888 34196
rect 10919 34156 11888 34184
rect 10919 34153 10931 34156
rect 10873 34147 10931 34153
rect 11882 34144 11888 34156
rect 11940 34144 11946 34196
rect 27522 34184 27528 34196
rect 27483 34156 27528 34184
rect 27522 34144 27528 34156
rect 27580 34144 27586 34196
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33980 10839 33983
rect 12526 33980 12532 33992
rect 10827 33952 12532 33980
rect 10827 33949 10839 33952
rect 10781 33943 10839 33949
rect 12526 33940 12532 33952
rect 12584 33940 12590 33992
rect 22094 33940 22100 33992
rect 22152 33980 22158 33992
rect 22649 33983 22707 33989
rect 22649 33980 22661 33983
rect 22152 33952 22661 33980
rect 22152 33940 22158 33952
rect 22649 33949 22661 33952
rect 22695 33949 22707 33983
rect 22649 33943 22707 33949
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33980 24639 33983
rect 24762 33980 24768 33992
rect 24627 33952 24768 33980
rect 24627 33949 24639 33952
rect 24581 33943 24639 33949
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 26878 33940 26884 33992
rect 26936 33980 26942 33992
rect 27709 33983 27767 33989
rect 27709 33980 27721 33983
rect 26936 33952 27721 33980
rect 26936 33940 26942 33952
rect 27709 33949 27721 33952
rect 27755 33949 27767 33983
rect 27709 33943 27767 33949
rect 23566 33872 23572 33924
rect 23624 33912 23630 33924
rect 24673 33915 24731 33921
rect 24673 33912 24685 33915
rect 23624 33884 24685 33912
rect 23624 33872 23630 33884
rect 24673 33881 24685 33884
rect 24719 33881 24731 33915
rect 24673 33875 24731 33881
rect 22741 33847 22799 33853
rect 22741 33813 22753 33847
rect 22787 33844 22799 33847
rect 23658 33844 23664 33856
rect 22787 33816 23664 33844
rect 22787 33813 22799 33816
rect 22741 33807 22799 33813
rect 23658 33804 23664 33816
rect 23716 33804 23722 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 23477 33643 23535 33649
rect 23477 33609 23489 33643
rect 23523 33640 23535 33643
rect 24578 33640 24584 33652
rect 23523 33612 24584 33640
rect 23523 33609 23535 33612
rect 23477 33603 23535 33609
rect 24578 33600 24584 33612
rect 24636 33600 24642 33652
rect 106 33464 112 33516
rect 164 33504 170 33516
rect 1765 33507 1823 33513
rect 1765 33504 1777 33507
rect 164 33476 1777 33504
rect 164 33464 170 33476
rect 1765 33473 1777 33476
rect 1811 33473 1823 33507
rect 1765 33467 1823 33473
rect 2409 33507 2467 33513
rect 2409 33473 2421 33507
rect 2455 33473 2467 33507
rect 23658 33504 23664 33516
rect 23619 33476 23664 33504
rect 2409 33467 2467 33473
rect 14 33396 20 33448
rect 72 33436 78 33448
rect 2424 33436 2452 33467
rect 23658 33464 23664 33476
rect 23716 33464 23722 33516
rect 30377 33507 30435 33513
rect 30377 33473 30389 33507
rect 30423 33504 30435 33507
rect 34514 33504 34520 33516
rect 30423 33476 34520 33504
rect 30423 33473 30435 33476
rect 30377 33467 30435 33473
rect 34514 33464 34520 33476
rect 34572 33464 34578 33516
rect 38102 33504 38108 33516
rect 38063 33476 38108 33504
rect 38102 33464 38108 33476
rect 38160 33464 38166 33516
rect 72 33408 2452 33436
rect 72 33396 78 33408
rect 1581 33371 1639 33377
rect 1581 33337 1593 33371
rect 1627 33368 1639 33371
rect 3418 33368 3424 33380
rect 1627 33340 3424 33368
rect 1627 33337 1639 33340
rect 1581 33331 1639 33337
rect 3418 33328 3424 33340
rect 3476 33328 3482 33380
rect 20438 33328 20444 33380
rect 20496 33368 20502 33380
rect 30469 33371 30527 33377
rect 30469 33368 30481 33371
rect 20496 33340 30481 33368
rect 20496 33328 20502 33340
rect 30469 33337 30481 33340
rect 30515 33337 30527 33371
rect 38289 33371 38347 33377
rect 38289 33368 38301 33371
rect 30469 33331 30527 33337
rect 35866 33340 38301 33368
rect 2225 33303 2283 33309
rect 2225 33269 2237 33303
rect 2271 33300 2283 33303
rect 3970 33300 3976 33312
rect 2271 33272 3976 33300
rect 2271 33269 2283 33272
rect 2225 33263 2283 33269
rect 3970 33260 3976 33272
rect 4028 33260 4034 33312
rect 21174 33260 21180 33312
rect 21232 33300 21238 33312
rect 35866 33300 35894 33340
rect 38289 33337 38301 33340
rect 38335 33337 38347 33371
rect 38289 33331 38347 33337
rect 21232 33272 35894 33300
rect 21232 33260 21238 33272
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 2961 33099 3019 33105
rect 2961 33096 2973 33099
rect 2924 33068 2973 33096
rect 2924 33056 2930 33068
rect 2961 33065 2973 33068
rect 3007 33065 3019 33099
rect 2961 33059 3019 33065
rect 1118 32988 1124 33040
rect 1176 33028 1182 33040
rect 2317 33031 2375 33037
rect 2317 33028 2329 33031
rect 1176 33000 2329 33028
rect 1176 32988 1182 33000
rect 2317 32997 2329 33000
rect 2363 32997 2375 33031
rect 2317 32991 2375 32997
rect 1486 32920 1492 32972
rect 1544 32960 1550 32972
rect 1544 32932 2544 32960
rect 1544 32920 1550 32932
rect 2516 32901 2544 32932
rect 1581 32895 1639 32901
rect 1581 32861 1593 32895
rect 1627 32892 1639 32895
rect 2501 32895 2559 32901
rect 1627 32864 2268 32892
rect 1627 32861 1639 32864
rect 1581 32855 1639 32861
rect 2240 32768 2268 32864
rect 2501 32861 2513 32895
rect 2547 32861 2559 32895
rect 2501 32855 2559 32861
rect 2682 32852 2688 32904
rect 2740 32892 2746 32904
rect 3145 32895 3203 32901
rect 3145 32892 3157 32895
rect 2740 32864 3157 32892
rect 2740 32852 2746 32864
rect 3145 32861 3157 32864
rect 3191 32861 3203 32895
rect 3145 32855 3203 32861
rect 6822 32852 6828 32904
rect 6880 32892 6886 32904
rect 6917 32895 6975 32901
rect 6917 32892 6929 32895
rect 6880 32864 6929 32892
rect 6880 32852 6886 32864
rect 6917 32861 6929 32864
rect 6963 32861 6975 32895
rect 6917 32855 6975 32861
rect 29733 32895 29791 32901
rect 29733 32861 29745 32895
rect 29779 32892 29791 32895
rect 36170 32892 36176 32904
rect 29779 32864 36176 32892
rect 29779 32861 29791 32864
rect 29733 32855 29791 32861
rect 36170 32852 36176 32864
rect 36228 32852 36234 32904
rect 1762 32756 1768 32768
rect 1723 32728 1768 32756
rect 1762 32716 1768 32728
rect 1820 32716 1826 32768
rect 2222 32756 2228 32768
rect 2183 32728 2228 32756
rect 2222 32716 2228 32728
rect 2280 32716 2286 32768
rect 7009 32759 7067 32765
rect 7009 32725 7021 32759
rect 7055 32756 7067 32759
rect 7190 32756 7196 32768
rect 7055 32728 7196 32756
rect 7055 32725 7067 32728
rect 7009 32719 7067 32725
rect 7190 32716 7196 32728
rect 7248 32716 7254 32768
rect 25314 32716 25320 32768
rect 25372 32756 25378 32768
rect 29825 32759 29883 32765
rect 29825 32756 29837 32759
rect 25372 32728 29837 32756
rect 25372 32716 25378 32728
rect 29825 32725 29837 32728
rect 29871 32725 29883 32759
rect 29825 32719 29883 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 2222 32512 2228 32564
rect 2280 32552 2286 32564
rect 22554 32552 22560 32564
rect 2280 32524 22560 32552
rect 2280 32512 2286 32524
rect 22554 32512 22560 32524
rect 22612 32512 22618 32564
rect 5350 32444 5356 32496
rect 5408 32484 5414 32496
rect 27154 32484 27160 32496
rect 5408 32456 27160 32484
rect 5408 32444 5414 32456
rect 27154 32444 27160 32456
rect 27212 32444 27218 32496
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32385 1639 32419
rect 3050 32416 3056 32428
rect 3011 32388 3056 32416
rect 1581 32379 1639 32385
rect 1596 32348 1624 32379
rect 3050 32376 3056 32388
rect 3108 32376 3114 32428
rect 3694 32416 3700 32428
rect 3655 32388 3700 32416
rect 3694 32376 3700 32388
rect 3752 32376 3758 32428
rect 28534 32416 28540 32428
rect 28495 32388 28540 32416
rect 28534 32376 28540 32388
rect 28592 32376 28598 32428
rect 33778 32376 33784 32428
rect 33836 32416 33842 32428
rect 37737 32419 37795 32425
rect 37737 32416 37749 32419
rect 33836 32388 37749 32416
rect 33836 32376 33842 32388
rect 37737 32385 37749 32388
rect 37783 32385 37795 32419
rect 37737 32379 37795 32385
rect 4982 32348 4988 32360
rect 1596 32320 4988 32348
rect 4982 32308 4988 32320
rect 5040 32308 5046 32360
rect 37458 32348 37464 32360
rect 37419 32320 37464 32348
rect 37458 32308 37464 32320
rect 37516 32308 37522 32360
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 1946 32172 1952 32224
rect 2004 32212 2010 32224
rect 2682 32212 2688 32224
rect 2004 32184 2688 32212
rect 2004 32172 2010 32184
rect 2682 32172 2688 32184
rect 2740 32212 2746 32224
rect 2869 32215 2927 32221
rect 2869 32212 2881 32215
rect 2740 32184 2881 32212
rect 2740 32172 2746 32184
rect 2869 32181 2881 32184
rect 2915 32181 2927 32215
rect 2869 32175 2927 32181
rect 3513 32215 3571 32221
rect 3513 32181 3525 32215
rect 3559 32212 3571 32215
rect 6638 32212 6644 32224
rect 3559 32184 6644 32212
rect 3559 32181 3571 32184
rect 3513 32175 3571 32181
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 28534 32172 28540 32224
rect 28592 32212 28598 32224
rect 28629 32215 28687 32221
rect 28629 32212 28641 32215
rect 28592 32184 28641 32212
rect 28592 32172 28598 32184
rect 28629 32181 28641 32184
rect 28675 32181 28687 32215
rect 28629 32175 28687 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 2958 32008 2964 32020
rect 2919 31980 2964 32008
rect 2958 31968 2964 31980
rect 3016 31968 3022 32020
rect 35526 32008 35532 32020
rect 35487 31980 35532 32008
rect 35526 31968 35532 31980
rect 35584 31968 35590 32020
rect 1673 31943 1731 31949
rect 1673 31909 1685 31943
rect 1719 31940 1731 31943
rect 3786 31940 3792 31952
rect 1719 31912 3792 31940
rect 1719 31909 1731 31912
rect 1673 31903 1731 31909
rect 3786 31900 3792 31912
rect 3844 31900 3850 31952
rect 5626 31940 5632 31952
rect 3988 31912 5632 31940
rect 2409 31875 2467 31881
rect 2409 31872 2421 31875
rect 1872 31844 2421 31872
rect 842 31764 848 31816
rect 900 31804 906 31816
rect 1872 31813 1900 31844
rect 2409 31841 2421 31844
rect 2455 31841 2467 31875
rect 3988 31872 4016 31912
rect 5626 31900 5632 31912
rect 5684 31900 5690 31952
rect 2409 31835 2467 31841
rect 2516 31844 4016 31872
rect 4065 31875 4123 31881
rect 1857 31807 1915 31813
rect 900 31776 1808 31804
rect 900 31764 906 31776
rect 1780 31736 1808 31776
rect 1857 31773 1869 31807
rect 1903 31773 1915 31807
rect 1857 31767 1915 31773
rect 2317 31807 2375 31813
rect 2317 31773 2329 31807
rect 2363 31804 2375 31807
rect 2516 31804 2544 31844
rect 4065 31841 4077 31875
rect 4111 31872 4123 31875
rect 5442 31872 5448 31884
rect 4111 31844 5448 31872
rect 4111 31841 4123 31844
rect 4065 31835 4123 31841
rect 5442 31832 5448 31844
rect 5500 31832 5506 31884
rect 3145 31807 3203 31813
rect 3145 31804 3157 31807
rect 2363 31776 2544 31804
rect 2608 31776 3157 31804
rect 2363 31773 2375 31776
rect 2317 31767 2375 31773
rect 2608 31736 2636 31776
rect 3145 31773 3157 31776
rect 3191 31804 3203 31807
rect 3973 31807 4031 31813
rect 3191 31776 3924 31804
rect 3191 31773 3203 31776
rect 3145 31767 3203 31773
rect 1780 31708 2636 31736
rect 3896 31736 3924 31776
rect 3973 31773 3985 31807
rect 4019 31804 4031 31807
rect 17954 31804 17960 31816
rect 4019 31776 7328 31804
rect 17915 31776 17960 31804
rect 4019 31773 4031 31776
rect 3973 31767 4031 31773
rect 7300 31748 7328 31776
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18049 31807 18107 31813
rect 18049 31773 18061 31807
rect 18095 31804 18107 31807
rect 19334 31804 19340 31816
rect 18095 31776 19340 31804
rect 18095 31773 18107 31776
rect 18049 31767 18107 31773
rect 19334 31764 19340 31776
rect 19392 31764 19398 31816
rect 33870 31764 33876 31816
rect 33928 31804 33934 31816
rect 35713 31807 35771 31813
rect 35713 31804 35725 31807
rect 33928 31776 35725 31804
rect 33928 31764 33934 31776
rect 35713 31773 35725 31776
rect 35759 31773 35771 31807
rect 35713 31767 35771 31773
rect 37182 31764 37188 31816
rect 37240 31804 37246 31816
rect 37461 31807 37519 31813
rect 37461 31804 37473 31807
rect 37240 31776 37473 31804
rect 37240 31764 37246 31776
rect 37461 31773 37473 31776
rect 37507 31773 37519 31807
rect 37461 31767 37519 31773
rect 37550 31764 37556 31816
rect 37608 31804 37614 31816
rect 37737 31807 37795 31813
rect 37737 31804 37749 31807
rect 37608 31776 37749 31804
rect 37608 31764 37614 31776
rect 37737 31773 37749 31776
rect 37783 31773 37795 31807
rect 37737 31767 37795 31773
rect 5074 31736 5080 31748
rect 3896 31708 5080 31736
rect 5074 31696 5080 31708
rect 5132 31696 5138 31748
rect 7282 31696 7288 31748
rect 7340 31696 7346 31748
rect 11698 31628 11704 31680
rect 11756 31668 11762 31680
rect 11793 31671 11851 31677
rect 11793 31668 11805 31671
rect 11756 31640 11805 31668
rect 11756 31628 11762 31640
rect 11793 31637 11805 31640
rect 11839 31637 11851 31671
rect 11793 31631 11851 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 4982 31464 4988 31476
rect 4943 31436 4988 31464
rect 4982 31424 4988 31436
rect 5040 31424 5046 31476
rect 19426 31424 19432 31476
rect 19484 31464 19490 31476
rect 20441 31467 20499 31473
rect 20441 31464 20453 31467
rect 19484 31436 20453 31464
rect 19484 31424 19490 31436
rect 20441 31433 20453 31436
rect 20487 31433 20499 31467
rect 20441 31427 20499 31433
rect 750 31356 756 31408
rect 808 31396 814 31408
rect 4065 31399 4123 31405
rect 4065 31396 4077 31399
rect 808 31368 4077 31396
rect 808 31356 814 31368
rect 4065 31365 4077 31368
rect 4111 31365 4123 31399
rect 4065 31359 4123 31365
rect 1394 31288 1400 31340
rect 1452 31328 1458 31340
rect 1857 31331 1915 31337
rect 1857 31328 1869 31331
rect 1452 31300 1869 31328
rect 1452 31288 1458 31300
rect 1857 31297 1869 31300
rect 1903 31297 1915 31331
rect 1857 31291 1915 31297
rect 3237 31331 3295 31337
rect 3237 31297 3249 31331
rect 3283 31328 3295 31331
rect 3510 31328 3516 31340
rect 3283 31300 3516 31328
rect 3283 31297 3295 31300
rect 3237 31291 3295 31297
rect 3510 31288 3516 31300
rect 3568 31288 3574 31340
rect 3973 31331 4031 31337
rect 3973 31297 3985 31331
rect 4019 31297 4031 31331
rect 3973 31291 4031 31297
rect 5169 31331 5227 31337
rect 5169 31297 5181 31331
rect 5215 31328 5227 31331
rect 6546 31328 6552 31340
rect 5215 31300 6552 31328
rect 5215 31297 5227 31300
rect 5169 31291 5227 31297
rect 2501 31263 2559 31269
rect 2501 31229 2513 31263
rect 2547 31229 2559 31263
rect 3988 31260 4016 31291
rect 6546 31288 6552 31300
rect 6604 31288 6610 31340
rect 11701 31331 11759 31337
rect 11701 31297 11713 31331
rect 11747 31328 11759 31331
rect 12066 31328 12072 31340
rect 11747 31300 12072 31328
rect 11747 31297 11759 31300
rect 11701 31291 11759 31297
rect 12066 31288 12072 31300
rect 12124 31288 12130 31340
rect 18690 31328 18696 31340
rect 18651 31300 18696 31328
rect 18690 31288 18696 31300
rect 18748 31288 18754 31340
rect 19337 31331 19395 31337
rect 19337 31297 19349 31331
rect 19383 31297 19395 31331
rect 20622 31328 20628 31340
rect 20583 31300 20628 31328
rect 19337 31291 19395 31297
rect 9122 31260 9128 31272
rect 3988 31232 9128 31260
rect 2501 31223 2559 31229
rect 1854 31152 1860 31204
rect 1912 31192 1918 31204
rect 2516 31192 2544 31223
rect 9122 31220 9128 31232
rect 9180 31220 9186 31272
rect 12434 31220 12440 31272
rect 12492 31260 12498 31272
rect 12492 31232 12537 31260
rect 12492 31220 12498 31232
rect 17586 31220 17592 31272
rect 17644 31260 17650 31272
rect 19352 31260 19380 31291
rect 20622 31288 20628 31300
rect 20680 31288 20686 31340
rect 17644 31232 19380 31260
rect 17644 31220 17650 31232
rect 1912 31164 2544 31192
rect 18785 31195 18843 31201
rect 1912 31152 1918 31164
rect 18785 31161 18797 31195
rect 18831 31192 18843 31195
rect 20346 31192 20352 31204
rect 18831 31164 20352 31192
rect 18831 31161 18843 31164
rect 18785 31155 18843 31161
rect 20346 31152 20352 31164
rect 20404 31152 20410 31204
rect 1026 31084 1032 31136
rect 1084 31124 1090 31136
rect 1949 31127 2007 31133
rect 1949 31124 1961 31127
rect 1084 31096 1961 31124
rect 1084 31084 1090 31096
rect 1949 31093 1961 31096
rect 1995 31093 2007 31127
rect 1949 31087 2007 31093
rect 3329 31127 3387 31133
rect 3329 31093 3341 31127
rect 3375 31124 3387 31127
rect 4706 31124 4712 31136
rect 3375 31096 4712 31124
rect 3375 31093 3387 31096
rect 3329 31087 3387 31093
rect 4706 31084 4712 31096
rect 4764 31084 4770 31136
rect 10226 31084 10232 31136
rect 10284 31124 10290 31136
rect 11793 31127 11851 31133
rect 11793 31124 11805 31127
rect 10284 31096 11805 31124
rect 10284 31084 10290 31096
rect 11793 31093 11805 31096
rect 11839 31093 11851 31127
rect 11793 31087 11851 31093
rect 19429 31127 19487 31133
rect 19429 31093 19441 31127
rect 19475 31124 19487 31127
rect 19978 31124 19984 31136
rect 19475 31096 19984 31124
rect 19475 31093 19487 31096
rect 19429 31087 19487 31093
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 6546 30920 6552 30932
rect 6507 30892 6552 30920
rect 6546 30880 6552 30892
rect 6604 30880 6610 30932
rect 12250 30880 12256 30932
rect 12308 30920 12314 30932
rect 13357 30923 13415 30929
rect 13357 30920 13369 30923
rect 12308 30892 13369 30920
rect 12308 30880 12314 30892
rect 13357 30889 13369 30892
rect 13403 30889 13415 30923
rect 13357 30883 13415 30889
rect 7837 30855 7895 30861
rect 7837 30821 7849 30855
rect 7883 30852 7895 30855
rect 12710 30852 12716 30864
rect 7883 30824 12716 30852
rect 7883 30821 7895 30824
rect 7837 30815 7895 30821
rect 12710 30812 12716 30824
rect 12768 30812 12774 30864
rect 1210 30744 1216 30796
rect 1268 30784 1274 30796
rect 2685 30787 2743 30793
rect 2685 30784 2697 30787
rect 1268 30756 2697 30784
rect 1268 30744 1274 30756
rect 2685 30753 2697 30756
rect 2731 30753 2743 30787
rect 2685 30747 2743 30753
rect 6730 30744 6736 30796
rect 6788 30784 6794 30796
rect 11698 30784 11704 30796
rect 6788 30756 9352 30784
rect 11659 30756 11704 30784
rect 6788 30744 6794 30756
rect 658 30676 664 30728
rect 716 30716 722 30728
rect 2593 30719 2651 30725
rect 2593 30716 2605 30719
rect 716 30688 2605 30716
rect 716 30676 722 30688
rect 2593 30685 2605 30688
rect 2639 30685 2651 30719
rect 3418 30716 3424 30728
rect 3379 30688 3424 30716
rect 2593 30679 2651 30685
rect 3418 30676 3424 30688
rect 3476 30676 3482 30728
rect 5074 30716 5080 30728
rect 5035 30688 5080 30716
rect 5074 30676 5080 30688
rect 5132 30676 5138 30728
rect 5810 30716 5816 30728
rect 5771 30688 5816 30716
rect 5810 30676 5816 30688
rect 5868 30676 5874 30728
rect 6454 30716 6460 30728
rect 6415 30688 6460 30716
rect 6454 30676 6460 30688
rect 6512 30676 6518 30728
rect 6638 30676 6644 30728
rect 6696 30716 6702 30728
rect 7745 30719 7803 30725
rect 7745 30716 7757 30719
rect 6696 30688 7757 30716
rect 6696 30676 6702 30688
rect 7745 30685 7757 30688
rect 7791 30685 7803 30719
rect 7745 30679 7803 30685
rect 9030 30676 9036 30728
rect 9088 30716 9094 30728
rect 9125 30719 9183 30725
rect 9125 30716 9137 30719
rect 9088 30688 9137 30716
rect 9088 30676 9094 30688
rect 9125 30685 9137 30688
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 1949 30651 2007 30657
rect 1949 30617 1961 30651
rect 1995 30648 2007 30651
rect 2130 30648 2136 30660
rect 1995 30620 2136 30648
rect 1995 30617 2007 30620
rect 1949 30611 2007 30617
rect 2130 30608 2136 30620
rect 2188 30608 2194 30660
rect 5534 30608 5540 30660
rect 5592 30648 5598 30660
rect 9217 30651 9275 30657
rect 9217 30648 9229 30651
rect 5592 30620 9229 30648
rect 5592 30608 5598 30620
rect 9217 30617 9229 30620
rect 9263 30617 9275 30651
rect 9324 30648 9352 30756
rect 11698 30744 11704 30756
rect 11756 30744 11762 30796
rect 19889 30787 19947 30793
rect 19889 30753 19901 30787
rect 19935 30784 19947 30787
rect 21358 30784 21364 30796
rect 19935 30756 21364 30784
rect 19935 30753 19947 30756
rect 19889 30747 19947 30753
rect 21358 30744 21364 30756
rect 21416 30744 21422 30796
rect 23017 30787 23075 30793
rect 23017 30784 23029 30787
rect 22066 30756 23029 30784
rect 9769 30719 9827 30725
rect 9769 30685 9781 30719
rect 9815 30716 9827 30719
rect 10410 30716 10416 30728
rect 9815 30688 10416 30716
rect 9815 30685 9827 30688
rect 9769 30679 9827 30685
rect 10410 30676 10416 30688
rect 10468 30676 10474 30728
rect 10962 30716 10968 30728
rect 10923 30688 10968 30716
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 12894 30676 12900 30728
rect 12952 30716 12958 30728
rect 13265 30719 13323 30725
rect 13265 30716 13277 30719
rect 12952 30688 13277 30716
rect 12952 30676 12958 30688
rect 13265 30685 13277 30688
rect 13311 30685 13323 30719
rect 15010 30716 15016 30728
rect 14971 30688 15016 30716
rect 13265 30679 13323 30685
rect 15010 30676 15016 30688
rect 15068 30676 15074 30728
rect 11793 30651 11851 30657
rect 11793 30648 11805 30651
rect 9324 30620 11805 30648
rect 9217 30611 9275 30617
rect 11793 30617 11805 30620
rect 11839 30617 11851 30651
rect 11793 30611 11851 30617
rect 12526 30608 12532 30660
rect 12584 30648 12590 30660
rect 12713 30651 12771 30657
rect 12713 30648 12725 30651
rect 12584 30620 12725 30648
rect 12584 30608 12590 30620
rect 12713 30617 12725 30620
rect 12759 30648 12771 30651
rect 12802 30648 12808 30660
rect 12759 30620 12808 30648
rect 12759 30617 12771 30620
rect 12713 30611 12771 30617
rect 12802 30608 12808 30620
rect 12860 30608 12866 30660
rect 15378 30608 15384 30660
rect 15436 30648 15442 30660
rect 15436 30620 19932 30648
rect 15436 30608 15442 30620
rect 2038 30580 2044 30592
rect 1999 30552 2044 30580
rect 2038 30540 2044 30552
rect 2096 30540 2102 30592
rect 2958 30540 2964 30592
rect 3016 30580 3022 30592
rect 3237 30583 3295 30589
rect 3237 30580 3249 30583
rect 3016 30552 3249 30580
rect 3016 30540 3022 30552
rect 3237 30549 3249 30552
rect 3283 30549 3295 30583
rect 4430 30580 4436 30592
rect 4391 30552 4436 30580
rect 3237 30543 3295 30549
rect 4430 30540 4436 30552
rect 4488 30540 4494 30592
rect 5166 30580 5172 30592
rect 5127 30552 5172 30580
rect 5166 30540 5172 30552
rect 5224 30540 5230 30592
rect 5905 30583 5963 30589
rect 5905 30549 5917 30583
rect 5951 30580 5963 30583
rect 6914 30580 6920 30592
rect 5951 30552 6920 30580
rect 5951 30549 5963 30552
rect 5905 30543 5963 30549
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 7098 30580 7104 30592
rect 7059 30552 7104 30580
rect 7098 30540 7104 30552
rect 7156 30540 7162 30592
rect 8386 30580 8392 30592
rect 8347 30552 8392 30580
rect 8386 30540 8392 30552
rect 8444 30540 8450 30592
rect 9490 30540 9496 30592
rect 9548 30580 9554 30592
rect 9861 30583 9919 30589
rect 9861 30580 9873 30583
rect 9548 30552 9873 30580
rect 9548 30540 9554 30552
rect 9861 30549 9873 30552
rect 9907 30549 9919 30583
rect 9861 30543 9919 30549
rect 11057 30583 11115 30589
rect 11057 30549 11069 30583
rect 11103 30580 11115 30583
rect 11238 30580 11244 30592
rect 11103 30552 11244 30580
rect 11103 30549 11115 30552
rect 11057 30543 11115 30549
rect 11238 30540 11244 30552
rect 11296 30540 11302 30592
rect 15105 30583 15163 30589
rect 15105 30549 15117 30583
rect 15151 30580 15163 30583
rect 18782 30580 18788 30592
rect 15151 30552 18788 30580
rect 15151 30549 15163 30552
rect 15105 30543 15163 30549
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 19904 30580 19932 30620
rect 19978 30608 19984 30660
rect 20036 30648 20042 30660
rect 20901 30651 20959 30657
rect 20036 30620 20081 30648
rect 20036 30608 20042 30620
rect 20901 30617 20913 30651
rect 20947 30648 20959 30651
rect 22066 30648 22094 30756
rect 23017 30753 23029 30756
rect 23063 30753 23075 30787
rect 23017 30747 23075 30753
rect 20947 30620 22094 30648
rect 22741 30651 22799 30657
rect 20947 30617 20959 30620
rect 20901 30611 20959 30617
rect 22741 30617 22753 30651
rect 22787 30617 22799 30651
rect 22741 30611 22799 30617
rect 20916 30580 20944 30611
rect 19904 30552 20944 30580
rect 22756 30580 22784 30611
rect 22830 30608 22836 30660
rect 22888 30648 22894 30660
rect 38102 30648 38108 30660
rect 22888 30620 22933 30648
rect 38063 30620 38108 30648
rect 22888 30608 22894 30620
rect 38102 30608 38108 30620
rect 38160 30608 38166 30660
rect 25314 30580 25320 30592
rect 22756 30552 25320 30580
rect 25314 30540 25320 30552
rect 25372 30540 25378 30592
rect 38194 30580 38200 30592
rect 38155 30552 38200 30580
rect 38194 30540 38200 30552
rect 38252 30540 38258 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 10686 30376 10692 30388
rect 8312 30348 10692 30376
rect 5166 30308 5172 30320
rect 3344 30280 5172 30308
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30209 1639 30243
rect 2682 30240 2688 30252
rect 2643 30212 2688 30240
rect 1581 30203 1639 30209
rect 1596 30172 1624 30203
rect 2682 30200 2688 30212
rect 2740 30200 2746 30252
rect 3344 30249 3372 30280
rect 5166 30268 5172 30280
rect 5224 30268 5230 30320
rect 8312 30308 8340 30348
rect 10686 30336 10692 30348
rect 10744 30336 10750 30388
rect 10778 30336 10784 30388
rect 10836 30336 10842 30388
rect 12618 30376 12624 30388
rect 11624 30348 12624 30376
rect 7208 30280 8340 30308
rect 3329 30243 3387 30249
rect 3329 30209 3341 30243
rect 3375 30209 3387 30243
rect 3970 30240 3976 30252
rect 3931 30212 3976 30240
rect 3329 30203 3387 30209
rect 3970 30200 3976 30212
rect 4028 30200 4034 30252
rect 5261 30243 5319 30249
rect 5261 30209 5273 30243
rect 5307 30240 5319 30243
rect 5534 30240 5540 30252
rect 5307 30212 5540 30240
rect 5307 30209 5319 30212
rect 5261 30203 5319 30209
rect 5534 30200 5540 30212
rect 5592 30200 5598 30252
rect 7208 30249 7236 30280
rect 8386 30268 8392 30320
rect 8444 30308 8450 30320
rect 8849 30311 8907 30317
rect 8849 30308 8861 30311
rect 8444 30280 8861 30308
rect 8444 30268 8450 30280
rect 8849 30277 8861 30280
rect 8895 30277 8907 30311
rect 8849 30271 8907 30277
rect 8938 30268 8944 30320
rect 8996 30308 9002 30320
rect 8996 30280 9041 30308
rect 8996 30268 9002 30280
rect 9214 30268 9220 30320
rect 9272 30308 9278 30320
rect 9950 30308 9956 30320
rect 9272 30280 9956 30308
rect 9272 30268 9278 30280
rect 9950 30268 9956 30280
rect 10008 30268 10014 30320
rect 10796 30308 10824 30336
rect 10520 30280 10824 30308
rect 7193 30243 7251 30249
rect 7193 30209 7205 30243
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 7653 30243 7711 30249
rect 7653 30209 7665 30243
rect 7699 30209 7711 30243
rect 7653 30203 7711 30209
rect 3421 30175 3479 30181
rect 1596 30144 2774 30172
rect 1762 30104 1768 30116
rect 1723 30076 1768 30104
rect 1762 30064 1768 30076
rect 1820 30064 1826 30116
rect 2746 30104 2774 30144
rect 3421 30141 3433 30175
rect 3467 30172 3479 30175
rect 4614 30172 4620 30184
rect 3467 30144 4620 30172
rect 3467 30141 3479 30144
rect 3421 30135 3479 30141
rect 4614 30132 4620 30144
rect 4672 30132 4678 30184
rect 5718 30172 5724 30184
rect 5679 30144 5724 30172
rect 5718 30132 5724 30144
rect 5776 30132 5782 30184
rect 7668 30172 7696 30203
rect 10134 30200 10140 30252
rect 10192 30246 10198 30252
rect 10313 30249 10371 30255
rect 10313 30246 10325 30249
rect 10192 30218 10325 30246
rect 10192 30200 10198 30218
rect 10313 30215 10325 30218
rect 10359 30215 10371 30249
rect 10313 30209 10371 30215
rect 10413 30243 10471 30249
rect 10413 30209 10425 30243
rect 10459 30240 10471 30243
rect 10520 30240 10548 30280
rect 10459 30212 10548 30240
rect 10459 30209 10471 30212
rect 10413 30203 10471 30209
rect 10594 30200 10600 30252
rect 10652 30240 10658 30252
rect 10965 30243 11023 30249
rect 10965 30240 10977 30243
rect 10652 30212 10977 30240
rect 10652 30200 10658 30212
rect 10965 30209 10977 30212
rect 11011 30240 11023 30243
rect 11624 30240 11652 30348
rect 12618 30336 12624 30348
rect 12676 30336 12682 30388
rect 16114 30376 16120 30388
rect 16075 30348 16120 30376
rect 16114 30336 16120 30348
rect 16172 30336 16178 30388
rect 13354 30308 13360 30320
rect 13315 30280 13360 30308
rect 13354 30268 13360 30280
rect 13412 30268 13418 30320
rect 13449 30311 13507 30317
rect 13449 30277 13461 30311
rect 13495 30308 13507 30311
rect 15565 30311 15623 30317
rect 15565 30308 15577 30311
rect 13495 30280 15577 30308
rect 13495 30277 13507 30280
rect 13449 30271 13507 30277
rect 15565 30277 15577 30280
rect 15611 30277 15623 30311
rect 18506 30308 18512 30320
rect 15565 30271 15623 30277
rect 16132 30280 18512 30308
rect 11882 30240 11888 30252
rect 11011 30212 11652 30240
rect 11843 30212 11888 30240
rect 11011 30209 11023 30212
rect 10965 30203 11023 30209
rect 11882 30200 11888 30212
rect 11940 30200 11946 30252
rect 12250 30200 12256 30252
rect 12308 30240 12314 30252
rect 12345 30243 12403 30249
rect 12345 30240 12357 30243
rect 12308 30212 12357 30240
rect 12308 30200 12314 30212
rect 12345 30209 12357 30212
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 14829 30243 14887 30249
rect 14829 30209 14841 30243
rect 14875 30240 14887 30243
rect 15473 30243 15531 30249
rect 14875 30212 15424 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 8846 30172 8852 30184
rect 7668 30144 8852 30172
rect 5077 30107 5135 30113
rect 5077 30104 5089 30107
rect 2746 30076 5089 30104
rect 5077 30073 5089 30076
rect 5123 30073 5135 30107
rect 7668 30104 7696 30144
rect 8846 30132 8852 30144
rect 8904 30132 8910 30184
rect 9214 30172 9220 30184
rect 9175 30144 9220 30172
rect 9214 30132 9220 30144
rect 9272 30132 9278 30184
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 12437 30175 12495 30181
rect 12437 30172 12449 30175
rect 9364 30144 12449 30172
rect 9364 30132 9370 30144
rect 12437 30141 12449 30144
rect 12483 30141 12495 30175
rect 12437 30135 12495 30141
rect 14366 30132 14372 30184
rect 14424 30172 14430 30184
rect 15396 30172 15424 30212
rect 15473 30209 15485 30243
rect 15519 30240 15531 30243
rect 16132 30240 16160 30280
rect 18506 30268 18512 30280
rect 18564 30268 18570 30320
rect 19613 30311 19671 30317
rect 19613 30277 19625 30311
rect 19659 30308 19671 30311
rect 20162 30308 20168 30320
rect 19659 30280 20168 30308
rect 19659 30277 19671 30280
rect 19613 30271 19671 30277
rect 20162 30268 20168 30280
rect 20220 30268 20226 30320
rect 21358 30308 21364 30320
rect 21319 30280 21364 30308
rect 21358 30268 21364 30280
rect 21416 30268 21422 30320
rect 22554 30308 22560 30320
rect 22515 30280 22560 30308
rect 22554 30268 22560 30280
rect 22612 30268 22618 30320
rect 16298 30240 16304 30252
rect 15519 30212 16160 30240
rect 16259 30212 16304 30240
rect 15519 30209 15531 30212
rect 15473 30203 15531 30209
rect 16298 30200 16304 30212
rect 16356 30200 16362 30252
rect 21266 30240 21272 30252
rect 21227 30212 21272 30240
rect 21266 30200 21272 30212
rect 21324 30200 21330 30252
rect 22373 30243 22431 30249
rect 22373 30209 22385 30243
rect 22419 30240 22431 30243
rect 27430 30240 27436 30252
rect 22419 30212 27436 30240
rect 22419 30209 22431 30212
rect 22373 30203 22431 30209
rect 27430 30200 27436 30212
rect 27488 30200 27494 30252
rect 16482 30172 16488 30184
rect 14424 30144 14469 30172
rect 15396 30144 16488 30172
rect 14424 30132 14430 30144
rect 16482 30132 16488 30144
rect 16540 30132 16546 30184
rect 18785 30175 18843 30181
rect 18785 30141 18797 30175
rect 18831 30172 18843 30175
rect 19521 30175 19579 30181
rect 19521 30172 19533 30175
rect 18831 30144 19533 30172
rect 18831 30141 18843 30144
rect 18785 30135 18843 30141
rect 19521 30141 19533 30144
rect 19567 30141 19579 30175
rect 19521 30135 19579 30141
rect 19797 30175 19855 30181
rect 19797 30141 19809 30175
rect 19843 30172 19855 30175
rect 22094 30172 22100 30184
rect 19843 30144 22100 30172
rect 19843 30141 19855 30144
rect 19797 30135 19855 30141
rect 5077 30067 5135 30073
rect 5184 30076 7696 30104
rect 1670 29996 1676 30048
rect 1728 30036 1734 30048
rect 2777 30039 2835 30045
rect 2777 30036 2789 30039
rect 1728 30008 2789 30036
rect 1728 29996 1734 30008
rect 2777 30005 2789 30008
rect 2823 30005 2835 30039
rect 2777 29999 2835 30005
rect 3326 29996 3332 30048
rect 3384 30036 3390 30048
rect 4065 30039 4123 30045
rect 4065 30036 4077 30039
rect 3384 30008 4077 30036
rect 3384 29996 3390 30008
rect 4065 30005 4077 30008
rect 4111 30005 4123 30039
rect 4065 29999 4123 30005
rect 4154 29996 4160 30048
rect 4212 30036 4218 30048
rect 5184 30036 5212 30076
rect 8754 30064 8760 30116
rect 8812 30104 8818 30116
rect 8812 30076 12112 30104
rect 8812 30064 8818 30076
rect 7006 30036 7012 30048
rect 4212 30008 5212 30036
rect 6967 30008 7012 30036
rect 4212 29996 4218 30008
rect 7006 29996 7012 30008
rect 7064 29996 7070 30048
rect 7742 30036 7748 30048
rect 7703 30008 7748 30036
rect 7742 29996 7748 30008
rect 7800 29996 7806 30048
rect 8110 29996 8116 30048
rect 8168 30036 8174 30048
rect 11057 30039 11115 30045
rect 11057 30036 11069 30039
rect 8168 30008 11069 30036
rect 8168 29996 8174 30008
rect 11057 30005 11069 30008
rect 11103 30005 11115 30039
rect 11698 30036 11704 30048
rect 11659 30008 11704 30036
rect 11057 29999 11115 30005
rect 11698 29996 11704 30008
rect 11756 29996 11762 30048
rect 12084 30036 12112 30076
rect 12526 30036 12532 30048
rect 12084 30008 12532 30036
rect 12526 29996 12532 30008
rect 12584 29996 12590 30048
rect 12618 29996 12624 30048
rect 12676 30036 12682 30048
rect 14734 30036 14740 30048
rect 12676 30008 14740 30036
rect 12676 29996 12682 30008
rect 14734 29996 14740 30008
rect 14792 29996 14798 30048
rect 14918 30036 14924 30048
rect 14879 30008 14924 30036
rect 14918 29996 14924 30008
rect 14976 29996 14982 30048
rect 15470 29996 15476 30048
rect 15528 30036 15534 30048
rect 19812 30036 19840 30135
rect 22094 30132 22100 30144
rect 22152 30132 22158 30184
rect 15528 30008 19840 30036
rect 15528 29996 15534 30008
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 2685 29835 2743 29841
rect 2685 29801 2697 29835
rect 2731 29832 2743 29835
rect 7558 29832 7564 29844
rect 2731 29804 7564 29832
rect 2731 29801 2743 29804
rect 2685 29795 2743 29801
rect 7558 29792 7564 29804
rect 7616 29792 7622 29844
rect 8202 29792 8208 29844
rect 8260 29832 8266 29844
rect 8260 29804 14320 29832
rect 8260 29792 8266 29804
rect 11698 29764 11704 29776
rect 1596 29736 11704 29764
rect 1596 29637 1624 29736
rect 11698 29724 11704 29736
rect 11756 29724 11762 29776
rect 11790 29724 11796 29776
rect 11848 29764 11854 29776
rect 13906 29764 13912 29776
rect 11848 29736 13912 29764
rect 11848 29724 11854 29736
rect 13906 29724 13912 29736
rect 13964 29724 13970 29776
rect 6178 29656 6184 29708
rect 6236 29696 6242 29708
rect 9766 29696 9772 29708
rect 6236 29668 9772 29696
rect 6236 29656 6242 29668
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 10502 29656 10508 29708
rect 10560 29696 10566 29708
rect 11054 29696 11060 29708
rect 10560 29668 10605 29696
rect 11015 29668 11060 29696
rect 10560 29656 10566 29668
rect 11054 29656 11060 29668
rect 11112 29656 11118 29708
rect 12434 29656 12440 29708
rect 12492 29696 12498 29708
rect 12894 29696 12900 29708
rect 12492 29668 12537 29696
rect 12855 29668 12900 29696
rect 12492 29656 12498 29668
rect 12894 29656 12900 29668
rect 12952 29656 12958 29708
rect 14292 29696 14320 29804
rect 14366 29792 14372 29844
rect 14424 29832 14430 29844
rect 15378 29832 15384 29844
rect 14424 29804 15384 29832
rect 14424 29792 14430 29804
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 15562 29792 15568 29844
rect 15620 29832 15626 29844
rect 16393 29835 16451 29841
rect 16393 29832 16405 29835
rect 15620 29804 16405 29832
rect 15620 29792 15626 29804
rect 16393 29801 16405 29804
rect 16439 29801 16451 29835
rect 16393 29795 16451 29801
rect 18690 29792 18696 29844
rect 18748 29832 18754 29844
rect 22097 29835 22155 29841
rect 18748 29804 21036 29832
rect 18748 29792 18754 29804
rect 15286 29724 15292 29776
rect 15344 29764 15350 29776
rect 20073 29767 20131 29773
rect 20073 29764 20085 29767
rect 15344 29736 20085 29764
rect 15344 29724 15350 29736
rect 20073 29733 20085 29736
rect 20119 29764 20131 29767
rect 20714 29764 20720 29776
rect 20119 29736 20720 29764
rect 20119 29733 20131 29736
rect 20073 29727 20131 29733
rect 20714 29724 20720 29736
rect 20772 29724 20778 29776
rect 18322 29696 18328 29708
rect 14292 29668 18328 29696
rect 18322 29656 18328 29668
rect 18380 29656 18386 29708
rect 18874 29656 18880 29708
rect 18932 29696 18938 29708
rect 20809 29699 20867 29705
rect 20809 29696 20821 29699
rect 18932 29668 20821 29696
rect 18932 29656 18938 29668
rect 20809 29665 20821 29668
rect 20855 29665 20867 29699
rect 20809 29659 20867 29665
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29597 1639 29631
rect 2590 29628 2596 29640
rect 2551 29600 2596 29628
rect 1581 29591 1639 29597
rect 2590 29588 2596 29600
rect 2648 29588 2654 29640
rect 3237 29631 3295 29637
rect 3237 29597 3249 29631
rect 3283 29628 3295 29631
rect 4062 29628 4068 29640
rect 3283 29600 4068 29628
rect 3283 29597 3295 29600
rect 3237 29591 3295 29597
rect 4062 29588 4068 29600
rect 4120 29588 4126 29640
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29628 4583 29631
rect 4798 29628 4804 29640
rect 4571 29600 4804 29628
rect 4571 29597 4583 29600
rect 4525 29591 4583 29597
rect 4798 29588 4804 29600
rect 4856 29628 4862 29640
rect 5169 29631 5227 29637
rect 5169 29628 5181 29631
rect 4856 29600 5181 29628
rect 4856 29588 4862 29600
rect 5169 29597 5181 29600
rect 5215 29628 5227 29631
rect 5813 29631 5871 29637
rect 5813 29628 5825 29631
rect 5215 29600 5825 29628
rect 5215 29597 5227 29600
rect 5169 29591 5227 29597
rect 5813 29597 5825 29600
rect 5859 29597 5871 29631
rect 5813 29591 5871 29597
rect 6086 29588 6092 29640
rect 6144 29628 6150 29640
rect 6457 29631 6515 29637
rect 6457 29628 6469 29631
rect 6144 29600 6469 29628
rect 6144 29588 6150 29600
rect 6457 29597 6469 29600
rect 6503 29628 6515 29631
rect 7101 29631 7159 29637
rect 7101 29628 7113 29631
rect 6503 29600 7113 29628
rect 6503 29597 6515 29600
rect 6457 29591 6515 29597
rect 7101 29597 7113 29600
rect 7147 29628 7159 29631
rect 7745 29631 7803 29637
rect 7745 29628 7757 29631
rect 7147 29600 7757 29628
rect 7147 29597 7159 29600
rect 7101 29591 7159 29597
rect 7745 29597 7757 29600
rect 7791 29597 7803 29631
rect 7745 29591 7803 29597
rect 8389 29631 8447 29637
rect 8389 29597 8401 29631
rect 8435 29628 8447 29631
rect 8662 29628 8668 29640
rect 8435 29600 8668 29628
rect 8435 29597 8447 29600
rect 8389 29591 8447 29597
rect 3602 29520 3608 29572
rect 3660 29560 3666 29572
rect 4617 29563 4675 29569
rect 4617 29560 4629 29563
rect 3660 29532 4629 29560
rect 3660 29520 3666 29532
rect 4617 29529 4629 29532
rect 4663 29529 4675 29563
rect 4617 29523 4675 29529
rect 4982 29520 4988 29572
rect 5040 29560 5046 29572
rect 6549 29563 6607 29569
rect 6549 29560 6561 29563
rect 5040 29532 6561 29560
rect 5040 29520 5046 29532
rect 6549 29529 6561 29532
rect 6595 29529 6607 29563
rect 7760 29560 7788 29591
rect 8662 29588 8668 29600
rect 8720 29588 8726 29640
rect 8754 29588 8760 29640
rect 8812 29628 8818 29640
rect 9125 29631 9183 29637
rect 9125 29628 9137 29631
rect 8812 29600 9137 29628
rect 8812 29588 8818 29600
rect 9125 29597 9137 29600
rect 9171 29597 9183 29631
rect 9125 29591 9183 29597
rect 9953 29630 10011 29633
rect 9953 29628 10088 29630
rect 10134 29628 10140 29640
rect 9953 29627 10140 29628
rect 9953 29593 9965 29627
rect 9999 29602 10140 29627
rect 9999 29593 10011 29602
rect 10060 29600 10140 29602
rect 9953 29587 10011 29593
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 14550 29628 14556 29640
rect 14511 29600 14556 29628
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 15657 29631 15715 29637
rect 15657 29628 15669 29631
rect 14792 29600 15669 29628
rect 14792 29588 14798 29600
rect 15657 29597 15669 29600
rect 15703 29597 15715 29631
rect 15657 29591 15715 29597
rect 16301 29631 16359 29637
rect 16301 29597 16313 29631
rect 16347 29628 16359 29631
rect 16482 29628 16488 29640
rect 16347 29600 16488 29628
rect 16347 29597 16359 29600
rect 16301 29591 16359 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 18690 29628 18696 29640
rect 18651 29600 18696 29628
rect 18690 29588 18696 29600
rect 18748 29588 18754 29640
rect 20717 29631 20775 29637
rect 20717 29597 20729 29631
rect 20763 29628 20775 29631
rect 20898 29628 20904 29640
rect 20763 29600 20904 29628
rect 20763 29597 20775 29600
rect 20717 29591 20775 29597
rect 20898 29588 20904 29600
rect 20956 29588 20962 29640
rect 21008 29628 21036 29804
rect 22097 29801 22109 29835
rect 22143 29832 22155 29835
rect 22830 29832 22836 29844
rect 22143 29804 22836 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 26145 29835 26203 29841
rect 26145 29801 26157 29835
rect 26191 29832 26203 29835
rect 27798 29832 27804 29844
rect 26191 29804 27804 29832
rect 26191 29801 26203 29804
rect 26145 29795 26203 29801
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 22005 29631 22063 29637
rect 22005 29628 22017 29631
rect 21008 29600 22017 29628
rect 22005 29597 22017 29600
rect 22051 29597 22063 29631
rect 22005 29591 22063 29597
rect 24486 29588 24492 29640
rect 24544 29628 24550 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 24544 29600 24593 29628
rect 24544 29588 24550 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 26050 29628 26056 29640
rect 26011 29600 26056 29628
rect 24581 29591 24639 29597
rect 26050 29588 26056 29600
rect 26108 29588 26114 29640
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29628 26755 29631
rect 26970 29628 26976 29640
rect 26743 29600 26976 29628
rect 26743 29597 26755 29600
rect 26697 29591 26755 29597
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 38286 29628 38292 29640
rect 38247 29600 38292 29628
rect 38286 29588 38292 29600
rect 38344 29588 38350 29640
rect 9858 29560 9864 29572
rect 7760 29532 9864 29560
rect 6549 29523 6607 29529
rect 9858 29520 9864 29532
rect 9916 29520 9922 29572
rect 10594 29520 10600 29572
rect 10652 29569 10658 29572
rect 10652 29560 10664 29569
rect 10652 29532 10697 29560
rect 10652 29523 10664 29532
rect 10652 29520 10658 29523
rect 10778 29520 10784 29572
rect 10836 29560 10842 29572
rect 12529 29563 12587 29569
rect 12529 29560 12541 29563
rect 10836 29532 12541 29560
rect 10836 29520 10842 29532
rect 12529 29529 12541 29532
rect 12575 29529 12587 29563
rect 12529 29523 12587 29529
rect 12618 29520 12624 29572
rect 12676 29560 12682 29572
rect 14274 29560 14280 29572
rect 12676 29532 14280 29560
rect 12676 29520 12682 29532
rect 14274 29520 14280 29532
rect 14332 29520 14338 29572
rect 19518 29560 19524 29572
rect 19479 29532 19524 29560
rect 19518 29520 19524 29532
rect 19576 29520 19582 29572
rect 19613 29563 19671 29569
rect 19613 29529 19625 29563
rect 19659 29529 19671 29563
rect 19613 29523 19671 29529
rect 1762 29492 1768 29504
rect 1723 29464 1768 29492
rect 1762 29452 1768 29464
rect 1820 29452 1826 29504
rect 3329 29495 3387 29501
rect 3329 29461 3341 29495
rect 3375 29492 3387 29495
rect 3786 29492 3792 29504
rect 3375 29464 3792 29492
rect 3375 29461 3387 29464
rect 3329 29455 3387 29461
rect 3786 29452 3792 29464
rect 3844 29452 3850 29504
rect 5261 29495 5319 29501
rect 5261 29461 5273 29495
rect 5307 29492 5319 29495
rect 5350 29492 5356 29504
rect 5307 29464 5356 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 5350 29452 5356 29464
rect 5408 29452 5414 29504
rect 5905 29495 5963 29501
rect 5905 29461 5917 29495
rect 5951 29492 5963 29495
rect 6362 29492 6368 29504
rect 5951 29464 6368 29492
rect 5951 29461 5963 29464
rect 5905 29455 5963 29461
rect 6362 29452 6368 29464
rect 6420 29452 6426 29504
rect 7193 29495 7251 29501
rect 7193 29461 7205 29495
rect 7239 29492 7251 29495
rect 7466 29492 7472 29504
rect 7239 29464 7472 29492
rect 7239 29461 7251 29464
rect 7193 29455 7251 29461
rect 7466 29452 7472 29464
rect 7524 29452 7530 29504
rect 7834 29492 7840 29504
rect 7795 29464 7840 29492
rect 7834 29452 7840 29464
rect 7892 29452 7898 29504
rect 7926 29452 7932 29504
rect 7984 29492 7990 29504
rect 8481 29495 8539 29501
rect 8481 29492 8493 29495
rect 7984 29464 8493 29492
rect 7984 29452 7990 29464
rect 8481 29461 8493 29464
rect 8527 29461 8539 29495
rect 8481 29455 8539 29461
rect 9122 29452 9128 29504
rect 9180 29492 9186 29504
rect 9217 29495 9275 29501
rect 9217 29492 9229 29495
rect 9180 29464 9229 29492
rect 9180 29452 9186 29464
rect 9217 29461 9229 29464
rect 9263 29461 9275 29495
rect 9766 29492 9772 29504
rect 9727 29464 9772 29492
rect 9217 29455 9275 29461
rect 9766 29452 9772 29464
rect 9824 29452 9830 29504
rect 14458 29452 14464 29504
rect 14516 29492 14522 29504
rect 14645 29495 14703 29501
rect 14645 29492 14657 29495
rect 14516 29464 14657 29492
rect 14516 29452 14522 29464
rect 14645 29461 14657 29464
rect 14691 29461 14703 29495
rect 15746 29492 15752 29504
rect 15707 29464 15752 29492
rect 14645 29455 14703 29461
rect 15746 29452 15752 29464
rect 15804 29452 15810 29504
rect 18785 29495 18843 29501
rect 18785 29461 18797 29495
rect 18831 29492 18843 29495
rect 19628 29492 19656 29523
rect 18831 29464 19656 29492
rect 23753 29495 23811 29501
rect 18831 29461 18843 29464
rect 18785 29455 18843 29461
rect 23753 29461 23765 29495
rect 23799 29492 23811 29495
rect 23934 29492 23940 29504
rect 23799 29464 23940 29492
rect 23799 29461 23811 29464
rect 23753 29455 23811 29461
rect 23934 29452 23940 29464
rect 23992 29452 23998 29504
rect 24026 29452 24032 29504
rect 24084 29492 24090 29504
rect 24673 29495 24731 29501
rect 24673 29492 24685 29495
rect 24084 29464 24685 29492
rect 24084 29452 24090 29464
rect 24673 29461 24685 29464
rect 24719 29461 24731 29495
rect 24673 29455 24731 29461
rect 26510 29452 26516 29504
rect 26568 29492 26574 29504
rect 26789 29495 26847 29501
rect 26789 29492 26801 29495
rect 26568 29464 26801 29492
rect 26568 29452 26574 29464
rect 26789 29461 26801 29464
rect 26835 29461 26847 29495
rect 26789 29455 26847 29461
rect 36998 29452 37004 29504
rect 37056 29492 37062 29504
rect 38105 29495 38163 29501
rect 38105 29492 38117 29495
rect 37056 29464 38117 29492
rect 37056 29452 37062 29464
rect 38105 29461 38117 29464
rect 38151 29461 38163 29495
rect 38105 29455 38163 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 566 29248 572 29300
rect 624 29288 630 29300
rect 8389 29291 8447 29297
rect 624 29260 7788 29288
rect 624 29248 630 29260
rect 2130 29180 2136 29232
rect 2188 29220 2194 29232
rect 2188 29192 5764 29220
rect 2188 29180 2194 29192
rect 1857 29155 1915 29161
rect 1857 29121 1869 29155
rect 1903 29152 1915 29155
rect 2406 29152 2412 29164
rect 1903 29124 2412 29152
rect 1903 29121 1915 29124
rect 1857 29115 1915 29121
rect 2406 29112 2412 29124
rect 2464 29112 2470 29164
rect 2501 29155 2559 29161
rect 2501 29121 2513 29155
rect 2547 29152 2559 29155
rect 2866 29152 2872 29164
rect 2547 29124 2872 29152
rect 2547 29121 2559 29124
rect 2501 29115 2559 29121
rect 2866 29112 2872 29124
rect 2924 29152 2930 29164
rect 3237 29155 3295 29161
rect 3237 29152 3249 29155
rect 2924 29124 3249 29152
rect 2924 29112 2930 29124
rect 3237 29121 3249 29124
rect 3283 29152 3295 29155
rect 3878 29152 3884 29164
rect 3283 29124 3884 29152
rect 3283 29121 3295 29124
rect 3237 29115 3295 29121
rect 3878 29112 3884 29124
rect 3936 29112 3942 29164
rect 3973 29155 4031 29161
rect 3973 29121 3985 29155
rect 4019 29121 4031 29155
rect 3973 29115 4031 29121
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29152 4675 29155
rect 5074 29152 5080 29164
rect 4663 29124 5080 29152
rect 4663 29121 4675 29124
rect 4617 29115 4675 29121
rect 1949 29087 2007 29093
rect 1949 29053 1961 29087
rect 1995 29084 2007 29087
rect 2774 29084 2780 29096
rect 1995 29056 2780 29084
rect 1995 29053 2007 29056
rect 1949 29047 2007 29053
rect 2774 29044 2780 29056
rect 2832 29044 2838 29096
rect 3988 29084 4016 29115
rect 5074 29112 5080 29124
rect 5132 29112 5138 29164
rect 5736 29161 5764 29192
rect 7190 29180 7196 29232
rect 7248 29220 7254 29232
rect 7650 29220 7656 29232
rect 7248 29192 7656 29220
rect 7248 29180 7254 29192
rect 7650 29180 7656 29192
rect 7708 29180 7714 29232
rect 7760 29220 7788 29260
rect 8389 29257 8401 29291
rect 8435 29288 8447 29291
rect 8938 29288 8944 29300
rect 8435 29260 8944 29288
rect 8435 29257 8447 29260
rect 8389 29251 8447 29257
rect 8938 29248 8944 29260
rect 8996 29248 9002 29300
rect 9493 29291 9551 29297
rect 9493 29257 9505 29291
rect 9539 29288 9551 29291
rect 11790 29288 11796 29300
rect 9539 29260 11796 29288
rect 9539 29257 9551 29260
rect 9493 29251 9551 29257
rect 11790 29248 11796 29260
rect 11848 29248 11854 29300
rect 11900 29260 12940 29288
rect 9306 29220 9312 29232
rect 7760 29192 9312 29220
rect 9306 29180 9312 29192
rect 9364 29180 9370 29232
rect 10226 29220 10232 29232
rect 10187 29192 10232 29220
rect 10226 29180 10232 29192
rect 10284 29180 10290 29232
rect 5721 29155 5779 29161
rect 5721 29121 5733 29155
rect 5767 29121 5779 29155
rect 5721 29115 5779 29121
rect 6914 29112 6920 29164
rect 6972 29112 6978 29164
rect 7101 29155 7159 29161
rect 7101 29121 7113 29155
rect 7147 29152 7159 29155
rect 8202 29152 8208 29164
rect 7147 29124 8208 29152
rect 7147 29121 7159 29124
rect 7101 29115 7159 29121
rect 8202 29112 8208 29124
rect 8260 29112 8266 29164
rect 8294 29112 8300 29164
rect 8352 29152 8358 29164
rect 9398 29152 9404 29164
rect 8352 29124 8397 29152
rect 9359 29124 9404 29152
rect 8352 29112 8358 29124
rect 9398 29112 9404 29124
rect 9456 29112 9462 29164
rect 4798 29084 4804 29096
rect 3988 29056 4804 29084
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 5813 29087 5871 29093
rect 5813 29053 5825 29087
rect 5859 29084 5871 29087
rect 6822 29084 6828 29096
rect 5859 29056 6828 29084
rect 5859 29053 5871 29056
rect 5813 29047 5871 29053
rect 6822 29044 6828 29056
rect 6880 29044 6886 29096
rect 6932 29084 6960 29112
rect 10137 29087 10195 29093
rect 10137 29084 10149 29087
rect 6932 29056 10149 29084
rect 10137 29053 10149 29056
rect 10183 29053 10195 29087
rect 10778 29084 10784 29096
rect 10739 29056 10784 29084
rect 10137 29047 10195 29053
rect 10778 29044 10784 29056
rect 10836 29044 10842 29096
rect 1302 28976 1308 29028
rect 1360 29016 1366 29028
rect 2593 29019 2651 29025
rect 2593 29016 2605 29019
rect 1360 28988 2605 29016
rect 1360 28976 1366 28988
rect 2593 28985 2605 28988
rect 2639 28985 2651 29019
rect 2593 28979 2651 28985
rect 3142 28976 3148 29028
rect 3200 29016 3206 29028
rect 3329 29019 3387 29025
rect 3329 29016 3341 29019
rect 3200 28988 3341 29016
rect 3200 28976 3206 28988
rect 3329 28985 3341 28988
rect 3375 28985 3387 29019
rect 3329 28979 3387 28985
rect 3970 28976 3976 29028
rect 4028 29016 4034 29028
rect 4065 29019 4123 29025
rect 4065 29016 4077 29019
rect 4028 28988 4077 29016
rect 4028 28976 4034 28988
rect 4065 28985 4077 28988
rect 4111 28985 4123 29019
rect 4065 28979 4123 28985
rect 4709 29019 4767 29025
rect 4709 28985 4721 29019
rect 4755 29016 4767 29019
rect 6914 29016 6920 29028
rect 4755 28988 6920 29016
rect 4755 28985 4767 28988
rect 4709 28979 4767 28985
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 7190 29016 7196 29028
rect 7151 28988 7196 29016
rect 7190 28976 7196 28988
rect 7248 28976 7254 29028
rect 7558 28976 7564 29028
rect 7616 29016 7622 29028
rect 11900 29016 11928 29260
rect 12069 29223 12127 29229
rect 12069 29189 12081 29223
rect 12115 29220 12127 29223
rect 12805 29223 12863 29229
rect 12805 29220 12817 29223
rect 12115 29192 12817 29220
rect 12115 29189 12127 29192
rect 12069 29183 12127 29189
rect 12805 29189 12817 29192
rect 12851 29189 12863 29223
rect 12912 29220 12940 29260
rect 14274 29248 14280 29300
rect 14332 29288 14338 29300
rect 19518 29288 19524 29300
rect 14332 29260 19524 29288
rect 14332 29248 14338 29260
rect 19518 29248 19524 29260
rect 19576 29248 19582 29300
rect 14642 29220 14648 29232
rect 12912 29192 14648 29220
rect 12805 29183 12863 29189
rect 14642 29180 14648 29192
rect 14700 29180 14706 29232
rect 14737 29223 14795 29229
rect 14737 29189 14749 29223
rect 14783 29220 14795 29223
rect 15562 29220 15568 29232
rect 14783 29192 15568 29220
rect 14783 29189 14795 29192
rect 14737 29183 14795 29189
rect 15562 29180 15568 29192
rect 15620 29180 15626 29232
rect 18966 29220 18972 29232
rect 18927 29192 18972 29220
rect 18966 29180 18972 29192
rect 19024 29180 19030 29232
rect 19426 29180 19432 29232
rect 19484 29220 19490 29232
rect 20438 29220 20444 29232
rect 19484 29192 20444 29220
rect 19484 29180 19490 29192
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 20533 29223 20591 29229
rect 20533 29189 20545 29223
rect 20579 29220 20591 29223
rect 20622 29220 20628 29232
rect 20579 29192 20628 29220
rect 20579 29189 20591 29192
rect 20533 29183 20591 29189
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 23566 29220 23572 29232
rect 23527 29192 23572 29220
rect 23566 29180 23572 29192
rect 23624 29180 23630 29232
rect 23658 29180 23664 29232
rect 23716 29220 23722 29232
rect 23716 29192 23761 29220
rect 23716 29180 23722 29192
rect 23934 29180 23940 29232
rect 23992 29220 23998 29232
rect 25133 29223 25191 29229
rect 25133 29220 25145 29223
rect 23992 29192 25145 29220
rect 23992 29180 23998 29192
rect 25133 29189 25145 29192
rect 25179 29189 25191 29223
rect 25133 29183 25191 29189
rect 25222 29180 25228 29232
rect 25280 29220 25286 29232
rect 25280 29192 25325 29220
rect 25280 29180 25286 29192
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29152 12035 29155
rect 14366 29152 14372 29164
rect 12023 29124 12434 29152
rect 12023 29121 12035 29124
rect 11977 29115 12035 29121
rect 7616 28988 11928 29016
rect 12406 29016 12434 29124
rect 13556 29124 14372 29152
rect 12710 29084 12716 29096
rect 12671 29056 12716 29084
rect 12710 29044 12716 29056
rect 12768 29044 12774 29096
rect 13556 29084 13584 29124
rect 14366 29112 14372 29124
rect 14424 29112 14430 29164
rect 15286 29112 15292 29164
rect 15344 29152 15350 29164
rect 15344 29124 15389 29152
rect 15344 29112 15350 29124
rect 15654 29112 15660 29164
rect 15712 29152 15718 29164
rect 15749 29155 15807 29161
rect 15749 29152 15761 29155
rect 15712 29124 15761 29152
rect 15712 29112 15718 29124
rect 15749 29121 15761 29124
rect 15795 29121 15807 29155
rect 15749 29115 15807 29121
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29152 15899 29155
rect 15930 29152 15936 29164
rect 15887 29124 15936 29152
rect 15887 29121 15899 29124
rect 15841 29115 15899 29121
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 16850 29152 16856 29164
rect 16811 29124 16856 29152
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 18141 29155 18199 29161
rect 18141 29121 18153 29155
rect 18187 29121 18199 29155
rect 18141 29115 18199 29121
rect 12820 29056 13584 29084
rect 12820 29016 12848 29056
rect 13630 29044 13636 29096
rect 13688 29084 13694 29096
rect 13688 29056 13733 29084
rect 13688 29044 13694 29056
rect 13906 29044 13912 29096
rect 13964 29084 13970 29096
rect 14645 29087 14703 29093
rect 14645 29084 14657 29087
rect 13964 29056 14657 29084
rect 13964 29044 13970 29056
rect 14645 29053 14657 29056
rect 14691 29053 14703 29087
rect 18156 29084 18184 29115
rect 18874 29084 18880 29096
rect 14645 29047 14703 29053
rect 14752 29056 18184 29084
rect 18835 29056 18880 29084
rect 12406 28988 12848 29016
rect 7616 28976 7622 28988
rect 13078 28976 13084 29028
rect 13136 29016 13142 29028
rect 14752 29016 14780 29056
rect 18874 29044 18880 29056
rect 18932 29044 18938 29096
rect 19334 29084 19340 29096
rect 19295 29056 19340 29084
rect 19334 29044 19340 29056
rect 19392 29044 19398 29096
rect 21082 29084 21088 29096
rect 21043 29056 21088 29084
rect 21082 29044 21088 29056
rect 21140 29044 21146 29096
rect 23934 29084 23940 29096
rect 23895 29056 23940 29084
rect 23934 29044 23940 29056
rect 23992 29044 23998 29096
rect 25409 29087 25467 29093
rect 25409 29053 25421 29087
rect 25455 29084 25467 29087
rect 26050 29084 26056 29096
rect 25455 29056 26056 29084
rect 25455 29053 25467 29056
rect 25409 29047 25467 29053
rect 16945 29019 17003 29025
rect 16945 29016 16957 29019
rect 13136 28988 14780 29016
rect 15304 28988 16957 29016
rect 13136 28976 13142 28988
rect 1578 28908 1584 28960
rect 1636 28948 1642 28960
rect 9766 28948 9772 28960
rect 1636 28920 9772 28948
rect 1636 28908 1642 28920
rect 9766 28908 9772 28920
rect 9824 28908 9830 28960
rect 13814 28908 13820 28960
rect 13872 28948 13878 28960
rect 15304 28948 15332 28988
rect 16945 28985 16957 28988
rect 16991 28985 17003 29019
rect 16945 28979 17003 28985
rect 18322 28976 18328 29028
rect 18380 29016 18386 29028
rect 18380 28988 19288 29016
rect 18380 28976 18386 28988
rect 13872 28920 15332 28948
rect 18233 28951 18291 28957
rect 13872 28908 13878 28920
rect 18233 28917 18245 28951
rect 18279 28948 18291 28951
rect 18598 28948 18604 28960
rect 18279 28920 18604 28948
rect 18279 28917 18291 28920
rect 18233 28911 18291 28917
rect 18598 28908 18604 28920
rect 18656 28908 18662 28960
rect 19260 28948 19288 28988
rect 19978 28976 19984 29028
rect 20036 29016 20042 29028
rect 25424 29016 25452 29047
rect 26050 29044 26056 29056
rect 26108 29044 26114 29096
rect 37182 29044 37188 29096
rect 37240 29084 37246 29096
rect 37461 29087 37519 29093
rect 37461 29084 37473 29087
rect 37240 29056 37473 29084
rect 37240 29044 37246 29056
rect 37461 29053 37473 29056
rect 37507 29053 37519 29087
rect 37461 29047 37519 29053
rect 37737 29087 37795 29093
rect 37737 29053 37749 29087
rect 37783 29053 37795 29087
rect 37737 29047 37795 29053
rect 20036 28988 25452 29016
rect 20036 28976 20042 28988
rect 27430 28976 27436 29028
rect 27488 29016 27494 29028
rect 37752 29016 37780 29047
rect 27488 28988 37780 29016
rect 27488 28976 27494 28988
rect 20806 28948 20812 28960
rect 19260 28920 20812 28948
rect 20806 28908 20812 28920
rect 20864 28908 20870 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 5166 28704 5172 28756
rect 5224 28744 5230 28756
rect 5224 28716 14504 28744
rect 5224 28704 5230 28716
rect 2590 28636 2596 28688
rect 2648 28676 2654 28688
rect 6086 28676 6092 28688
rect 2648 28648 6092 28676
rect 2648 28636 2654 28648
rect 6086 28636 6092 28648
rect 6144 28636 6150 28688
rect 9398 28676 9404 28688
rect 6840 28648 9404 28676
rect 2746 28580 4660 28608
rect 1946 28540 1952 28552
rect 1907 28512 1952 28540
rect 1946 28500 1952 28512
rect 2004 28500 2010 28552
rect 2593 28543 2651 28549
rect 2593 28509 2605 28543
rect 2639 28540 2651 28543
rect 2746 28540 2774 28580
rect 2639 28512 2774 28540
rect 3237 28543 3295 28549
rect 2639 28509 2651 28512
rect 2593 28503 2651 28509
rect 3237 28509 3249 28543
rect 3283 28509 3295 28543
rect 3237 28503 3295 28509
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28540 4031 28543
rect 4062 28540 4068 28552
rect 4019 28512 4068 28540
rect 4019 28509 4031 28512
rect 3973 28503 4031 28509
rect 3252 28472 3280 28503
rect 4062 28500 4068 28512
rect 4120 28500 4126 28552
rect 4632 28549 4660 28580
rect 4617 28543 4675 28549
rect 4617 28509 4629 28543
rect 4663 28540 4675 28543
rect 4890 28540 4896 28552
rect 4663 28512 4896 28540
rect 4663 28509 4675 28512
rect 4617 28503 4675 28509
rect 4890 28500 4896 28512
rect 4948 28540 4954 28552
rect 6104 28549 6132 28636
rect 6840 28549 6868 28648
rect 9398 28636 9404 28648
rect 9456 28636 9462 28688
rect 7837 28611 7895 28617
rect 7837 28577 7849 28611
rect 7883 28608 7895 28611
rect 10870 28608 10876 28620
rect 7883 28580 10876 28608
rect 7883 28577 7895 28580
rect 7837 28571 7895 28577
rect 10870 28568 10876 28580
rect 10928 28568 10934 28620
rect 14476 28608 14504 28716
rect 16850 28704 16856 28756
rect 16908 28744 16914 28756
rect 18785 28747 18843 28753
rect 16908 28716 17724 28744
rect 16908 28704 16914 28716
rect 15194 28636 15200 28688
rect 15252 28676 15258 28688
rect 17589 28679 17647 28685
rect 17589 28676 17601 28679
rect 15252 28648 17601 28676
rect 15252 28636 15258 28648
rect 17589 28645 17601 28648
rect 17635 28645 17647 28679
rect 17696 28676 17724 28716
rect 18785 28713 18797 28747
rect 18831 28744 18843 28747
rect 18966 28744 18972 28756
rect 18831 28716 18972 28744
rect 18831 28713 18843 28716
rect 18785 28707 18843 28713
rect 18966 28704 18972 28716
rect 19024 28704 19030 28756
rect 20070 28704 20076 28756
rect 20128 28744 20134 28756
rect 20165 28747 20223 28753
rect 20165 28744 20177 28747
rect 20128 28716 20177 28744
rect 20128 28704 20134 28716
rect 20165 28713 20177 28716
rect 20211 28713 20223 28747
rect 20165 28707 20223 28713
rect 23382 28704 23388 28756
rect 23440 28744 23446 28756
rect 24581 28747 24639 28753
rect 24581 28744 24593 28747
rect 23440 28716 24593 28744
rect 23440 28704 23446 28716
rect 24581 28713 24593 28716
rect 24627 28713 24639 28747
rect 26878 28744 26884 28756
rect 26839 28716 26884 28744
rect 24581 28707 24639 28713
rect 26878 28704 26884 28716
rect 26936 28704 26942 28756
rect 19058 28676 19064 28688
rect 17696 28648 19064 28676
rect 17589 28639 17647 28645
rect 19058 28636 19064 28648
rect 19116 28636 19122 28688
rect 20254 28636 20260 28688
rect 20312 28676 20318 28688
rect 21910 28676 21916 28688
rect 20312 28648 21916 28676
rect 20312 28636 20318 28648
rect 21910 28636 21916 28648
rect 21968 28636 21974 28688
rect 23477 28679 23535 28685
rect 23477 28645 23489 28679
rect 23523 28676 23535 28679
rect 32398 28676 32404 28688
rect 23523 28648 32404 28676
rect 23523 28645 23535 28648
rect 23477 28639 23535 28645
rect 32398 28636 32404 28648
rect 32456 28636 32462 28688
rect 24302 28608 24308 28620
rect 14476 28580 24308 28608
rect 24302 28568 24308 28580
rect 24360 28568 24366 28620
rect 25314 28608 25320 28620
rect 25275 28580 25320 28608
rect 25314 28568 25320 28580
rect 25372 28568 25378 28620
rect 25498 28568 25504 28620
rect 25556 28608 25562 28620
rect 25593 28611 25651 28617
rect 25593 28608 25605 28611
rect 25556 28580 25605 28608
rect 25556 28568 25562 28580
rect 25593 28577 25605 28580
rect 25639 28577 25651 28611
rect 25593 28571 25651 28577
rect 5261 28543 5319 28549
rect 5261 28540 5273 28543
rect 4948 28512 5273 28540
rect 4948 28500 4954 28512
rect 5261 28509 5273 28512
rect 5307 28509 5319 28543
rect 5261 28503 5319 28509
rect 6089 28543 6147 28549
rect 6089 28509 6101 28543
rect 6135 28509 6147 28543
rect 6089 28503 6147 28509
rect 6825 28543 6883 28549
rect 6825 28509 6837 28543
rect 6871 28509 6883 28543
rect 6825 28503 6883 28509
rect 7558 28500 7564 28552
rect 7616 28540 7622 28552
rect 7745 28543 7803 28549
rect 7745 28540 7757 28543
rect 7616 28512 7757 28540
rect 7616 28500 7622 28512
rect 7745 28509 7757 28512
rect 7791 28509 7803 28543
rect 7745 28503 7803 28509
rect 8389 28543 8447 28549
rect 8389 28509 8401 28543
rect 8435 28540 8447 28543
rect 9217 28543 9275 28549
rect 8435 28512 9168 28540
rect 8435 28509 8447 28512
rect 8389 28503 8447 28509
rect 6546 28472 6552 28484
rect 3252 28444 6552 28472
rect 6546 28432 6552 28444
rect 6604 28432 6610 28484
rect 7006 28472 7012 28484
rect 6967 28444 7012 28472
rect 7006 28432 7012 28444
rect 7064 28432 7070 28484
rect 8294 28432 8300 28484
rect 8352 28472 8358 28484
rect 9140 28472 9168 28512
rect 9217 28509 9229 28543
rect 9263 28540 9275 28543
rect 9398 28540 9404 28552
rect 9263 28512 9404 28540
rect 9263 28509 9275 28512
rect 9217 28503 9275 28509
rect 9398 28500 9404 28512
rect 9456 28540 9462 28552
rect 9858 28540 9864 28552
rect 9456 28512 9864 28540
rect 9456 28500 9462 28512
rect 9858 28500 9864 28512
rect 9916 28500 9922 28552
rect 10229 28543 10287 28549
rect 10229 28509 10241 28543
rect 10275 28540 10287 28543
rect 10318 28540 10324 28552
rect 10275 28512 10324 28540
rect 10275 28509 10287 28512
rect 10229 28503 10287 28509
rect 10318 28500 10324 28512
rect 10376 28500 10382 28552
rect 10781 28543 10839 28549
rect 10781 28509 10793 28543
rect 10827 28509 10839 28543
rect 10781 28503 10839 28509
rect 8352 28444 9076 28472
rect 9140 28444 9444 28472
rect 8352 28432 8358 28444
rect 2041 28407 2099 28413
rect 2041 28373 2053 28407
rect 2087 28404 2099 28407
rect 2222 28404 2228 28416
rect 2087 28376 2228 28404
rect 2087 28373 2099 28376
rect 2041 28367 2099 28373
rect 2222 28364 2228 28376
rect 2280 28364 2286 28416
rect 2682 28404 2688 28416
rect 2643 28376 2688 28404
rect 2682 28364 2688 28376
rect 2740 28364 2746 28416
rect 3329 28407 3387 28413
rect 3329 28373 3341 28407
rect 3375 28404 3387 28407
rect 3878 28404 3884 28416
rect 3375 28376 3884 28404
rect 3375 28373 3387 28376
rect 3329 28367 3387 28373
rect 3878 28364 3884 28376
rect 3936 28364 3942 28416
rect 4062 28404 4068 28416
rect 4023 28376 4068 28404
rect 4062 28364 4068 28376
rect 4120 28364 4126 28416
rect 4614 28364 4620 28416
rect 4672 28404 4678 28416
rect 4709 28407 4767 28413
rect 4709 28404 4721 28407
rect 4672 28376 4721 28404
rect 4672 28364 4678 28376
rect 4709 28373 4721 28376
rect 4755 28373 4767 28407
rect 4709 28367 4767 28373
rect 5258 28364 5264 28416
rect 5316 28404 5322 28416
rect 5353 28407 5411 28413
rect 5353 28404 5365 28407
rect 5316 28376 5365 28404
rect 5316 28364 5322 28376
rect 5353 28373 5365 28376
rect 5399 28373 5411 28407
rect 5353 28367 5411 28373
rect 6086 28364 6092 28416
rect 6144 28404 6150 28416
rect 6181 28407 6239 28413
rect 6181 28404 6193 28407
rect 6144 28376 6193 28404
rect 6144 28364 6150 28376
rect 6181 28373 6193 28376
rect 6227 28373 6239 28407
rect 6181 28367 6239 28373
rect 8481 28407 8539 28413
rect 8481 28373 8493 28407
rect 8527 28404 8539 28407
rect 8754 28404 8760 28416
rect 8527 28376 8760 28404
rect 8527 28373 8539 28376
rect 8481 28367 8539 28373
rect 8754 28364 8760 28376
rect 8812 28364 8818 28416
rect 9048 28404 9076 28444
rect 9309 28407 9367 28413
rect 9309 28404 9321 28407
rect 9048 28376 9321 28404
rect 9309 28373 9321 28376
rect 9355 28373 9367 28407
rect 9416 28404 9444 28444
rect 9582 28432 9588 28484
rect 9640 28472 9646 28484
rect 10796 28472 10824 28503
rect 11514 28500 11520 28552
rect 11572 28540 11578 28552
rect 11609 28543 11667 28549
rect 11609 28540 11621 28543
rect 11572 28512 11621 28540
rect 11572 28500 11578 28512
rect 11609 28509 11621 28512
rect 11655 28509 11667 28543
rect 16206 28540 16212 28552
rect 16167 28512 16212 28540
rect 11609 28503 11667 28509
rect 16206 28500 16212 28512
rect 16264 28500 16270 28552
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 16758 28540 16764 28552
rect 16632 28512 16764 28540
rect 16632 28500 16638 28512
rect 16758 28500 16764 28512
rect 16816 28540 16822 28552
rect 16853 28543 16911 28549
rect 16853 28540 16865 28543
rect 16816 28512 16865 28540
rect 16816 28500 16822 28512
rect 16853 28509 16865 28512
rect 16899 28509 16911 28543
rect 16853 28503 16911 28509
rect 17402 28500 17408 28552
rect 17460 28540 17466 28552
rect 17497 28543 17555 28549
rect 17497 28540 17509 28543
rect 17460 28512 17509 28540
rect 17460 28500 17466 28512
rect 17497 28509 17509 28512
rect 17543 28540 17555 28543
rect 17586 28540 17592 28552
rect 17543 28512 17592 28540
rect 17543 28509 17555 28512
rect 17497 28503 17555 28509
rect 17586 28500 17592 28512
rect 17644 28500 17650 28552
rect 18693 28543 18751 28549
rect 18693 28509 18705 28543
rect 18739 28509 18751 28543
rect 18693 28503 18751 28509
rect 12342 28472 12348 28484
rect 9640 28444 10824 28472
rect 12303 28444 12348 28472
rect 9640 28432 9646 28444
rect 12342 28432 12348 28444
rect 12400 28432 12406 28484
rect 12437 28475 12495 28481
rect 12437 28441 12449 28475
rect 12483 28441 12495 28475
rect 13354 28472 13360 28484
rect 13315 28444 13360 28472
rect 12437 28435 12495 28441
rect 9766 28404 9772 28416
rect 9416 28376 9772 28404
rect 9309 28367 9367 28373
rect 9766 28364 9772 28376
rect 9824 28364 9830 28416
rect 10042 28404 10048 28416
rect 10003 28376 10048 28404
rect 10042 28364 10048 28376
rect 10100 28364 10106 28416
rect 10410 28364 10416 28416
rect 10468 28404 10474 28416
rect 10873 28407 10931 28413
rect 10873 28404 10885 28407
rect 10468 28376 10885 28404
rect 10468 28364 10474 28376
rect 10873 28373 10885 28376
rect 10919 28373 10931 28407
rect 10873 28367 10931 28373
rect 11701 28407 11759 28413
rect 11701 28373 11713 28407
rect 11747 28404 11759 28407
rect 12452 28404 12480 28435
rect 13354 28432 13360 28444
rect 13412 28432 13418 28484
rect 13722 28432 13728 28484
rect 13780 28472 13786 28484
rect 14369 28475 14427 28481
rect 14369 28472 14381 28475
rect 13780 28444 14381 28472
rect 13780 28432 13786 28444
rect 14369 28441 14381 28444
rect 14415 28441 14427 28475
rect 14369 28435 14427 28441
rect 14461 28475 14519 28481
rect 14461 28441 14473 28475
rect 14507 28472 14519 28475
rect 14918 28472 14924 28484
rect 14507 28444 14924 28472
rect 14507 28441 14519 28444
rect 14461 28435 14519 28441
rect 14918 28432 14924 28444
rect 14976 28432 14982 28484
rect 15378 28472 15384 28484
rect 15339 28444 15384 28472
rect 15378 28432 15384 28444
rect 15436 28432 15442 28484
rect 18708 28472 18736 28503
rect 19058 28500 19064 28552
rect 19116 28540 19122 28552
rect 19429 28543 19487 28549
rect 19429 28540 19441 28543
rect 19116 28512 19441 28540
rect 19116 28500 19122 28512
rect 19429 28509 19441 28512
rect 19475 28509 19487 28543
rect 20346 28540 20352 28552
rect 20307 28512 20352 28540
rect 19429 28503 19487 28509
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 20806 28540 20812 28552
rect 20767 28512 20812 28540
rect 20806 28500 20812 28512
rect 20864 28500 20870 28552
rect 21910 28540 21916 28552
rect 21871 28512 21916 28540
rect 21910 28500 21916 28512
rect 21968 28540 21974 28552
rect 23293 28543 23351 28549
rect 23293 28540 23305 28543
rect 21968 28512 23305 28540
rect 21968 28500 21974 28512
rect 23293 28509 23305 28512
rect 23339 28509 23351 28543
rect 23293 28503 23351 28509
rect 23842 28500 23848 28552
rect 23900 28540 23906 28552
rect 24765 28543 24823 28549
rect 24765 28540 24777 28543
rect 23900 28512 24777 28540
rect 23900 28500 23906 28512
rect 24765 28509 24777 28512
rect 24811 28509 24823 28543
rect 26789 28543 26847 28549
rect 26789 28540 26801 28543
rect 24765 28503 24823 28509
rect 26160 28512 26801 28540
rect 26160 28484 26188 28512
rect 26789 28509 26801 28512
rect 26835 28509 26847 28543
rect 27430 28540 27436 28552
rect 27391 28512 27436 28540
rect 26789 28503 26847 28509
rect 27430 28500 27436 28512
rect 27488 28500 27494 28552
rect 31941 28543 31999 28549
rect 31941 28509 31953 28543
rect 31987 28540 31999 28543
rect 36998 28540 37004 28552
rect 31987 28512 37004 28540
rect 31987 28509 31999 28512
rect 31941 28503 31999 28509
rect 36998 28500 37004 28512
rect 37056 28500 37062 28552
rect 15488 28444 18736 28472
rect 11747 28376 12480 28404
rect 11747 28373 11759 28376
rect 11701 28367 11759 28373
rect 12526 28364 12532 28416
rect 12584 28404 12590 28416
rect 15488 28404 15516 28444
rect 19150 28432 19156 28484
rect 19208 28472 19214 28484
rect 24946 28472 24952 28484
rect 19208 28444 24952 28472
rect 19208 28432 19214 28444
rect 24946 28432 24952 28444
rect 25004 28432 25010 28484
rect 25406 28432 25412 28484
rect 25464 28472 25470 28484
rect 25464 28444 25509 28472
rect 25464 28432 25470 28444
rect 26142 28432 26148 28484
rect 26200 28432 26206 28484
rect 12584 28376 15516 28404
rect 12584 28364 12590 28376
rect 15746 28364 15752 28416
rect 15804 28404 15810 28416
rect 16301 28407 16359 28413
rect 16301 28404 16313 28407
rect 15804 28376 16313 28404
rect 15804 28364 15810 28376
rect 16301 28373 16313 28376
rect 16347 28373 16359 28407
rect 16301 28367 16359 28373
rect 16945 28407 17003 28413
rect 16945 28373 16957 28407
rect 16991 28404 17003 28407
rect 19058 28404 19064 28416
rect 16991 28376 19064 28404
rect 16991 28373 17003 28376
rect 16945 28367 17003 28373
rect 19058 28364 19064 28376
rect 19116 28364 19122 28416
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 19521 28407 19579 28413
rect 19521 28404 19533 28407
rect 19392 28376 19533 28404
rect 19392 28364 19398 28376
rect 19521 28373 19533 28376
rect 19567 28373 19579 28407
rect 19521 28367 19579 28373
rect 20254 28364 20260 28416
rect 20312 28404 20318 28416
rect 20901 28407 20959 28413
rect 20901 28404 20913 28407
rect 20312 28376 20913 28404
rect 20312 28364 20318 28376
rect 20901 28373 20913 28376
rect 20947 28373 20959 28407
rect 20901 28367 20959 28373
rect 21542 28364 21548 28416
rect 21600 28404 21606 28416
rect 22005 28407 22063 28413
rect 22005 28404 22017 28407
rect 21600 28376 22017 28404
rect 21600 28364 21606 28376
rect 22005 28373 22017 28376
rect 22051 28373 22063 28407
rect 22005 28367 22063 28373
rect 25958 28364 25964 28416
rect 26016 28404 26022 28416
rect 27525 28407 27583 28413
rect 27525 28404 27537 28407
rect 26016 28376 27537 28404
rect 26016 28364 26022 28376
rect 27525 28373 27537 28376
rect 27571 28373 27583 28407
rect 32030 28404 32036 28416
rect 31991 28376 32036 28404
rect 27525 28367 27583 28373
rect 32030 28364 32036 28376
rect 32088 28364 32094 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3421 28203 3479 28209
rect 3421 28169 3433 28203
rect 3467 28200 3479 28203
rect 3467 28172 6592 28200
rect 3467 28169 3479 28172
rect 3421 28163 3479 28169
rect 3878 28092 3884 28144
rect 3936 28132 3942 28144
rect 5445 28135 5503 28141
rect 5445 28132 5457 28135
rect 3936 28104 5457 28132
rect 3936 28092 3942 28104
rect 5445 28101 5457 28104
rect 5491 28101 5503 28135
rect 5445 28095 5503 28101
rect 5810 28092 5816 28144
rect 5868 28132 5874 28144
rect 5997 28135 6055 28141
rect 5997 28132 6009 28135
rect 5868 28104 6009 28132
rect 5868 28092 5874 28104
rect 5997 28101 6009 28104
rect 6043 28132 6055 28135
rect 6454 28132 6460 28144
rect 6043 28104 6460 28132
rect 6043 28101 6055 28104
rect 5997 28095 6055 28101
rect 6454 28092 6460 28104
rect 6512 28092 6518 28144
rect 1578 28064 1584 28076
rect 1539 28036 1584 28064
rect 1578 28024 1584 28036
rect 1636 28024 1642 28076
rect 2685 28067 2743 28073
rect 2685 28033 2697 28067
rect 2731 28064 2743 28067
rect 2866 28064 2872 28076
rect 2731 28036 2872 28064
rect 2731 28033 2743 28036
rect 2685 28027 2743 28033
rect 2866 28024 2872 28036
rect 2924 28064 2930 28076
rect 3329 28067 3387 28073
rect 3329 28064 3341 28067
rect 2924 28036 3341 28064
rect 2924 28024 2930 28036
rect 3329 28033 3341 28036
rect 3375 28033 3387 28067
rect 3329 28027 3387 28033
rect 3418 28024 3424 28076
rect 3476 28064 3482 28076
rect 3973 28067 4031 28073
rect 3973 28064 3985 28067
rect 3476 28036 3985 28064
rect 3476 28024 3482 28036
rect 3973 28033 3985 28036
rect 4019 28033 4031 28067
rect 3973 28027 4031 28033
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28064 4675 28067
rect 4798 28064 4804 28076
rect 4663 28036 4804 28064
rect 4663 28033 4675 28036
rect 4617 28027 4675 28033
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 2777 27999 2835 28005
rect 2777 27965 2789 27999
rect 2823 27996 2835 27999
rect 5353 27999 5411 28005
rect 2823 27968 5304 27996
rect 2823 27965 2835 27968
rect 2777 27959 2835 27965
rect 1762 27928 1768 27940
rect 1723 27900 1768 27928
rect 1762 27888 1768 27900
rect 1820 27888 1826 27940
rect 3878 27888 3884 27940
rect 3936 27928 3942 27940
rect 4709 27931 4767 27937
rect 4709 27928 4721 27931
rect 3936 27900 4721 27928
rect 3936 27888 3942 27900
rect 4709 27897 4721 27900
rect 4755 27897 4767 27931
rect 5276 27928 5304 27968
rect 5353 27965 5365 27999
rect 5399 27996 5411 27999
rect 5718 27996 5724 28008
rect 5399 27968 5724 27996
rect 5399 27965 5411 27968
rect 5353 27959 5411 27965
rect 5718 27956 5724 27968
rect 5776 27956 5782 28008
rect 6564 27996 6592 28172
rect 6914 28160 6920 28212
rect 6972 28160 6978 28212
rect 9030 28200 9036 28212
rect 8036 28172 9036 28200
rect 6932 28132 6960 28160
rect 7101 28135 7159 28141
rect 7101 28132 7113 28135
rect 6932 28104 7113 28132
rect 7101 28101 7113 28104
rect 7147 28101 7159 28135
rect 7101 28095 7159 28101
rect 7374 28092 7380 28144
rect 7432 28132 7438 28144
rect 8036 28141 8064 28172
rect 9030 28160 9036 28172
rect 9088 28200 9094 28212
rect 10962 28200 10968 28212
rect 9088 28172 10968 28200
rect 9088 28160 9094 28172
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11977 28203 12035 28209
rect 11977 28169 11989 28203
rect 12023 28200 12035 28203
rect 17126 28200 17132 28212
rect 12023 28172 17132 28200
rect 12023 28169 12035 28172
rect 11977 28163 12035 28169
rect 17126 28160 17132 28172
rect 17184 28160 17190 28212
rect 19242 28160 19248 28212
rect 19300 28160 19306 28212
rect 23750 28160 23756 28212
rect 23808 28200 23814 28212
rect 24305 28203 24363 28209
rect 24305 28200 24317 28203
rect 23808 28172 24317 28200
rect 23808 28160 23814 28172
rect 24305 28169 24317 28172
rect 24351 28169 24363 28203
rect 24305 28163 24363 28169
rect 24949 28203 25007 28209
rect 24949 28169 24961 28203
rect 24995 28200 25007 28203
rect 25406 28200 25412 28212
rect 24995 28172 25412 28200
rect 24995 28169 25007 28172
rect 24949 28163 25007 28169
rect 25406 28160 25412 28172
rect 25464 28160 25470 28212
rect 25958 28200 25964 28212
rect 25608 28172 25964 28200
rect 8021 28135 8079 28141
rect 7432 28104 7880 28132
rect 7432 28092 7438 28104
rect 7852 28064 7880 28104
rect 8021 28101 8033 28135
rect 8067 28101 8079 28135
rect 9674 28132 9680 28144
rect 8021 28095 8079 28101
rect 8588 28104 9680 28132
rect 8478 28064 8484 28076
rect 7852 28036 8484 28064
rect 8478 28024 8484 28036
rect 8536 28024 8542 28076
rect 6380 27968 6592 27996
rect 7009 27999 7067 28005
rect 5534 27928 5540 27940
rect 5276 27900 5540 27928
rect 4709 27891 4767 27897
rect 5534 27888 5540 27900
rect 5592 27888 5598 27940
rect 4065 27863 4123 27869
rect 4065 27829 4077 27863
rect 4111 27860 4123 27863
rect 5902 27860 5908 27872
rect 4111 27832 5908 27860
rect 4111 27829 4123 27832
rect 4065 27823 4123 27829
rect 5902 27820 5908 27832
rect 5960 27820 5966 27872
rect 6380 27860 6408 27968
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 7098 27996 7104 28008
rect 7055 27968 7104 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 8588 27996 8616 28104
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 9766 28092 9772 28144
rect 9824 28132 9830 28144
rect 9824 28104 10180 28132
rect 9824 28092 9830 28104
rect 10152 28076 10180 28104
rect 11146 28092 11152 28144
rect 11204 28132 11210 28144
rect 13265 28135 13323 28141
rect 13265 28132 13277 28135
rect 11204 28104 13277 28132
rect 11204 28092 11210 28104
rect 13265 28101 13277 28104
rect 13311 28101 13323 28135
rect 13265 28095 13323 28101
rect 13357 28135 13415 28141
rect 13357 28101 13369 28135
rect 13403 28132 13415 28135
rect 13814 28132 13820 28144
rect 13403 28104 13820 28132
rect 13403 28101 13415 28104
rect 13357 28095 13415 28101
rect 13814 28092 13820 28104
rect 13872 28092 13878 28144
rect 18598 28132 18604 28144
rect 18559 28104 18604 28132
rect 18598 28092 18604 28104
rect 18656 28092 18662 28144
rect 18966 28092 18972 28144
rect 19024 28132 19030 28144
rect 19260 28132 19288 28160
rect 20070 28132 20076 28144
rect 19024 28104 20076 28132
rect 19024 28092 19030 28104
rect 20070 28092 20076 28104
rect 20128 28092 20134 28144
rect 20254 28092 20260 28144
rect 20312 28132 20318 28144
rect 20542 28135 20600 28141
rect 20542 28132 20554 28135
rect 20312 28104 20554 28132
rect 20312 28092 20318 28104
rect 20542 28101 20554 28104
rect 20588 28101 20600 28135
rect 22094 28132 22100 28144
rect 22055 28104 22100 28132
rect 20542 28095 20600 28101
rect 22094 28092 22100 28104
rect 22152 28092 22158 28144
rect 25608 28141 25636 28172
rect 25958 28160 25964 28172
rect 26016 28160 26022 28212
rect 22189 28135 22247 28141
rect 22189 28101 22201 28135
rect 22235 28132 22247 28135
rect 23661 28135 23719 28141
rect 23661 28132 23673 28135
rect 22235 28104 23673 28132
rect 22235 28101 22247 28104
rect 22189 28095 22247 28101
rect 23661 28101 23673 28104
rect 23707 28101 23719 28135
rect 23661 28095 23719 28101
rect 25593 28135 25651 28141
rect 25593 28101 25605 28135
rect 25639 28101 25651 28135
rect 25593 28095 25651 28101
rect 25685 28135 25743 28141
rect 25685 28101 25697 28135
rect 25731 28132 25743 28135
rect 27249 28135 27307 28141
rect 27249 28132 27261 28135
rect 25731 28104 27261 28132
rect 25731 28101 25743 28104
rect 25685 28095 25743 28101
rect 27249 28101 27261 28104
rect 27295 28101 27307 28135
rect 27249 28095 27307 28101
rect 8938 28024 8944 28076
rect 8996 28064 9002 28076
rect 9309 28070 9367 28073
rect 9232 28067 9367 28070
rect 9232 28064 9321 28067
rect 8996 28042 9321 28064
rect 8996 28036 9260 28042
rect 8996 28024 9002 28036
rect 9309 28033 9321 28042
rect 9355 28033 9367 28067
rect 9950 28064 9956 28076
rect 9911 28036 9956 28064
rect 9309 28027 9367 28033
rect 9950 28024 9956 28036
rect 10008 28024 10014 28076
rect 10134 28024 10140 28076
rect 10192 28064 10198 28076
rect 10597 28067 10655 28073
rect 10597 28064 10609 28067
rect 10192 28036 10609 28064
rect 10192 28024 10198 28036
rect 10597 28033 10609 28036
rect 10643 28033 10655 28067
rect 10597 28027 10655 28033
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12434 28064 12440 28076
rect 11931 28036 12440 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12434 28024 12440 28036
rect 12492 28024 12498 28076
rect 12529 28067 12587 28073
rect 12529 28033 12541 28067
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 7760 27968 8616 27996
rect 9401 27999 9459 28005
rect 7760 27940 7788 27968
rect 9401 27965 9413 27999
rect 9447 27996 9459 27999
rect 11422 27996 11428 28008
rect 9447 27984 9536 27996
rect 9646 27984 11428 27996
rect 9447 27968 11428 27984
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 9508 27956 9674 27968
rect 11422 27956 11428 27968
rect 11480 27956 11486 28008
rect 12544 27996 12572 28027
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 12676 28036 12721 28064
rect 12676 28024 12682 28036
rect 14182 28024 14188 28076
rect 14240 28064 14246 28076
rect 15197 28067 15255 28073
rect 15197 28064 15209 28067
rect 14240 28036 15209 28064
rect 14240 28024 14246 28036
rect 15197 28033 15209 28036
rect 15243 28033 15255 28067
rect 15197 28027 15255 28033
rect 15562 28024 15568 28076
rect 15620 28064 15626 28076
rect 16117 28067 16175 28073
rect 16117 28064 16129 28067
rect 15620 28036 16129 28064
rect 15620 28024 15626 28036
rect 16117 28033 16129 28036
rect 16163 28064 16175 28067
rect 16390 28064 16396 28076
rect 16163 28036 16396 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 16390 28024 16396 28036
rect 16448 28024 16454 28076
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28064 16911 28067
rect 17034 28064 17040 28076
rect 16899 28036 17040 28064
rect 16899 28033 16911 28036
rect 16853 28027 16911 28033
rect 17034 28024 17040 28036
rect 17092 28024 17098 28076
rect 17494 28064 17500 28076
rect 17455 28036 17500 28064
rect 17494 28024 17500 28036
rect 17552 28024 17558 28076
rect 23569 28067 23627 28073
rect 23569 28064 23581 28067
rect 22940 28036 23581 28064
rect 13630 27996 13636 28008
rect 12544 27968 13636 27996
rect 13630 27956 13636 27968
rect 13688 27956 13694 28008
rect 14093 27999 14151 28005
rect 14093 27965 14105 27999
rect 14139 27965 14151 27999
rect 14093 27959 14151 27965
rect 15289 27999 15347 28005
rect 15289 27965 15301 27999
rect 15335 27996 15347 27999
rect 16666 27996 16672 28008
rect 15335 27968 16672 27996
rect 15335 27965 15347 27968
rect 15289 27959 15347 27965
rect 7742 27888 7748 27940
rect 7800 27888 7806 27940
rect 8478 27888 8484 27940
rect 8536 27928 8542 27940
rect 10045 27931 10103 27937
rect 10045 27928 10057 27931
rect 8536 27900 10057 27928
rect 8536 27888 8542 27900
rect 10045 27897 10057 27900
rect 10091 27897 10103 27931
rect 13998 27928 14004 27940
rect 10045 27891 10103 27897
rect 10520 27900 14004 27928
rect 7098 27860 7104 27872
rect 6380 27832 7104 27860
rect 7098 27820 7104 27832
rect 7156 27820 7162 27872
rect 8386 27820 8392 27872
rect 8444 27860 8450 27872
rect 8573 27863 8631 27869
rect 8573 27860 8585 27863
rect 8444 27832 8585 27860
rect 8444 27820 8450 27832
rect 8573 27829 8585 27832
rect 8619 27829 8631 27863
rect 8573 27823 8631 27829
rect 8662 27820 8668 27872
rect 8720 27860 8726 27872
rect 10520 27860 10548 27900
rect 13998 27888 14004 27900
rect 14056 27888 14062 27940
rect 10686 27860 10692 27872
rect 8720 27832 10548 27860
rect 10647 27832 10692 27860
rect 8720 27820 8726 27832
rect 10686 27820 10692 27832
rect 10744 27820 10750 27872
rect 10962 27820 10968 27872
rect 11020 27860 11026 27872
rect 13078 27860 13084 27872
rect 11020 27832 13084 27860
rect 11020 27820 11026 27832
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 13170 27820 13176 27872
rect 13228 27860 13234 27872
rect 14108 27860 14136 27959
rect 16666 27956 16672 27968
rect 16724 27956 16730 28008
rect 17402 27956 17408 28008
rect 17460 27996 17466 28008
rect 18509 27999 18567 28005
rect 17460 27968 17724 27996
rect 17460 27956 17466 27968
rect 16114 27888 16120 27940
rect 16172 27928 16178 27940
rect 17589 27931 17647 27937
rect 17589 27928 17601 27931
rect 16172 27900 17601 27928
rect 16172 27888 16178 27900
rect 17589 27897 17601 27900
rect 17635 27897 17647 27931
rect 17696 27928 17724 27968
rect 18509 27965 18521 27999
rect 18555 27996 18567 27999
rect 19426 27996 19432 28008
rect 18555 27968 19432 27996
rect 18555 27965 18567 27968
rect 18509 27959 18567 27965
rect 19426 27956 19432 27968
rect 19484 27956 19490 28008
rect 19521 27999 19579 28005
rect 19521 27965 19533 27999
rect 19567 27965 19579 27999
rect 19521 27959 19579 27965
rect 20441 27999 20499 28005
rect 20441 27965 20453 27999
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 19536 27928 19564 27959
rect 17696 27900 19564 27928
rect 20464 27928 20492 27959
rect 20530 27956 20536 28008
rect 20588 27996 20594 28008
rect 20717 27999 20775 28005
rect 20717 27996 20729 27999
rect 20588 27968 20729 27996
rect 20588 27956 20594 27968
rect 20717 27965 20729 27968
rect 20763 27965 20775 27999
rect 20717 27959 20775 27965
rect 22462 27956 22468 28008
rect 22520 27996 22526 28008
rect 22940 27996 22968 28036
rect 23569 28033 23581 28036
rect 23615 28033 23627 28067
rect 24210 28064 24216 28076
rect 24171 28036 24216 28064
rect 23569 28027 23627 28033
rect 24210 28024 24216 28036
rect 24268 28024 24274 28076
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28064 24915 28067
rect 25130 28064 25136 28076
rect 24903 28036 25136 28064
rect 24903 28033 24915 28036
rect 24857 28027 24915 28033
rect 25130 28024 25136 28036
rect 25188 28024 25194 28076
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28064 27215 28067
rect 27798 28064 27804 28076
rect 27203 28036 27804 28064
rect 27203 28033 27215 28036
rect 27157 28027 27215 28033
rect 27798 28024 27804 28036
rect 27856 28024 27862 28076
rect 22520 27968 22968 27996
rect 23109 27999 23167 28005
rect 22520 27956 22526 27968
rect 23109 27965 23121 27999
rect 23155 27996 23167 27999
rect 24762 27996 24768 28008
rect 23155 27968 24768 27996
rect 23155 27965 23167 27968
rect 23109 27959 23167 27965
rect 24762 27956 24768 27968
rect 24820 27956 24826 28008
rect 24946 27956 24952 28008
rect 25004 27996 25010 28008
rect 26605 27999 26663 28005
rect 26605 27996 26617 27999
rect 25004 27968 26617 27996
rect 25004 27956 25010 27968
rect 26605 27965 26617 27968
rect 26651 27996 26663 27999
rect 27430 27996 27436 28008
rect 26651 27968 27436 27996
rect 26651 27965 26663 27968
rect 26605 27959 26663 27965
rect 27430 27956 27436 27968
rect 27488 27956 27494 28008
rect 30742 27928 30748 27940
rect 20464 27900 30748 27928
rect 17589 27891 17647 27897
rect 30742 27888 30748 27900
rect 30800 27888 30806 27940
rect 31726 27900 35894 27928
rect 13228 27832 14136 27860
rect 16209 27863 16267 27869
rect 13228 27820 13234 27832
rect 16209 27829 16221 27863
rect 16255 27860 16267 27863
rect 16298 27860 16304 27872
rect 16255 27832 16304 27860
rect 16255 27829 16267 27832
rect 16209 27823 16267 27829
rect 16298 27820 16304 27832
rect 16356 27820 16362 27872
rect 16942 27860 16948 27872
rect 16903 27832 16948 27860
rect 16942 27820 16948 27832
rect 17000 27820 17006 27872
rect 17494 27820 17500 27872
rect 17552 27860 17558 27872
rect 31726 27860 31754 27900
rect 17552 27832 31754 27860
rect 35866 27860 35894 27900
rect 37642 27860 37648 27872
rect 35866 27832 37648 27860
rect 17552 27820 17558 27832
rect 37642 27820 37648 27832
rect 37700 27820 37706 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 4798 27616 4804 27668
rect 4856 27656 4862 27668
rect 9766 27656 9772 27668
rect 4856 27628 9772 27656
rect 4856 27616 4862 27628
rect 9766 27616 9772 27628
rect 9824 27616 9830 27668
rect 9858 27616 9864 27668
rect 9916 27656 9922 27668
rect 9916 27628 12940 27656
rect 9916 27616 9922 27628
rect 10042 27588 10048 27600
rect 1596 27560 10048 27588
rect 1596 27461 1624 27560
rect 10042 27548 10048 27560
rect 10100 27548 10106 27600
rect 10318 27548 10324 27600
rect 10376 27588 10382 27600
rect 10962 27588 10968 27600
rect 10376 27560 10968 27588
rect 10376 27548 10382 27560
rect 10962 27548 10968 27560
rect 11020 27548 11026 27600
rect 5994 27520 6000 27532
rect 4264 27492 6000 27520
rect 1581 27455 1639 27461
rect 1581 27421 1593 27455
rect 1627 27421 1639 27455
rect 1581 27415 1639 27421
rect 2593 27455 2651 27461
rect 2593 27421 2605 27455
rect 2639 27452 2651 27455
rect 3234 27452 3240 27464
rect 2639 27424 3240 27452
rect 2639 27421 2651 27424
rect 2593 27415 2651 27421
rect 3234 27412 3240 27424
rect 3292 27412 3298 27464
rect 4264 27461 4292 27492
rect 5994 27480 6000 27492
rect 6052 27480 6058 27532
rect 6822 27480 6828 27532
rect 6880 27520 6886 27532
rect 8202 27520 8208 27532
rect 6880 27492 8208 27520
rect 6880 27480 6886 27492
rect 8202 27480 8208 27492
rect 8260 27480 8266 27532
rect 8481 27523 8539 27529
rect 8481 27489 8493 27523
rect 8527 27520 8539 27523
rect 9398 27520 9404 27532
rect 8527 27492 9404 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 9398 27480 9404 27492
rect 9456 27480 9462 27532
rect 9582 27520 9588 27532
rect 9543 27492 9588 27520
rect 9582 27480 9588 27492
rect 9640 27480 9646 27532
rect 10781 27523 10839 27529
rect 10781 27489 10793 27523
rect 10827 27520 10839 27523
rect 11054 27520 11060 27532
rect 10827 27492 11060 27520
rect 10827 27489 10839 27492
rect 10781 27483 10839 27489
rect 11054 27480 11060 27492
rect 11112 27480 11118 27532
rect 12345 27523 12403 27529
rect 12345 27489 12357 27523
rect 12391 27520 12403 27523
rect 12710 27520 12716 27532
rect 12391 27492 12716 27520
rect 12391 27489 12403 27492
rect 12345 27483 12403 27489
rect 12710 27480 12716 27492
rect 12768 27480 12774 27532
rect 4249 27455 4307 27461
rect 4249 27421 4261 27455
rect 4295 27421 4307 27455
rect 4249 27415 4307 27421
rect 4798 27412 4804 27464
rect 4856 27452 4862 27464
rect 4893 27455 4951 27461
rect 4893 27452 4905 27455
rect 4856 27424 4905 27452
rect 4856 27412 4862 27424
rect 4893 27421 4905 27424
rect 4939 27421 4951 27455
rect 4893 27415 4951 27421
rect 4982 27412 4988 27464
rect 5040 27412 5046 27464
rect 6564 27424 6868 27452
rect 2866 27344 2872 27396
rect 2924 27384 2930 27396
rect 5000 27384 5028 27412
rect 5626 27384 5632 27396
rect 2924 27356 5028 27384
rect 5587 27356 5632 27384
rect 2924 27344 2930 27356
rect 5626 27344 5632 27356
rect 5684 27344 5690 27396
rect 5721 27387 5779 27393
rect 5721 27353 5733 27387
rect 5767 27353 5779 27387
rect 5721 27347 5779 27353
rect 1762 27316 1768 27328
rect 1723 27288 1768 27316
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 2406 27276 2412 27328
rect 2464 27316 2470 27328
rect 2685 27319 2743 27325
rect 2685 27316 2697 27319
rect 2464 27288 2697 27316
rect 2464 27276 2470 27288
rect 2685 27285 2697 27288
rect 2731 27285 2743 27319
rect 3326 27316 3332 27328
rect 3287 27288 3332 27316
rect 2685 27279 2743 27285
rect 3326 27276 3332 27288
rect 3384 27276 3390 27328
rect 4341 27319 4399 27325
rect 4341 27285 4353 27319
rect 4387 27316 4399 27319
rect 4798 27316 4804 27328
rect 4387 27288 4804 27316
rect 4387 27285 4399 27288
rect 4341 27279 4399 27285
rect 4798 27276 4804 27288
rect 4856 27276 4862 27328
rect 4985 27319 5043 27325
rect 4985 27285 4997 27319
rect 5031 27316 5043 27319
rect 5166 27316 5172 27328
rect 5031 27288 5172 27316
rect 5031 27285 5043 27288
rect 4985 27279 5043 27285
rect 5166 27276 5172 27288
rect 5224 27276 5230 27328
rect 5442 27276 5448 27328
rect 5500 27316 5506 27328
rect 5736 27316 5764 27347
rect 5810 27344 5816 27396
rect 5868 27384 5874 27396
rect 6564 27384 6592 27424
rect 5868 27356 6592 27384
rect 6641 27387 6699 27393
rect 5868 27344 5874 27356
rect 6641 27353 6653 27387
rect 6687 27353 6699 27387
rect 6840 27384 6868 27424
rect 6914 27412 6920 27464
rect 6972 27452 6978 27464
rect 7469 27455 7527 27461
rect 7469 27452 7481 27455
rect 6972 27424 7481 27452
rect 6972 27412 6978 27424
rect 7469 27421 7481 27424
rect 7515 27421 7527 27455
rect 7469 27415 7527 27421
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27452 8447 27455
rect 8754 27452 8760 27464
rect 8435 27424 8760 27452
rect 8435 27421 8447 27424
rect 8389 27415 8447 27421
rect 8754 27412 8760 27424
rect 8812 27412 8818 27464
rect 11882 27412 11888 27464
rect 11940 27452 11946 27464
rect 12912 27461 12940 27628
rect 15102 27616 15108 27668
rect 15160 27656 15166 27668
rect 15160 27628 16344 27656
rect 15160 27616 15166 27628
rect 13078 27548 13084 27600
rect 13136 27588 13142 27600
rect 16206 27588 16212 27600
rect 13136 27560 16212 27588
rect 13136 27548 13142 27560
rect 16206 27548 16212 27560
rect 16264 27548 16270 27600
rect 16316 27588 16344 27628
rect 16390 27616 16396 27668
rect 16448 27656 16454 27668
rect 25130 27656 25136 27668
rect 16448 27628 25136 27656
rect 16448 27616 16454 27628
rect 25130 27616 25136 27628
rect 25188 27616 25194 27668
rect 16574 27588 16580 27600
rect 16316 27560 16580 27588
rect 16574 27548 16580 27560
rect 16632 27548 16638 27600
rect 20714 27588 20720 27600
rect 20675 27560 20720 27588
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 21450 27548 21456 27600
rect 21508 27588 21514 27600
rect 21910 27588 21916 27600
rect 21508 27560 21916 27588
rect 21508 27548 21514 27560
rect 21910 27548 21916 27560
rect 21968 27588 21974 27600
rect 21968 27560 22094 27588
rect 21968 27548 21974 27560
rect 12989 27523 13047 27529
rect 12989 27489 13001 27523
rect 13035 27520 13047 27523
rect 13998 27520 14004 27532
rect 13035 27492 14004 27520
rect 13035 27489 13047 27492
rect 12989 27483 13047 27489
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 20165 27523 20223 27529
rect 14752 27492 16988 27520
rect 12253 27455 12311 27461
rect 12253 27452 12265 27455
rect 11940 27424 12265 27452
rect 11940 27412 11946 27424
rect 12253 27421 12265 27424
rect 12299 27421 12311 27455
rect 12253 27415 12311 27421
rect 12897 27455 12955 27461
rect 12897 27421 12909 27455
rect 12943 27421 12955 27455
rect 13541 27455 13599 27461
rect 13541 27452 13553 27455
rect 12897 27415 12955 27421
rect 13004 27424 13553 27452
rect 13004 27396 13032 27424
rect 13541 27421 13553 27424
rect 13587 27421 13599 27455
rect 14752 27452 14780 27492
rect 13541 27415 13599 27421
rect 14200 27424 14780 27452
rect 7006 27384 7012 27396
rect 6840 27356 7012 27384
rect 6641 27347 6699 27353
rect 5500 27288 5764 27316
rect 6656 27316 6684 27347
rect 7006 27344 7012 27356
rect 7064 27344 7070 27396
rect 7561 27387 7619 27393
rect 7561 27353 7573 27387
rect 7607 27384 7619 27387
rect 9214 27384 9220 27396
rect 7607 27356 9076 27384
rect 9175 27356 9220 27384
rect 7607 27353 7619 27356
rect 7561 27347 7619 27353
rect 8386 27316 8392 27328
rect 6656 27288 8392 27316
rect 5500 27276 5506 27288
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 9048 27316 9076 27356
rect 9214 27344 9220 27356
rect 9272 27344 9278 27396
rect 9309 27387 9367 27393
rect 9309 27353 9321 27387
rect 9355 27384 9367 27387
rect 9674 27384 9680 27396
rect 9355 27356 9680 27384
rect 9355 27353 9367 27356
rect 9309 27347 9367 27353
rect 9674 27344 9680 27356
rect 9732 27344 9738 27396
rect 10873 27387 10931 27393
rect 10873 27353 10885 27387
rect 10919 27353 10931 27387
rect 10873 27347 10931 27353
rect 10888 27316 10916 27347
rect 10962 27344 10968 27396
rect 11020 27384 11026 27396
rect 11793 27387 11851 27393
rect 11793 27384 11805 27387
rect 11020 27356 11805 27384
rect 11020 27344 11026 27356
rect 11793 27353 11805 27356
rect 11839 27384 11851 27387
rect 12526 27384 12532 27396
rect 11839 27356 12532 27384
rect 11839 27353 11851 27356
rect 11793 27347 11851 27353
rect 12526 27344 12532 27356
rect 12584 27344 12590 27396
rect 12986 27344 12992 27396
rect 13044 27344 13050 27396
rect 14200 27384 14228 27424
rect 13096 27356 14228 27384
rect 9048 27288 10916 27316
rect 11054 27276 11060 27328
rect 11112 27316 11118 27328
rect 13096 27316 13124 27356
rect 14274 27344 14280 27396
rect 14332 27384 14338 27396
rect 14642 27384 14648 27396
rect 14332 27356 14648 27384
rect 14332 27344 14338 27356
rect 14642 27344 14648 27356
rect 14700 27384 14706 27396
rect 14921 27387 14979 27393
rect 14921 27384 14933 27387
rect 14700 27356 14933 27384
rect 14700 27344 14706 27356
rect 14921 27353 14933 27356
rect 14967 27353 14979 27387
rect 14921 27347 14979 27353
rect 15013 27387 15071 27393
rect 15013 27353 15025 27387
rect 15059 27384 15071 27387
rect 15194 27384 15200 27396
rect 15059 27356 15200 27384
rect 15059 27353 15071 27356
rect 15013 27347 15071 27353
rect 11112 27288 13124 27316
rect 13633 27319 13691 27325
rect 11112 27276 11118 27288
rect 13633 27285 13645 27319
rect 13679 27316 13691 27319
rect 14090 27316 14096 27328
rect 13679 27288 14096 27316
rect 13679 27285 13691 27288
rect 13633 27279 13691 27285
rect 14090 27276 14096 27288
rect 14148 27276 14154 27328
rect 14936 27316 14964 27347
rect 15194 27344 15200 27356
rect 15252 27344 15258 27396
rect 15286 27344 15292 27396
rect 15344 27384 15350 27396
rect 15565 27387 15623 27393
rect 15565 27384 15577 27387
rect 15344 27356 15577 27384
rect 15344 27344 15350 27356
rect 15565 27353 15577 27356
rect 15611 27353 15623 27387
rect 16114 27384 16120 27396
rect 16075 27356 16120 27384
rect 15565 27347 15623 27353
rect 16114 27344 16120 27356
rect 16172 27344 16178 27396
rect 16206 27344 16212 27396
rect 16264 27384 16270 27396
rect 16960 27384 16988 27492
rect 20165 27489 20177 27523
rect 20211 27520 20223 27523
rect 20806 27520 20812 27532
rect 20211 27492 20812 27520
rect 20211 27489 20223 27492
rect 20165 27483 20223 27489
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 21361 27523 21419 27529
rect 21361 27489 21373 27523
rect 21407 27520 21419 27523
rect 21542 27520 21548 27532
rect 21407 27492 21548 27520
rect 21407 27489 21419 27492
rect 21361 27483 21419 27489
rect 21542 27480 21548 27492
rect 21600 27480 21606 27532
rect 22066 27520 22094 27560
rect 24762 27548 24768 27600
rect 24820 27588 24826 27600
rect 24820 27560 26648 27588
rect 24820 27548 24826 27560
rect 22557 27523 22615 27529
rect 22557 27520 22569 27523
rect 22066 27492 22569 27520
rect 22557 27489 22569 27492
rect 22603 27489 22615 27523
rect 22557 27483 22615 27489
rect 23569 27523 23627 27529
rect 23569 27489 23581 27523
rect 23615 27520 23627 27523
rect 24854 27520 24860 27532
rect 23615 27492 24860 27520
rect 23615 27489 23627 27492
rect 23569 27483 23627 27489
rect 24854 27480 24860 27492
rect 24912 27520 24918 27532
rect 25498 27520 25504 27532
rect 24912 27492 25504 27520
rect 24912 27480 24918 27492
rect 25498 27480 25504 27492
rect 25556 27480 25562 27532
rect 25685 27523 25743 27529
rect 25685 27489 25697 27523
rect 25731 27520 25743 27523
rect 26510 27520 26516 27532
rect 25731 27492 26516 27520
rect 25731 27489 25743 27492
rect 25685 27483 25743 27489
rect 26510 27480 26516 27492
rect 26568 27480 26574 27532
rect 26620 27529 26648 27560
rect 26605 27523 26663 27529
rect 26605 27489 26617 27523
rect 26651 27489 26663 27523
rect 27617 27523 27675 27529
rect 27617 27520 27629 27523
rect 26605 27483 26663 27489
rect 26804 27492 27629 27520
rect 17034 27412 17040 27464
rect 17092 27452 17098 27464
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 17092 27424 17601 27452
rect 17092 27412 17098 27424
rect 17589 27421 17601 27424
rect 17635 27452 17647 27455
rect 17862 27452 17868 27464
rect 17635 27424 17868 27452
rect 17635 27421 17647 27424
rect 17589 27415 17647 27421
rect 17862 27412 17868 27424
rect 17920 27412 17926 27464
rect 18506 27412 18512 27464
rect 18564 27452 18570 27464
rect 18693 27455 18751 27461
rect 18693 27452 18705 27455
rect 18564 27424 18705 27452
rect 18564 27412 18570 27424
rect 18693 27421 18705 27424
rect 18739 27452 18751 27455
rect 19150 27452 19156 27464
rect 18739 27424 19156 27452
rect 18739 27421 18751 27424
rect 18693 27415 18751 27421
rect 19150 27412 19156 27424
rect 19208 27412 19214 27464
rect 19426 27452 19432 27464
rect 19387 27424 19432 27452
rect 19426 27412 19432 27424
rect 19484 27412 19490 27464
rect 17129 27387 17187 27393
rect 17129 27384 17141 27387
rect 16264 27356 16309 27384
rect 16960 27356 17141 27384
rect 16264 27344 16270 27356
rect 17129 27353 17141 27356
rect 17175 27384 17187 27387
rect 17402 27384 17408 27396
rect 17175 27356 17408 27384
rect 17175 27353 17187 27356
rect 17129 27347 17187 27353
rect 17402 27344 17408 27356
rect 17460 27344 17466 27396
rect 18046 27384 18052 27396
rect 17512 27356 18052 27384
rect 17512 27316 17540 27356
rect 18046 27344 18052 27356
rect 18104 27344 18110 27396
rect 18785 27387 18843 27393
rect 18785 27353 18797 27387
rect 18831 27384 18843 27387
rect 20257 27387 20315 27393
rect 18831 27356 20116 27384
rect 18831 27353 18843 27356
rect 18785 27347 18843 27353
rect 17678 27316 17684 27328
rect 14936 27288 17540 27316
rect 17639 27288 17684 27316
rect 17678 27276 17684 27288
rect 17736 27276 17742 27328
rect 19521 27319 19579 27325
rect 19521 27285 19533 27319
rect 19567 27316 19579 27319
rect 19978 27316 19984 27328
rect 19567 27288 19984 27316
rect 19567 27285 19579 27288
rect 19521 27279 19579 27285
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 20088 27316 20116 27356
rect 20257 27353 20269 27387
rect 20303 27353 20315 27387
rect 20257 27347 20315 27353
rect 20272 27316 20300 27347
rect 21450 27344 21456 27396
rect 21508 27384 21514 27396
rect 22005 27387 22063 27393
rect 21508 27356 21553 27384
rect 21508 27344 21514 27356
rect 22005 27353 22017 27387
rect 22051 27384 22063 27387
rect 22051 27356 22085 27384
rect 22051 27353 22063 27356
rect 22005 27347 22063 27353
rect 20088 27288 20300 27316
rect 21358 27276 21364 27328
rect 21416 27316 21422 27328
rect 22020 27316 22048 27347
rect 22370 27344 22376 27396
rect 22428 27384 22434 27396
rect 22649 27387 22707 27393
rect 22649 27384 22661 27387
rect 22428 27356 22661 27384
rect 22428 27344 22434 27356
rect 22649 27353 22661 27356
rect 22695 27353 22707 27387
rect 22649 27347 22707 27353
rect 25777 27387 25835 27393
rect 25777 27353 25789 27387
rect 25823 27384 25835 27387
rect 25866 27384 25872 27396
rect 25823 27356 25872 27384
rect 25823 27353 25835 27356
rect 25777 27347 25835 27353
rect 25866 27344 25872 27356
rect 25924 27344 25930 27396
rect 26050 27316 26056 27328
rect 21416 27288 26056 27316
rect 21416 27276 21422 27288
rect 26050 27276 26056 27288
rect 26108 27316 26114 27328
rect 26804 27316 26832 27492
rect 27617 27489 27629 27492
rect 27663 27489 27675 27523
rect 27617 27483 27675 27489
rect 37366 27480 37372 27532
rect 37424 27520 37430 27532
rect 37737 27523 37795 27529
rect 37737 27520 37749 27523
rect 37424 27492 37749 27520
rect 37424 27480 37430 27492
rect 37737 27489 37749 27492
rect 37783 27489 37795 27523
rect 37737 27483 37795 27489
rect 27890 27412 27896 27464
rect 27948 27452 27954 27464
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 27948 27424 28365 27452
rect 27948 27412 27954 27424
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 37458 27452 37464 27464
rect 37419 27424 37464 27452
rect 28353 27415 28411 27421
rect 37458 27412 37464 27424
rect 37516 27412 37522 27464
rect 27246 27384 27252 27396
rect 27207 27356 27252 27384
rect 27246 27344 27252 27356
rect 27304 27344 27310 27396
rect 27341 27387 27399 27393
rect 27341 27353 27353 27387
rect 27387 27353 27399 27387
rect 27341 27347 27399 27353
rect 26108 27288 26832 27316
rect 27356 27316 27384 27347
rect 28445 27319 28503 27325
rect 28445 27316 28457 27319
rect 27356 27288 28457 27316
rect 26108 27276 26114 27288
rect 28445 27285 28457 27288
rect 28491 27285 28503 27319
rect 28445 27279 28503 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 4890 27072 4896 27124
rect 4948 27112 4954 27124
rect 9214 27112 9220 27124
rect 4948 27084 8892 27112
rect 9127 27084 9220 27112
rect 4948 27072 4954 27084
rect 934 27004 940 27056
rect 992 27044 998 27056
rect 992 27016 6868 27044
rect 992 27004 998 27016
rect 1949 26979 2007 26985
rect 1949 26945 1961 26979
rect 1995 26976 2007 26979
rect 2130 26976 2136 26988
rect 1995 26948 2136 26976
rect 1995 26945 2007 26948
rect 1949 26939 2007 26945
rect 2130 26936 2136 26948
rect 2188 26936 2194 26988
rect 2590 26976 2596 26988
rect 2551 26948 2596 26976
rect 2590 26936 2596 26948
rect 2648 26936 2654 26988
rect 3234 26976 3240 26988
rect 3195 26948 3240 26976
rect 3234 26936 3240 26948
rect 3292 26936 3298 26988
rect 3881 26979 3939 26985
rect 3881 26945 3893 26979
rect 3927 26945 3939 26979
rect 3881 26939 3939 26945
rect 1578 26868 1584 26920
rect 1636 26908 1642 26920
rect 3896 26908 3924 26939
rect 4062 26936 4068 26988
rect 4120 26976 4126 26988
rect 4525 26979 4583 26985
rect 4525 26976 4537 26979
rect 4120 26948 4537 26976
rect 4120 26936 4126 26948
rect 4525 26945 4537 26948
rect 4571 26945 4583 26979
rect 4525 26939 4583 26945
rect 5169 26979 5227 26985
rect 5169 26945 5181 26979
rect 5215 26976 5227 26979
rect 5718 26976 5724 26988
rect 5215 26948 5724 26976
rect 5215 26945 5227 26948
rect 5169 26939 5227 26945
rect 5718 26936 5724 26948
rect 5776 26936 5782 26988
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 6641 26979 6699 26985
rect 6641 26945 6653 26979
rect 6687 26976 6699 26979
rect 6730 26976 6736 26988
rect 6687 26948 6736 26976
rect 6687 26945 6699 26948
rect 6641 26939 6699 26945
rect 1636 26880 3924 26908
rect 3973 26911 4031 26917
rect 1636 26868 1642 26880
rect 3973 26877 3985 26911
rect 4019 26908 4031 26911
rect 5442 26908 5448 26920
rect 4019 26880 5448 26908
rect 4019 26877 4031 26880
rect 3973 26871 4031 26877
rect 5442 26868 5448 26880
rect 5500 26868 5506 26920
rect 5828 26908 5856 26939
rect 6730 26936 6736 26948
rect 6788 26936 6794 26988
rect 6840 26976 6868 27016
rect 7190 27004 7196 27056
rect 7248 27044 7254 27056
rect 8864 27053 8892 27084
rect 9214 27072 9220 27084
rect 9272 27112 9278 27124
rect 11238 27112 11244 27124
rect 9272 27084 11244 27112
rect 9272 27072 9278 27084
rect 11238 27072 11244 27084
rect 11296 27072 11302 27124
rect 12710 27072 12716 27124
rect 12768 27112 12774 27124
rect 14274 27112 14280 27124
rect 12768 27084 14280 27112
rect 12768 27072 12774 27084
rect 14274 27072 14280 27084
rect 14332 27072 14338 27124
rect 14642 27072 14648 27124
rect 14700 27112 14706 27124
rect 21266 27112 21272 27124
rect 14700 27084 21272 27112
rect 14700 27072 14706 27084
rect 21266 27072 21272 27084
rect 21324 27072 21330 27124
rect 21361 27115 21419 27121
rect 21361 27081 21373 27115
rect 21407 27112 21419 27115
rect 21450 27112 21456 27124
rect 21407 27084 21456 27112
rect 21407 27081 21419 27084
rect 21361 27075 21419 27081
rect 21450 27072 21456 27084
rect 21508 27072 21514 27124
rect 25866 27112 25872 27124
rect 25827 27084 25872 27112
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 27246 27072 27252 27124
rect 27304 27112 27310 27124
rect 30742 27112 30748 27124
rect 27304 27084 28764 27112
rect 30703 27084 30748 27112
rect 27304 27072 27310 27084
rect 8297 27047 8355 27053
rect 8297 27044 8309 27047
rect 7248 27016 8309 27044
rect 7248 27004 7254 27016
rect 8297 27013 8309 27016
rect 8343 27013 8355 27047
rect 8297 27007 8355 27013
rect 8849 27047 8907 27053
rect 8849 27013 8861 27047
rect 8895 27013 8907 27047
rect 8849 27007 8907 27013
rect 7285 26979 7343 26985
rect 7285 26976 7297 26979
rect 6840 26948 7297 26976
rect 7285 26945 7297 26948
rect 7331 26976 7343 26979
rect 7374 26976 7380 26988
rect 7331 26948 7380 26976
rect 7331 26945 7343 26948
rect 7285 26939 7343 26945
rect 7374 26936 7380 26948
rect 7432 26936 7438 26988
rect 8202 26908 8208 26920
rect 5828 26880 6644 26908
rect 6638 26856 6644 26880
rect 6696 26856 6702 26908
rect 8163 26880 8208 26908
rect 8202 26868 8208 26880
rect 8260 26868 8266 26920
rect 3329 26843 3387 26849
rect 3329 26809 3341 26843
rect 3375 26840 3387 26843
rect 4982 26840 4988 26852
rect 3375 26812 4988 26840
rect 3375 26809 3387 26812
rect 3329 26803 3387 26809
rect 4982 26800 4988 26812
rect 5040 26800 5046 26852
rect 5261 26843 5319 26849
rect 5261 26809 5273 26843
rect 5307 26840 5319 26843
rect 6178 26840 6184 26852
rect 5307 26812 6184 26840
rect 5307 26809 5319 26812
rect 5261 26803 5319 26809
rect 6178 26800 6184 26812
rect 6236 26800 6242 26852
rect 6733 26843 6791 26849
rect 6733 26809 6745 26843
rect 6779 26840 6791 26843
rect 8864 26840 8892 27007
rect 9232 26908 9260 27072
rect 9490 27044 9496 27056
rect 9451 27016 9496 27044
rect 9490 27004 9496 27016
rect 9548 27004 9554 27056
rect 10870 27004 10876 27056
rect 10928 27044 10934 27056
rect 11885 27047 11943 27053
rect 11885 27044 11897 27047
rect 10928 27016 11897 27044
rect 10928 27004 10934 27016
rect 11885 27013 11897 27016
rect 11931 27013 11943 27047
rect 11885 27007 11943 27013
rect 12434 27004 12440 27056
rect 12492 27044 12498 27056
rect 12492 27016 12664 27044
rect 12492 27004 12498 27016
rect 10962 26976 10968 26988
rect 10923 26948 10968 26976
rect 10962 26936 10968 26948
rect 11020 26936 11026 26988
rect 12636 26976 12664 27016
rect 13170 27004 13176 27056
rect 13228 27044 13234 27056
rect 13228 27016 14872 27044
rect 13228 27004 13234 27016
rect 13354 26976 13360 26988
rect 12636 26948 13360 26976
rect 13354 26936 13360 26948
rect 13412 26936 13418 26988
rect 13538 26976 13544 26988
rect 13499 26948 13544 26976
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 14182 26976 14188 26988
rect 14143 26948 14188 26976
rect 14182 26936 14188 26948
rect 14240 26936 14246 26988
rect 14844 26985 14872 27016
rect 18506 27004 18512 27056
rect 18564 27044 18570 27056
rect 19058 27044 19064 27056
rect 18564 27016 19064 27044
rect 18564 27004 18570 27016
rect 19058 27004 19064 27016
rect 19116 27004 19122 27056
rect 19153 27047 19211 27053
rect 19153 27013 19165 27047
rect 19199 27044 19211 27047
rect 19334 27044 19340 27056
rect 19199 27016 19340 27044
rect 19199 27013 19211 27016
rect 19153 27007 19211 27013
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 19426 27004 19432 27056
rect 19484 27044 19490 27056
rect 22462 27044 22468 27056
rect 19484 27016 22468 27044
rect 19484 27004 19490 27016
rect 22462 27004 22468 27016
rect 22520 27004 22526 27056
rect 22738 27044 22744 27056
rect 22699 27016 22744 27044
rect 22738 27004 22744 27016
rect 22796 27004 22802 27056
rect 23290 27004 23296 27056
rect 23348 27044 23354 27056
rect 27709 27047 27767 27053
rect 27709 27044 27721 27047
rect 23348 27016 27721 27044
rect 23348 27004 23354 27016
rect 27709 27013 27721 27016
rect 27755 27013 27767 27047
rect 27709 27007 27767 27013
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 15654 26976 15660 26988
rect 15615 26948 15660 26976
rect 14829 26939 14887 26945
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 16022 26936 16028 26988
rect 16080 26976 16086 26988
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16080 26948 16865 26976
rect 16080 26936 16086 26948
rect 16853 26945 16865 26948
rect 16899 26976 16911 26979
rect 17310 26976 17316 26988
rect 16899 26948 17316 26976
rect 16899 26945 16911 26948
rect 16853 26939 16911 26945
rect 17310 26936 17316 26948
rect 17368 26936 17374 26988
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26976 17555 26979
rect 17586 26976 17592 26988
rect 17543 26948 17592 26976
rect 17543 26945 17555 26948
rect 17497 26939 17555 26945
rect 17586 26936 17592 26948
rect 17644 26936 17650 26988
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26976 18199 26979
rect 18690 26976 18696 26988
rect 18187 26948 18696 26976
rect 18187 26945 18199 26948
rect 18141 26939 18199 26945
rect 18690 26936 18696 26948
rect 18748 26936 18754 26988
rect 20162 26976 20168 26988
rect 19904 26948 20168 26976
rect 9401 26911 9459 26917
rect 9401 26908 9413 26911
rect 9232 26880 9413 26908
rect 9401 26877 9413 26880
rect 9447 26877 9459 26911
rect 9401 26871 9459 26877
rect 9677 26911 9735 26917
rect 9677 26877 9689 26911
rect 9723 26877 9735 26911
rect 9677 26871 9735 26877
rect 11793 26911 11851 26917
rect 11793 26877 11805 26911
rect 11839 26908 11851 26911
rect 12434 26908 12440 26920
rect 11839 26880 12440 26908
rect 11839 26877 11851 26880
rect 11793 26871 11851 26877
rect 9692 26840 9720 26871
rect 12434 26868 12440 26880
rect 12492 26868 12498 26920
rect 12805 26911 12863 26917
rect 12805 26877 12817 26911
rect 12851 26908 12863 26911
rect 12894 26908 12900 26920
rect 12851 26880 12900 26908
rect 12851 26877 12863 26880
rect 12805 26871 12863 26877
rect 12894 26868 12900 26880
rect 12952 26908 12958 26920
rect 13262 26908 13268 26920
rect 12952 26880 13268 26908
rect 12952 26868 12958 26880
rect 13262 26868 13268 26880
rect 13320 26868 13326 26920
rect 14277 26911 14335 26917
rect 14277 26877 14289 26911
rect 14323 26908 14335 26911
rect 19904 26908 19932 26948
rect 20162 26936 20168 26948
rect 20220 26936 20226 26988
rect 20346 26936 20352 26988
rect 20404 26976 20410 26988
rect 20533 26979 20591 26985
rect 20533 26976 20545 26979
rect 20404 26948 20545 26976
rect 20404 26936 20410 26948
rect 20533 26945 20545 26948
rect 20579 26976 20591 26979
rect 21269 26979 21327 26985
rect 20579 26948 21036 26976
rect 20579 26945 20591 26948
rect 20533 26939 20591 26945
rect 14323 26880 19932 26908
rect 20073 26911 20131 26917
rect 14323 26877 14335 26880
rect 14277 26871 14335 26877
rect 20073 26877 20085 26911
rect 20119 26908 20131 26911
rect 20714 26908 20720 26920
rect 20119 26880 20720 26908
rect 20119 26877 20131 26880
rect 20073 26871 20131 26877
rect 20714 26868 20720 26880
rect 20772 26868 20778 26920
rect 9858 26840 9864 26852
rect 6779 26812 7972 26840
rect 6779 26809 6791 26812
rect 6733 26803 6791 26809
rect 2038 26772 2044 26784
rect 1999 26744 2044 26772
rect 2038 26732 2044 26744
rect 2096 26732 2102 26784
rect 2590 26732 2596 26784
rect 2648 26772 2654 26784
rect 2685 26775 2743 26781
rect 2685 26772 2697 26775
rect 2648 26744 2697 26772
rect 2648 26732 2654 26744
rect 2685 26741 2697 26744
rect 2731 26741 2743 26775
rect 2685 26735 2743 26741
rect 4617 26775 4675 26781
rect 4617 26741 4629 26775
rect 4663 26772 4675 26775
rect 5074 26772 5080 26784
rect 4663 26744 5080 26772
rect 4663 26741 4675 26744
rect 4617 26735 4675 26741
rect 5074 26732 5080 26744
rect 5132 26732 5138 26784
rect 5905 26775 5963 26781
rect 5905 26741 5917 26775
rect 5951 26772 5963 26775
rect 6638 26772 6644 26784
rect 5951 26744 6644 26772
rect 5951 26741 5963 26744
rect 5905 26735 5963 26741
rect 6638 26732 6644 26744
rect 6696 26732 6702 26784
rect 7006 26732 7012 26784
rect 7064 26772 7070 26784
rect 7190 26772 7196 26784
rect 7064 26744 7196 26772
rect 7064 26732 7070 26744
rect 7190 26732 7196 26744
rect 7248 26732 7254 26784
rect 7374 26772 7380 26784
rect 7335 26744 7380 26772
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 7944 26772 7972 26812
rect 8128 26812 8708 26840
rect 8864 26812 9864 26840
rect 8128 26772 8156 26812
rect 7944 26744 8156 26772
rect 8680 26772 8708 26812
rect 9858 26800 9864 26812
rect 9916 26800 9922 26852
rect 12250 26800 12256 26852
rect 12308 26840 12314 26852
rect 15562 26840 15568 26852
rect 12308 26812 15568 26840
rect 12308 26800 12314 26812
rect 15562 26800 15568 26812
rect 15620 26800 15626 26852
rect 10686 26772 10692 26784
rect 8680 26744 10692 26772
rect 10686 26732 10692 26744
rect 10744 26732 10750 26784
rect 11054 26772 11060 26784
rect 11015 26744 11060 26772
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 13446 26732 13452 26784
rect 13504 26772 13510 26784
rect 13633 26775 13691 26781
rect 13633 26772 13645 26775
rect 13504 26744 13645 26772
rect 13504 26732 13510 26744
rect 13633 26741 13645 26744
rect 13679 26741 13691 26775
rect 14918 26772 14924 26784
rect 14879 26744 14924 26772
rect 13633 26735 13691 26741
rect 14918 26732 14924 26744
rect 14976 26732 14982 26784
rect 15194 26732 15200 26784
rect 15252 26772 15258 26784
rect 15749 26775 15807 26781
rect 15749 26772 15761 26775
rect 15252 26744 15761 26772
rect 15252 26732 15258 26744
rect 15749 26741 15761 26744
rect 15795 26741 15807 26775
rect 16942 26772 16948 26784
rect 16903 26744 16948 26772
rect 15749 26735 15807 26741
rect 16942 26732 16948 26744
rect 17000 26732 17006 26784
rect 17586 26772 17592 26784
rect 17547 26744 17592 26772
rect 17586 26732 17592 26744
rect 17644 26732 17650 26784
rect 18230 26772 18236 26784
rect 18191 26744 18236 26772
rect 18230 26732 18236 26744
rect 18288 26732 18294 26784
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 20625 26775 20683 26781
rect 20625 26772 20637 26775
rect 20496 26744 20637 26772
rect 20496 26732 20502 26744
rect 20625 26741 20637 26744
rect 20671 26741 20683 26775
rect 21008 26772 21036 26948
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 22002 26976 22008 26988
rect 21315 26948 22008 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 25774 26976 25780 26988
rect 25735 26948 25780 26976
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 21910 26868 21916 26920
rect 21968 26908 21974 26920
rect 22649 26911 22707 26917
rect 22649 26908 22661 26911
rect 21968 26880 22661 26908
rect 21968 26868 21974 26880
rect 22649 26877 22661 26880
rect 22695 26877 22707 26911
rect 22649 26871 22707 26877
rect 22925 26911 22983 26917
rect 22925 26877 22937 26911
rect 22971 26877 22983 26911
rect 22925 26871 22983 26877
rect 27617 26911 27675 26917
rect 27617 26877 27629 26911
rect 27663 26908 27675 26911
rect 27706 26908 27712 26920
rect 27663 26880 27712 26908
rect 27663 26877 27675 26880
rect 27617 26871 27675 26877
rect 21818 26800 21824 26852
rect 21876 26840 21882 26852
rect 22940 26840 22968 26871
rect 27706 26868 27712 26880
rect 27764 26868 27770 26920
rect 28629 26911 28687 26917
rect 28629 26877 28641 26911
rect 28675 26877 28687 26911
rect 28736 26908 28764 27084
rect 30742 27072 30748 27084
rect 30800 27072 30806 27124
rect 30834 27072 30840 27124
rect 30892 27112 30898 27124
rect 30892 27084 35894 27112
rect 30892 27072 30898 27084
rect 28810 27004 28816 27056
rect 28868 27044 28874 27056
rect 29273 27047 29331 27053
rect 29273 27044 29285 27047
rect 28868 27016 29285 27044
rect 28868 27004 28874 27016
rect 29273 27013 29285 27016
rect 29319 27013 29331 27047
rect 35866 27044 35894 27084
rect 38194 27044 38200 27056
rect 35866 27016 38200 27044
rect 29273 27007 29331 27013
rect 38194 27004 38200 27016
rect 38252 27004 38258 27056
rect 30653 26979 30711 26985
rect 30653 26945 30665 26979
rect 30699 26976 30711 26979
rect 38286 26976 38292 26988
rect 30699 26948 35894 26976
rect 38247 26948 38292 26976
rect 30699 26945 30711 26948
rect 30653 26939 30711 26945
rect 29181 26911 29239 26917
rect 29181 26908 29193 26911
rect 28736 26880 29193 26908
rect 28629 26871 28687 26877
rect 29181 26877 29193 26880
rect 29227 26908 29239 26911
rect 32030 26908 32036 26920
rect 29227 26880 32036 26908
rect 29227 26877 29239 26880
rect 29181 26871 29239 26877
rect 21876 26812 22968 26840
rect 28644 26840 28672 26871
rect 32030 26868 32036 26880
rect 32088 26868 32094 26920
rect 28644 26812 28764 26840
rect 21876 26800 21882 26812
rect 25866 26772 25872 26784
rect 21008 26744 25872 26772
rect 20625 26735 20683 26741
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 28736 26772 28764 26812
rect 28902 26800 28908 26852
rect 28960 26840 28966 26852
rect 29733 26843 29791 26849
rect 29733 26840 29745 26843
rect 28960 26812 29745 26840
rect 28960 26800 28966 26812
rect 29733 26809 29745 26812
rect 29779 26809 29791 26843
rect 35866 26840 35894 26948
rect 38286 26936 38292 26948
rect 38344 26936 38350 26988
rect 38105 26843 38163 26849
rect 38105 26840 38117 26843
rect 35866 26812 38117 26840
rect 29733 26803 29791 26809
rect 38105 26809 38117 26812
rect 38151 26809 38163 26843
rect 38105 26803 38163 26809
rect 28994 26772 29000 26784
rect 28736 26744 29000 26772
rect 28994 26732 29000 26744
rect 29052 26772 29058 26784
rect 29822 26772 29828 26784
rect 29052 26744 29828 26772
rect 29052 26732 29058 26744
rect 29822 26732 29828 26744
rect 29880 26732 29886 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 3326 26528 3332 26580
rect 3384 26568 3390 26580
rect 9306 26568 9312 26580
rect 3384 26540 9312 26568
rect 3384 26528 3390 26540
rect 9306 26528 9312 26540
rect 9364 26528 9370 26580
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 18785 26571 18843 26577
rect 18785 26568 18797 26571
rect 10100 26540 18797 26568
rect 10100 26528 10106 26540
rect 18785 26537 18797 26540
rect 18831 26537 18843 26571
rect 22186 26568 22192 26580
rect 18785 26531 18843 26537
rect 20640 26540 22192 26568
rect 4338 26500 4344 26512
rect 4080 26472 4344 26500
rect 2958 26432 2964 26444
rect 1596 26404 2964 26432
rect 1596 26373 1624 26404
rect 2958 26392 2964 26404
rect 3016 26392 3022 26444
rect 4080 26441 4108 26472
rect 4338 26460 4344 26472
rect 4396 26500 4402 26512
rect 4890 26500 4896 26512
rect 4396 26472 4896 26500
rect 4396 26460 4402 26472
rect 4890 26460 4896 26472
rect 4948 26460 4954 26512
rect 5074 26460 5080 26512
rect 5132 26500 5138 26512
rect 5132 26472 11836 26500
rect 5132 26460 5138 26472
rect 4065 26435 4123 26441
rect 4065 26401 4077 26435
rect 4111 26401 4123 26435
rect 4065 26395 4123 26401
rect 4154 26392 4160 26444
rect 4212 26432 4218 26444
rect 4706 26432 4712 26444
rect 4212 26404 4712 26432
rect 4212 26392 4218 26404
rect 4706 26392 4712 26404
rect 4764 26392 4770 26444
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26432 5319 26435
rect 10134 26432 10140 26444
rect 5307 26404 10140 26432
rect 5307 26401 5319 26404
rect 5261 26395 5319 26401
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 10778 26392 10784 26444
rect 10836 26432 10842 26444
rect 10965 26435 11023 26441
rect 10965 26432 10977 26435
rect 10836 26404 10977 26432
rect 10836 26392 10842 26404
rect 10965 26401 10977 26404
rect 11011 26401 11023 26435
rect 10965 26395 11023 26401
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26333 1639 26367
rect 1581 26327 1639 26333
rect 4890 26324 4896 26376
rect 4948 26364 4954 26376
rect 5169 26367 5227 26373
rect 5169 26364 5181 26367
rect 4948 26336 5181 26364
rect 4948 26324 4954 26336
rect 5169 26333 5181 26336
rect 5215 26333 5227 26367
rect 5810 26364 5816 26376
rect 5771 26336 5816 26364
rect 5169 26327 5227 26333
rect 5810 26324 5816 26336
rect 5868 26324 5874 26376
rect 6178 26324 6184 26376
rect 6236 26364 6242 26376
rect 6641 26367 6699 26373
rect 6641 26364 6653 26367
rect 6236 26336 6653 26364
rect 6236 26324 6242 26336
rect 6641 26333 6653 26336
rect 6687 26333 6699 26367
rect 9030 26364 9036 26376
rect 6641 26327 6699 26333
rect 8312 26336 9036 26364
rect 2685 26299 2743 26305
rect 2685 26265 2697 26299
rect 2731 26265 2743 26299
rect 2685 26259 2743 26265
rect 1762 26228 1768 26240
rect 1723 26200 1768 26228
rect 1762 26188 1768 26200
rect 1820 26188 1826 26240
rect 2700 26228 2728 26259
rect 2774 26256 2780 26308
rect 2832 26296 2838 26308
rect 3329 26299 3387 26305
rect 2832 26268 2877 26296
rect 2832 26256 2838 26268
rect 3329 26265 3341 26299
rect 3375 26296 3387 26299
rect 3375 26268 4108 26296
rect 3375 26265 3387 26268
rect 3329 26259 3387 26265
rect 2958 26228 2964 26240
rect 2700 26200 2964 26228
rect 2958 26188 2964 26200
rect 3016 26188 3022 26240
rect 4080 26228 4108 26268
rect 4154 26256 4160 26308
rect 4212 26296 4218 26308
rect 4709 26299 4767 26305
rect 4709 26296 4721 26299
rect 4212 26268 4257 26296
rect 4356 26268 4721 26296
rect 4212 26256 4218 26268
rect 4356 26228 4384 26268
rect 4709 26265 4721 26268
rect 4755 26296 4767 26299
rect 5718 26296 5724 26308
rect 4755 26268 5724 26296
rect 4755 26265 4767 26268
rect 4709 26259 4767 26265
rect 5718 26256 5724 26268
rect 5776 26256 5782 26308
rect 5905 26299 5963 26305
rect 5905 26265 5917 26299
rect 5951 26296 5963 26299
rect 7006 26296 7012 26308
rect 5951 26268 7012 26296
rect 5951 26265 5963 26268
rect 5905 26259 5963 26265
rect 7006 26256 7012 26268
rect 7064 26256 7070 26308
rect 7469 26299 7527 26305
rect 7469 26265 7481 26299
rect 7515 26265 7527 26299
rect 7469 26259 7527 26265
rect 7561 26299 7619 26305
rect 7561 26265 7573 26299
rect 7607 26296 7619 26299
rect 7926 26296 7932 26308
rect 7607 26268 7932 26296
rect 7607 26265 7619 26268
rect 7561 26259 7619 26265
rect 4080 26200 4384 26228
rect 6546 26188 6552 26240
rect 6604 26228 6610 26240
rect 6733 26231 6791 26237
rect 6733 26228 6745 26231
rect 6604 26200 6745 26228
rect 6604 26188 6610 26200
rect 6733 26197 6745 26200
rect 6779 26197 6791 26231
rect 7484 26228 7512 26259
rect 7926 26256 7932 26268
rect 7984 26256 7990 26308
rect 8018 26256 8024 26308
rect 8076 26296 8082 26308
rect 8312 26296 8340 26336
rect 9030 26324 9036 26336
rect 9088 26324 9094 26376
rect 9858 26324 9864 26376
rect 9916 26364 9922 26376
rect 11808 26364 11836 26472
rect 12434 26460 12440 26512
rect 12492 26500 12498 26512
rect 12492 26472 13400 26500
rect 12492 26460 12498 26472
rect 11974 26432 11980 26444
rect 11935 26404 11980 26432
rect 11974 26392 11980 26404
rect 12032 26392 12038 26444
rect 13081 26435 13139 26441
rect 13081 26401 13093 26435
rect 13127 26432 13139 26435
rect 13262 26432 13268 26444
rect 13127 26404 13268 26432
rect 13127 26401 13139 26404
rect 13081 26395 13139 26401
rect 13262 26392 13268 26404
rect 13320 26392 13326 26444
rect 13372 26441 13400 26472
rect 13998 26460 14004 26512
rect 14056 26500 14062 26512
rect 14056 26472 15056 26500
rect 14056 26460 14062 26472
rect 13357 26435 13415 26441
rect 13357 26401 13369 26435
rect 13403 26432 13415 26435
rect 14642 26432 14648 26444
rect 13403 26404 14648 26432
rect 13403 26401 13415 26404
rect 13357 26395 13415 26401
rect 14642 26392 14648 26404
rect 14700 26392 14706 26444
rect 12710 26364 12716 26376
rect 9916 26336 9961 26364
rect 11808 26336 12716 26364
rect 9916 26324 9922 26336
rect 12710 26324 12716 26336
rect 12768 26324 12774 26376
rect 8076 26268 8340 26296
rect 8481 26299 8539 26305
rect 8076 26256 8082 26268
rect 8481 26265 8493 26299
rect 8527 26265 8539 26299
rect 9048 26296 9076 26324
rect 9217 26299 9275 26305
rect 9217 26296 9229 26299
rect 9048 26268 9229 26296
rect 8481 26259 8539 26265
rect 9217 26265 9229 26268
rect 9263 26265 9275 26299
rect 9217 26259 9275 26265
rect 8036 26228 8064 26256
rect 7484 26200 8064 26228
rect 8496 26228 8524 26259
rect 9306 26256 9312 26308
rect 9364 26296 9370 26308
rect 9364 26268 9409 26296
rect 9364 26256 9370 26268
rect 10686 26256 10692 26308
rect 10744 26296 10750 26308
rect 11057 26299 11115 26305
rect 11057 26296 11069 26299
rect 10744 26268 11069 26296
rect 10744 26256 10750 26268
rect 11057 26265 11069 26268
rect 11103 26265 11115 26299
rect 11057 26259 11115 26265
rect 11790 26256 11796 26308
rect 11848 26296 11854 26308
rect 12434 26296 12440 26308
rect 11848 26268 12440 26296
rect 11848 26256 11854 26268
rect 12434 26256 12440 26268
rect 12492 26256 12498 26308
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 13173 26299 13231 26305
rect 13173 26296 13185 26299
rect 12584 26268 13185 26296
rect 12584 26256 12590 26268
rect 13173 26265 13185 26268
rect 13219 26265 13231 26299
rect 13173 26259 13231 26265
rect 13262 26256 13268 26308
rect 13320 26296 13326 26308
rect 13814 26296 13820 26308
rect 13320 26268 13820 26296
rect 13320 26256 13326 26268
rect 13814 26256 13820 26268
rect 13872 26256 13878 26308
rect 14366 26296 14372 26308
rect 14327 26268 14372 26296
rect 14366 26256 14372 26268
rect 14424 26256 14430 26308
rect 14458 26256 14464 26308
rect 14516 26296 14522 26308
rect 15028 26296 15056 26472
rect 15838 26460 15844 26512
rect 15896 26500 15902 26512
rect 15896 26472 16252 26500
rect 15896 26460 15902 26472
rect 15654 26392 15660 26444
rect 15712 26432 15718 26444
rect 16114 26432 16120 26444
rect 15712 26404 16120 26432
rect 15712 26392 15718 26404
rect 16114 26392 16120 26404
rect 16172 26392 16178 26444
rect 16224 26441 16252 26472
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26401 16267 26435
rect 16209 26395 16267 26401
rect 16574 26392 16580 26444
rect 16632 26432 16638 26444
rect 17770 26432 17776 26444
rect 16632 26404 17776 26432
rect 16632 26392 16638 26404
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 18138 26392 18144 26444
rect 18196 26432 18202 26444
rect 18782 26432 18788 26444
rect 18196 26404 18788 26432
rect 18196 26392 18202 26404
rect 18782 26392 18788 26404
rect 18840 26432 18846 26444
rect 20640 26441 20668 26540
rect 22186 26528 22192 26540
rect 22244 26528 22250 26580
rect 22370 26568 22376 26580
rect 22331 26540 22376 26568
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 26418 26528 26424 26580
rect 26476 26568 26482 26580
rect 26513 26571 26571 26577
rect 26513 26568 26525 26571
rect 26476 26540 26525 26568
rect 26476 26528 26482 26540
rect 26513 26537 26525 26540
rect 26559 26537 26571 26571
rect 27614 26568 27620 26580
rect 26513 26531 26571 26537
rect 26620 26540 27620 26568
rect 20806 26460 20812 26512
rect 20864 26500 20870 26512
rect 23017 26503 23075 26509
rect 23017 26500 23029 26503
rect 20864 26472 23029 26500
rect 20864 26460 20870 26472
rect 23017 26469 23029 26472
rect 23063 26469 23075 26503
rect 23017 26463 23075 26469
rect 19613 26435 19671 26441
rect 19613 26432 19625 26435
rect 18840 26404 19625 26432
rect 18840 26392 18846 26404
rect 19613 26401 19625 26404
rect 19659 26401 19671 26435
rect 19613 26395 19671 26401
rect 20625 26435 20683 26441
rect 20625 26401 20637 26435
rect 20671 26401 20683 26435
rect 20625 26395 20683 26401
rect 21177 26435 21235 26441
rect 21177 26401 21189 26435
rect 21223 26432 21235 26435
rect 22094 26432 22100 26444
rect 21223 26404 22100 26432
rect 21223 26401 21235 26404
rect 21177 26395 21235 26401
rect 22094 26392 22100 26404
rect 22152 26392 22158 26444
rect 22186 26392 22192 26444
rect 22244 26432 22250 26444
rect 23198 26432 23204 26444
rect 22244 26404 23204 26432
rect 22244 26392 22250 26404
rect 23198 26392 23204 26404
rect 23256 26392 23262 26444
rect 25774 26432 25780 26444
rect 25332 26404 25780 26432
rect 17129 26367 17187 26373
rect 17129 26364 17141 26367
rect 16592 26336 17141 26364
rect 16592 26308 16620 26336
rect 17129 26333 17141 26336
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17310 26324 17316 26376
rect 17368 26364 17374 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 17368 26336 18061 26364
rect 17368 26324 17374 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18690 26364 18696 26376
rect 18651 26336 18696 26364
rect 18049 26327 18107 26333
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 22278 26364 22284 26376
rect 22239 26336 22284 26364
rect 22278 26324 22284 26336
rect 22336 26324 22342 26376
rect 22922 26364 22928 26376
rect 22883 26336 22928 26364
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 25332 26373 25360 26404
rect 25774 26392 25780 26404
rect 25832 26432 25838 26444
rect 26620 26432 26648 26540
rect 27614 26528 27620 26540
rect 27672 26528 27678 26580
rect 28810 26568 28816 26580
rect 28771 26540 28816 26568
rect 28810 26528 28816 26540
rect 28868 26528 28874 26580
rect 37734 26568 37740 26580
rect 35866 26540 37740 26568
rect 35866 26500 35894 26540
rect 37734 26528 37740 26540
rect 37792 26528 37798 26580
rect 25832 26404 26648 26432
rect 27080 26472 35894 26500
rect 36357 26503 36415 26509
rect 25832 26392 25838 26404
rect 27080 26373 27108 26472
rect 36357 26469 36369 26503
rect 36403 26469 36415 26503
rect 38194 26500 38200 26512
rect 38155 26472 38200 26500
rect 36357 26463 36415 26469
rect 27706 26432 27712 26444
rect 27667 26404 27712 26432
rect 27706 26392 27712 26404
rect 27764 26392 27770 26444
rect 36372 26432 36400 26463
rect 38194 26460 38200 26472
rect 38252 26460 38258 26512
rect 36372 26404 38056 26432
rect 25317 26367 25375 26373
rect 25317 26333 25329 26367
rect 25363 26333 25375 26367
rect 25317 26327 25375 26333
rect 26421 26367 26479 26373
rect 26421 26333 26433 26367
rect 26467 26364 26479 26367
rect 27065 26367 27123 26373
rect 27065 26364 27077 26367
rect 26467 26336 27077 26364
rect 26467 26333 26479 26336
rect 26421 26327 26479 26333
rect 27065 26333 27077 26336
rect 27111 26333 27123 26367
rect 28718 26364 28724 26376
rect 28679 26336 28724 26364
rect 27065 26327 27123 26333
rect 28718 26324 28724 26336
rect 28776 26324 28782 26376
rect 36538 26364 36544 26376
rect 36499 26336 36544 26364
rect 36538 26324 36544 26336
rect 36596 26324 36602 26376
rect 38028 26373 38056 26404
rect 38013 26367 38071 26373
rect 38013 26333 38025 26367
rect 38059 26333 38071 26367
rect 38013 26327 38071 26333
rect 15749 26299 15807 26305
rect 15749 26296 15761 26299
rect 14516 26268 14561 26296
rect 15028 26268 15761 26296
rect 14516 26256 14522 26268
rect 15749 26265 15761 26268
rect 15795 26265 15807 26299
rect 15749 26259 15807 26265
rect 16574 26256 16580 26308
rect 16632 26256 16638 26308
rect 18141 26299 18199 26305
rect 18141 26265 18153 26299
rect 18187 26296 18199 26299
rect 19242 26296 19248 26308
rect 18187 26268 19248 26296
rect 18187 26265 18199 26268
rect 18141 26259 18199 26265
rect 19242 26256 19248 26268
rect 19300 26256 19306 26308
rect 19705 26299 19763 26305
rect 19705 26265 19717 26299
rect 19751 26296 19763 26299
rect 19978 26296 19984 26308
rect 19751 26268 19984 26296
rect 19751 26265 19763 26268
rect 19705 26259 19763 26265
rect 19978 26256 19984 26268
rect 20036 26256 20042 26308
rect 21269 26299 21327 26305
rect 21269 26265 21281 26299
rect 21315 26265 21327 26299
rect 21269 26259 21327 26265
rect 9030 26228 9036 26240
rect 8496 26200 9036 26228
rect 6733 26191 6791 26197
rect 9030 26188 9036 26200
rect 9088 26188 9094 26240
rect 9490 26188 9496 26240
rect 9548 26228 9554 26240
rect 13906 26228 13912 26240
rect 9548 26200 13912 26228
rect 9548 26188 9554 26200
rect 13906 26188 13912 26200
rect 13964 26188 13970 26240
rect 13998 26188 14004 26240
rect 14056 26228 14062 26240
rect 16592 26228 16620 26256
rect 17218 26228 17224 26240
rect 14056 26200 16620 26228
rect 17179 26200 17224 26228
rect 14056 26188 14062 26200
rect 17218 26188 17224 26200
rect 17276 26188 17282 26240
rect 21284 26228 21312 26259
rect 21358 26256 21364 26308
rect 21416 26296 21422 26308
rect 21821 26299 21879 26305
rect 21821 26296 21833 26299
rect 21416 26268 21833 26296
rect 21416 26256 21422 26268
rect 21821 26265 21833 26268
rect 21867 26265 21879 26299
rect 22940 26296 22968 26324
rect 30834 26296 30840 26308
rect 22940 26268 30840 26296
rect 21821 26259 21879 26265
rect 30834 26256 30840 26268
rect 30892 26256 30898 26308
rect 23382 26228 23388 26240
rect 21284 26200 23388 26228
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 25409 26231 25467 26237
rect 25409 26197 25421 26231
rect 25455 26228 25467 26231
rect 25590 26228 25596 26240
rect 25455 26200 25596 26228
rect 25455 26197 25467 26200
rect 25409 26191 25467 26197
rect 25590 26188 25596 26200
rect 25648 26188 25654 26240
rect 27157 26231 27215 26237
rect 27157 26197 27169 26231
rect 27203 26228 27215 26231
rect 27246 26228 27252 26240
rect 27203 26200 27252 26228
rect 27203 26197 27215 26200
rect 27157 26191 27215 26197
rect 27246 26188 27252 26200
rect 27304 26188 27310 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 2222 25984 2228 26036
rect 2280 26024 2286 26036
rect 2774 26024 2780 26036
rect 2280 25996 2780 26024
rect 2280 25984 2286 25996
rect 2774 25984 2780 25996
rect 2832 25984 2838 26036
rect 5258 26024 5264 26036
rect 4172 25996 5264 26024
rect 2314 25956 2320 25968
rect 2275 25928 2320 25956
rect 2314 25916 2320 25928
rect 2372 25916 2378 25968
rect 3418 25916 3424 25968
rect 3476 25956 3482 25968
rect 4062 25956 4068 25968
rect 3476 25928 4068 25956
rect 3476 25916 3482 25928
rect 4062 25916 4068 25928
rect 4120 25916 4126 25968
rect 4172 25965 4200 25996
rect 5258 25984 5264 25996
rect 5316 25984 5322 26036
rect 6733 26027 6791 26033
rect 6733 25993 6745 26027
rect 6779 26024 6791 26027
rect 6779 25996 11928 26024
rect 6779 25993 6791 25996
rect 6733 25987 6791 25993
rect 4157 25959 4215 25965
rect 4157 25925 4169 25959
rect 4203 25925 4215 25959
rect 4157 25919 4215 25925
rect 4246 25916 4252 25968
rect 4304 25956 4310 25968
rect 4304 25928 4752 25956
rect 4304 25916 4310 25928
rect 2222 25820 2228 25832
rect 2183 25792 2228 25820
rect 2222 25780 2228 25792
rect 2280 25780 2286 25832
rect 3237 25823 3295 25829
rect 3237 25789 3249 25823
rect 3283 25820 3295 25823
rect 3326 25820 3332 25832
rect 3283 25792 3332 25820
rect 3283 25789 3295 25792
rect 3237 25783 3295 25789
rect 3326 25780 3332 25792
rect 3384 25780 3390 25832
rect 4065 25823 4123 25829
rect 4065 25789 4077 25823
rect 4111 25789 4123 25823
rect 4338 25820 4344 25832
rect 4299 25792 4344 25820
rect 4065 25783 4123 25789
rect 4080 25752 4108 25783
rect 4338 25780 4344 25792
rect 4396 25780 4402 25832
rect 4724 25820 4752 25928
rect 4798 25916 4804 25968
rect 4856 25956 4862 25968
rect 5353 25959 5411 25965
rect 5353 25956 5365 25959
rect 4856 25928 5365 25956
rect 4856 25916 4862 25928
rect 5353 25925 5365 25928
rect 5399 25925 5411 25959
rect 8018 25956 8024 25968
rect 7979 25928 8024 25956
rect 5353 25919 5411 25925
rect 8018 25916 8024 25928
rect 8076 25916 8082 25968
rect 8113 25959 8171 25965
rect 8113 25925 8125 25959
rect 8159 25956 8171 25959
rect 8294 25956 8300 25968
rect 8159 25928 8300 25956
rect 8159 25925 8171 25928
rect 8113 25919 8171 25925
rect 8294 25916 8300 25928
rect 8352 25916 8358 25968
rect 8570 25916 8576 25968
rect 8628 25956 8634 25968
rect 8846 25956 8852 25968
rect 8628 25928 8852 25956
rect 8628 25916 8634 25928
rect 8846 25916 8852 25928
rect 8904 25916 8910 25968
rect 10134 25956 10140 25968
rect 10095 25928 10140 25956
rect 10134 25916 10140 25928
rect 10192 25916 10198 25968
rect 11330 25916 11336 25968
rect 11388 25956 11394 25968
rect 11900 25965 11928 25996
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 15838 26024 15844 26036
rect 12492 25996 15844 26024
rect 12492 25984 12498 25996
rect 15838 25984 15844 25996
rect 15896 26024 15902 26036
rect 16482 26024 16488 26036
rect 15896 25996 16488 26024
rect 15896 25984 15902 25996
rect 16482 25984 16488 25996
rect 16540 25984 16546 26036
rect 18322 25984 18328 26036
rect 18380 26024 18386 26036
rect 22738 26024 22744 26036
rect 18380 25996 22140 26024
rect 22699 25996 22744 26024
rect 18380 25984 18386 25996
rect 11793 25959 11851 25965
rect 11793 25956 11805 25959
rect 11388 25928 11805 25956
rect 11388 25916 11394 25928
rect 11793 25925 11805 25928
rect 11839 25925 11851 25959
rect 11793 25919 11851 25925
rect 11885 25959 11943 25965
rect 11885 25925 11897 25959
rect 11931 25925 11943 25959
rect 13998 25956 14004 25968
rect 11885 25919 11943 25925
rect 13280 25928 14004 25956
rect 6641 25891 6699 25897
rect 6641 25857 6653 25891
rect 6687 25857 6699 25891
rect 7282 25888 7288 25900
rect 7243 25860 7288 25888
rect 6641 25851 6699 25857
rect 5261 25823 5319 25829
rect 5261 25820 5273 25823
rect 4724 25792 5273 25820
rect 5261 25789 5273 25792
rect 5307 25789 5319 25823
rect 5902 25820 5908 25832
rect 5863 25792 5908 25820
rect 5261 25783 5319 25789
rect 5902 25780 5908 25792
rect 5960 25780 5966 25832
rect 6656 25820 6684 25851
rect 7282 25848 7288 25860
rect 7340 25848 7346 25900
rect 13280 25897 13308 25928
rect 13998 25916 14004 25928
rect 14056 25916 14062 25968
rect 15378 25916 15384 25968
rect 15436 25956 15442 25968
rect 16022 25956 16028 25968
rect 15436 25928 16028 25956
rect 15436 25916 15442 25928
rect 16022 25916 16028 25928
rect 16080 25916 16086 25968
rect 17773 25959 17831 25965
rect 17773 25925 17785 25959
rect 17819 25956 17831 25959
rect 19521 25959 19579 25965
rect 19521 25956 19533 25959
rect 17819 25928 19533 25956
rect 17819 25925 17831 25928
rect 17773 25919 17831 25925
rect 19521 25925 19533 25928
rect 19567 25925 19579 25959
rect 19521 25919 19579 25925
rect 20254 25916 20260 25968
rect 20312 25956 20318 25968
rect 20441 25959 20499 25965
rect 20441 25956 20453 25959
rect 20312 25928 20453 25956
rect 20312 25916 20318 25928
rect 20441 25925 20453 25928
rect 20487 25925 20499 25959
rect 20441 25919 20499 25925
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25857 13323 25891
rect 13906 25888 13912 25900
rect 13867 25860 13912 25888
rect 13265 25851 13323 25857
rect 13906 25848 13912 25860
rect 13964 25848 13970 25900
rect 14550 25888 14556 25900
rect 14511 25860 14556 25888
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 14826 25848 14832 25900
rect 14884 25888 14890 25900
rect 15194 25888 15200 25900
rect 14884 25860 15200 25888
rect 14884 25848 14890 25860
rect 15194 25848 15200 25860
rect 15252 25888 15258 25900
rect 15841 25891 15899 25897
rect 15841 25888 15853 25891
rect 15252 25860 15853 25888
rect 15252 25848 15258 25860
rect 15841 25857 15853 25860
rect 15887 25888 15899 25891
rect 16853 25891 16911 25897
rect 16853 25888 16865 25891
rect 15887 25860 16865 25888
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16853 25857 16865 25860
rect 16899 25857 16911 25891
rect 17678 25888 17684 25900
rect 17639 25860 17684 25888
rect 16853 25851 16911 25857
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 18322 25888 18328 25900
rect 18283 25860 18328 25888
rect 18322 25848 18328 25860
rect 18380 25848 18386 25900
rect 20806 25888 20812 25900
rect 20364 25860 20812 25888
rect 6914 25820 6920 25832
rect 6656 25792 6920 25820
rect 6914 25780 6920 25792
rect 6972 25780 6978 25832
rect 8386 25820 8392 25832
rect 8347 25792 8392 25820
rect 8386 25780 8392 25792
rect 8444 25780 8450 25832
rect 9122 25780 9128 25832
rect 9180 25820 9186 25832
rect 9582 25820 9588 25832
rect 9180 25792 9588 25820
rect 9180 25780 9186 25792
rect 9582 25780 9588 25792
rect 9640 25820 9646 25832
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 9640 25792 10057 25820
rect 9640 25780 9646 25792
rect 10045 25789 10057 25792
rect 10091 25789 10103 25823
rect 10318 25820 10324 25832
rect 10279 25792 10324 25820
rect 10045 25783 10103 25789
rect 10318 25780 10324 25792
rect 10376 25780 10382 25832
rect 12802 25820 12808 25832
rect 12176 25792 12808 25820
rect 5350 25752 5356 25764
rect 4080 25724 5356 25752
rect 5350 25712 5356 25724
rect 5408 25752 5414 25764
rect 5626 25752 5632 25764
rect 5408 25724 5632 25752
rect 5408 25712 5414 25724
rect 5626 25712 5632 25724
rect 5684 25712 5690 25764
rect 8404 25752 8432 25780
rect 12176 25752 12204 25792
rect 12802 25780 12808 25792
rect 12860 25780 12866 25832
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 15289 25823 15347 25829
rect 15289 25820 15301 25823
rect 13780 25792 15301 25820
rect 13780 25780 13786 25792
rect 15289 25789 15301 25792
rect 15335 25789 15347 25823
rect 15289 25783 15347 25789
rect 15562 25780 15568 25832
rect 15620 25820 15626 25832
rect 16945 25823 17003 25829
rect 16945 25820 16957 25823
rect 15620 25792 16957 25820
rect 15620 25780 15626 25792
rect 16945 25789 16957 25792
rect 16991 25789 17003 25823
rect 17696 25820 17724 25848
rect 19429 25823 19487 25829
rect 17696 25792 19380 25820
rect 16945 25783 17003 25789
rect 19352 25764 19380 25792
rect 19429 25789 19441 25823
rect 19475 25820 19487 25823
rect 20364 25820 20392 25860
rect 20806 25848 20812 25860
rect 20864 25848 20870 25900
rect 20901 25891 20959 25897
rect 20901 25857 20913 25891
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 19475 25792 20392 25820
rect 20916 25820 20944 25851
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 21818 25888 21824 25900
rect 21232 25860 21824 25888
rect 21232 25848 21238 25860
rect 21818 25848 21824 25860
rect 21876 25888 21882 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21876 25860 22017 25888
rect 21876 25848 21882 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22112 25888 22140 25996
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 23382 26024 23388 26036
rect 23343 25996 23388 26024
rect 23382 25984 23388 25996
rect 23440 25984 23446 26036
rect 24118 25984 24124 26036
rect 24176 26024 24182 26036
rect 28718 26024 28724 26036
rect 24176 25996 28724 26024
rect 24176 25984 24182 25996
rect 28718 25984 28724 25996
rect 28776 25984 28782 26036
rect 30653 26027 30711 26033
rect 30653 25993 30665 26027
rect 30699 26024 30711 26027
rect 33870 26024 33876 26036
rect 30699 25996 33876 26024
rect 30699 25993 30711 25996
rect 30653 25987 30711 25993
rect 33870 25984 33876 25996
rect 33928 25984 33934 26036
rect 25590 25956 25596 25968
rect 25551 25928 25596 25956
rect 25590 25916 25596 25928
rect 25648 25916 25654 25968
rect 27338 25956 27344 25968
rect 27299 25928 27344 25956
rect 27338 25916 27344 25928
rect 27396 25916 27402 25968
rect 27893 25959 27951 25965
rect 27893 25925 27905 25959
rect 27939 25956 27951 25959
rect 28902 25956 28908 25968
rect 27939 25928 28908 25956
rect 27939 25925 27951 25928
rect 27893 25919 27951 25925
rect 28902 25916 28908 25928
rect 28960 25916 28966 25968
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22112 25860 22661 25888
rect 22005 25851 22063 25857
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 21634 25820 21640 25832
rect 20916 25792 21640 25820
rect 19475 25789 19487 25792
rect 19429 25783 19487 25789
rect 8404 25724 12204 25752
rect 13630 25712 13636 25764
rect 13688 25752 13694 25764
rect 13906 25752 13912 25764
rect 13688 25724 13912 25752
rect 13688 25712 13694 25724
rect 13906 25712 13912 25724
rect 13964 25712 13970 25764
rect 14645 25755 14703 25761
rect 14645 25721 14657 25755
rect 14691 25752 14703 25755
rect 14691 25724 19288 25752
rect 14691 25721 14703 25724
rect 14645 25715 14703 25721
rect 2958 25644 2964 25696
rect 3016 25684 3022 25696
rect 5258 25684 5264 25696
rect 3016 25656 5264 25684
rect 3016 25644 3022 25656
rect 5258 25644 5264 25656
rect 5316 25644 5322 25696
rect 7377 25687 7435 25693
rect 7377 25653 7389 25687
rect 7423 25684 7435 25687
rect 10134 25684 10140 25696
rect 7423 25656 10140 25684
rect 7423 25653 7435 25656
rect 7377 25647 7435 25653
rect 10134 25644 10140 25656
rect 10192 25644 10198 25696
rect 13354 25684 13360 25696
rect 13315 25656 13360 25684
rect 13354 25644 13360 25656
rect 13412 25644 13418 25696
rect 14001 25687 14059 25693
rect 14001 25653 14013 25687
rect 14047 25684 14059 25687
rect 15378 25684 15384 25696
rect 14047 25656 15384 25684
rect 14047 25653 14059 25656
rect 14001 25647 14059 25653
rect 15378 25644 15384 25656
rect 15436 25644 15442 25696
rect 15930 25684 15936 25696
rect 15891 25656 15936 25684
rect 15930 25644 15936 25656
rect 15988 25644 15994 25696
rect 18417 25687 18475 25693
rect 18417 25653 18429 25687
rect 18463 25684 18475 25687
rect 18874 25684 18880 25696
rect 18463 25656 18880 25684
rect 18463 25653 18475 25656
rect 18417 25647 18475 25653
rect 18874 25644 18880 25656
rect 18932 25644 18938 25696
rect 19260 25684 19288 25724
rect 19334 25712 19340 25764
rect 19392 25712 19398 25764
rect 19518 25712 19524 25764
rect 19576 25752 19582 25764
rect 20916 25752 20944 25792
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22664 25820 22692 25851
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 23293 25891 23351 25897
rect 23293 25888 23305 25891
rect 23164 25860 23305 25888
rect 23164 25848 23170 25860
rect 23293 25857 23305 25860
rect 23339 25888 23351 25891
rect 24210 25888 24216 25900
rect 23339 25860 24216 25888
rect 23339 25857 23351 25860
rect 23293 25851 23351 25857
rect 24210 25848 24216 25860
rect 24268 25848 24274 25900
rect 30561 25891 30619 25897
rect 30561 25857 30573 25891
rect 30607 25888 30619 25891
rect 30834 25888 30840 25900
rect 30607 25860 30840 25888
rect 30607 25857 30619 25860
rect 30561 25851 30619 25857
rect 30834 25848 30840 25860
rect 30892 25848 30898 25900
rect 23750 25820 23756 25832
rect 22664 25792 23756 25820
rect 23750 25780 23756 25792
rect 23808 25780 23814 25832
rect 25501 25823 25559 25829
rect 25501 25789 25513 25823
rect 25547 25820 25559 25823
rect 26329 25823 26387 25829
rect 25547 25792 26280 25820
rect 25547 25789 25559 25792
rect 25501 25783 25559 25789
rect 26252 25764 26280 25792
rect 26329 25789 26341 25823
rect 26375 25789 26387 25823
rect 27246 25820 27252 25832
rect 27207 25792 27252 25820
rect 26329 25783 26387 25789
rect 19576 25724 20944 25752
rect 19576 25712 19582 25724
rect 21082 25712 21088 25764
rect 21140 25752 21146 25764
rect 22646 25752 22652 25764
rect 21140 25724 22652 25752
rect 21140 25712 21146 25724
rect 22646 25712 22652 25724
rect 22704 25712 22710 25764
rect 26234 25712 26240 25764
rect 26292 25712 26298 25764
rect 19426 25684 19432 25696
rect 19260 25656 19432 25684
rect 19426 25644 19432 25656
rect 19484 25644 19490 25696
rect 20990 25684 20996 25696
rect 20951 25656 20996 25684
rect 20990 25644 20996 25656
rect 21048 25644 21054 25696
rect 22097 25687 22155 25693
rect 22097 25653 22109 25687
rect 22143 25684 22155 25687
rect 22186 25684 22192 25696
rect 22143 25656 22192 25684
rect 22143 25653 22155 25656
rect 22097 25647 22155 25653
rect 22186 25644 22192 25656
rect 22244 25644 22250 25696
rect 24394 25644 24400 25696
rect 24452 25684 24458 25696
rect 26344 25684 26372 25783
rect 27246 25780 27252 25792
rect 27304 25780 27310 25832
rect 24452 25656 26372 25684
rect 24452 25644 24458 25656
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1486 25440 1492 25492
rect 1544 25480 1550 25492
rect 1765 25483 1823 25489
rect 1765 25480 1777 25483
rect 1544 25452 1777 25480
rect 1544 25440 1550 25452
rect 1765 25449 1777 25452
rect 1811 25449 1823 25483
rect 1765 25443 1823 25449
rect 3326 25440 3332 25492
rect 3384 25480 3390 25492
rect 5718 25480 5724 25492
rect 3384 25452 5724 25480
rect 3384 25440 3390 25452
rect 5718 25440 5724 25452
rect 5776 25480 5782 25492
rect 6270 25480 6276 25492
rect 5776 25452 6276 25480
rect 5776 25440 5782 25452
rect 6270 25440 6276 25452
rect 6328 25440 6334 25492
rect 6730 25440 6736 25492
rect 6788 25480 6794 25492
rect 7282 25480 7288 25492
rect 6788 25452 7288 25480
rect 6788 25440 6794 25452
rect 7282 25440 7288 25452
rect 7340 25440 7346 25492
rect 9490 25440 9496 25492
rect 9548 25480 9554 25492
rect 15470 25480 15476 25492
rect 9548 25452 15476 25480
rect 9548 25440 9554 25452
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 15565 25483 15623 25489
rect 15565 25449 15577 25483
rect 15611 25480 15623 25483
rect 16206 25480 16212 25492
rect 15611 25452 16212 25480
rect 15611 25449 15623 25452
rect 15565 25443 15623 25449
rect 16206 25440 16212 25452
rect 16264 25440 16270 25492
rect 16482 25440 16488 25492
rect 16540 25480 16546 25492
rect 19794 25480 19800 25492
rect 16540 25452 19800 25480
rect 16540 25440 16546 25452
rect 19794 25440 19800 25452
rect 19852 25440 19858 25492
rect 22278 25440 22284 25492
rect 22336 25480 22342 25492
rect 27522 25480 27528 25492
rect 22336 25452 27528 25480
rect 22336 25440 22342 25452
rect 27522 25440 27528 25452
rect 27580 25440 27586 25492
rect 27614 25440 27620 25492
rect 27672 25480 27678 25492
rect 29454 25480 29460 25492
rect 27672 25452 29460 25480
rect 27672 25440 27678 25452
rect 29454 25440 29460 25452
rect 29512 25440 29518 25492
rect 29914 25480 29920 25492
rect 29875 25452 29920 25480
rect 29914 25440 29920 25452
rect 29972 25440 29978 25492
rect 5994 25412 6000 25424
rect 4908 25384 6000 25412
rect 4908 25353 4936 25384
rect 5994 25372 6000 25384
rect 6052 25372 6058 25424
rect 8110 25372 8116 25424
rect 8168 25412 8174 25424
rect 9306 25412 9312 25424
rect 8168 25384 9312 25412
rect 8168 25372 8174 25384
rect 9306 25372 9312 25384
rect 9364 25372 9370 25424
rect 10888 25384 11468 25412
rect 4893 25347 4951 25353
rect 4893 25313 4905 25347
rect 4939 25313 4951 25347
rect 4893 25307 4951 25313
rect 5258 25304 5264 25356
rect 5316 25344 5322 25356
rect 5905 25347 5963 25353
rect 5905 25344 5917 25347
rect 5316 25316 5917 25344
rect 5316 25304 5322 25316
rect 5905 25313 5917 25316
rect 5951 25313 5963 25347
rect 6012 25344 6040 25372
rect 9122 25344 9128 25356
rect 6012 25316 9128 25344
rect 5905 25307 5963 25313
rect 1946 25276 1952 25288
rect 1907 25248 1952 25276
rect 1946 25236 1952 25248
rect 2004 25236 2010 25288
rect 4154 25276 4160 25288
rect 4115 25248 4160 25276
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25276 4307 25279
rect 4706 25276 4712 25288
rect 4295 25248 4712 25276
rect 4295 25245 4307 25248
rect 4249 25239 4307 25245
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 5920 25276 5948 25307
rect 9122 25304 9128 25316
rect 9180 25304 9186 25356
rect 9678 25347 9736 25353
rect 9678 25313 9690 25347
rect 9724 25344 9736 25347
rect 10226 25344 10232 25356
rect 9724 25316 10232 25344
rect 9724 25313 9736 25316
rect 9678 25307 9736 25313
rect 10226 25304 10232 25316
rect 10284 25304 10290 25356
rect 6270 25276 6276 25288
rect 5920 25248 6276 25276
rect 6270 25236 6276 25248
rect 6328 25236 6334 25288
rect 6365 25279 6423 25285
rect 6365 25245 6377 25279
rect 6411 25245 6423 25279
rect 9490 25276 9496 25288
rect 7774 25248 9496 25276
rect 6365 25239 6423 25245
rect 2501 25211 2559 25217
rect 2501 25177 2513 25211
rect 2547 25177 2559 25211
rect 3234 25208 3240 25220
rect 3195 25180 3240 25208
rect 2501 25171 2559 25177
rect 2516 25140 2544 25171
rect 3234 25168 3240 25180
rect 3292 25168 3298 25220
rect 4982 25168 4988 25220
rect 5040 25208 5046 25220
rect 6380 25208 6408 25239
rect 9490 25236 9496 25248
rect 9548 25236 9554 25288
rect 10888 25276 10916 25384
rect 11440 25344 11468 25384
rect 12636 25384 15056 25412
rect 12636 25344 12664 25384
rect 11440 25316 12664 25344
rect 13998 25304 14004 25356
rect 14056 25344 14062 25356
rect 14660 25344 14872 25356
rect 14921 25347 14979 25353
rect 14921 25344 14933 25347
rect 14056 25328 14933 25344
rect 14056 25316 14688 25328
rect 14844 25316 14933 25328
rect 14056 25304 14062 25316
rect 14921 25313 14933 25316
rect 14967 25313 14979 25347
rect 15028 25344 15056 25384
rect 15194 25372 15200 25424
rect 15252 25412 15258 25424
rect 21085 25415 21143 25421
rect 15252 25384 21036 25412
rect 15252 25372 15258 25384
rect 15028 25316 18828 25344
rect 14921 25307 14979 25313
rect 11330 25276 11336 25288
rect 10612 25248 10916 25276
rect 11291 25248 11336 25276
rect 6641 25211 6699 25217
rect 5040 25180 5085 25208
rect 6380 25180 6500 25208
rect 5040 25168 5046 25180
rect 4522 25140 4528 25152
rect 2516 25112 4528 25140
rect 4522 25100 4528 25112
rect 4580 25100 4586 25152
rect 6472 25140 6500 25180
rect 6641 25177 6653 25211
rect 6687 25208 6699 25211
rect 8662 25208 8668 25220
rect 6687 25180 7052 25208
rect 6687 25177 6699 25180
rect 6641 25171 6699 25177
rect 6822 25140 6828 25152
rect 6472 25112 6828 25140
rect 6822 25100 6828 25112
rect 6880 25100 6886 25152
rect 7024 25140 7052 25180
rect 7944 25180 8668 25208
rect 7944 25140 7972 25180
rect 8662 25168 8668 25180
rect 8720 25168 8726 25220
rect 9762 25211 9820 25217
rect 9762 25208 9774 25211
rect 9416 25180 9774 25208
rect 8110 25140 8116 25152
rect 7024 25112 7972 25140
rect 8071 25112 8116 25140
rect 8110 25100 8116 25112
rect 8168 25100 8174 25152
rect 8202 25100 8208 25152
rect 8260 25140 8266 25152
rect 9416 25140 9444 25180
rect 9762 25177 9774 25180
rect 9808 25177 9820 25211
rect 9762 25171 9820 25177
rect 8260 25112 9444 25140
rect 8260 25100 8266 25112
rect 9490 25100 9496 25152
rect 9548 25140 9554 25152
rect 10612 25140 10640 25248
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 13538 25276 13544 25288
rect 13499 25248 13544 25276
rect 13538 25236 13544 25248
rect 13596 25236 13602 25288
rect 14826 25285 14832 25288
rect 14821 25276 14832 25285
rect 14787 25248 14832 25276
rect 14821 25239 14832 25248
rect 14826 25236 14832 25239
rect 14884 25236 14890 25288
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25276 15531 25279
rect 15838 25276 15844 25288
rect 15519 25248 15844 25276
rect 15519 25245 15531 25248
rect 15473 25239 15531 25245
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18049 25279 18107 25285
rect 18049 25276 18061 25279
rect 18012 25248 18061 25276
rect 18012 25236 18018 25248
rect 18049 25245 18061 25248
rect 18095 25245 18107 25279
rect 18690 25276 18696 25288
rect 18603 25248 18696 25276
rect 18049 25239 18107 25245
rect 18690 25236 18696 25248
rect 18748 25236 18754 25288
rect 18800 25276 18828 25316
rect 18966 25304 18972 25356
rect 19024 25344 19030 25356
rect 19521 25347 19579 25353
rect 19521 25344 19533 25347
rect 19024 25316 19533 25344
rect 19024 25304 19030 25316
rect 19521 25313 19533 25316
rect 19567 25313 19579 25347
rect 19794 25344 19800 25356
rect 19755 25316 19800 25344
rect 19521 25307 19579 25313
rect 19794 25304 19800 25316
rect 19852 25304 19858 25356
rect 21008 25285 21036 25384
rect 21085 25381 21097 25415
rect 21131 25412 21143 25415
rect 28626 25412 28632 25424
rect 21131 25384 28632 25412
rect 21131 25381 21143 25384
rect 21085 25375 21143 25381
rect 28626 25372 28632 25384
rect 28684 25372 28690 25424
rect 22097 25347 22155 25353
rect 22097 25313 22109 25347
rect 22143 25344 22155 25347
rect 22186 25344 22192 25356
rect 22143 25316 22192 25344
rect 22143 25313 22155 25316
rect 22097 25307 22155 25313
rect 22186 25304 22192 25316
rect 22244 25304 22250 25356
rect 22370 25344 22376 25356
rect 22331 25316 22376 25344
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 26234 25344 26240 25356
rect 26147 25316 26240 25344
rect 26234 25304 26240 25316
rect 26292 25344 26298 25356
rect 27246 25344 27252 25356
rect 26292 25316 27252 25344
rect 26292 25304 26298 25316
rect 27246 25304 27252 25316
rect 27304 25304 27310 25356
rect 36538 25344 36544 25356
rect 28552 25316 36544 25344
rect 28552 25285 28580 25316
rect 36538 25304 36544 25316
rect 36596 25304 36602 25356
rect 20993 25279 21051 25285
rect 18800 25248 19334 25276
rect 10689 25211 10747 25217
rect 10689 25177 10701 25211
rect 10735 25208 10747 25211
rect 10870 25208 10876 25220
rect 10735 25180 10876 25208
rect 10735 25177 10747 25180
rect 10689 25171 10747 25177
rect 10870 25168 10876 25180
rect 10928 25168 10934 25220
rect 11606 25208 11612 25220
rect 11567 25180 11612 25208
rect 11606 25168 11612 25180
rect 11664 25168 11670 25220
rect 15930 25208 15936 25220
rect 12834 25180 15936 25208
rect 15930 25168 15936 25180
rect 15988 25168 15994 25220
rect 16209 25211 16267 25217
rect 16209 25177 16221 25211
rect 16255 25177 16267 25211
rect 16209 25171 16267 25177
rect 9548 25112 10640 25140
rect 10888 25140 10916 25168
rect 12434 25140 12440 25152
rect 10888 25112 12440 25140
rect 9548 25100 9554 25112
rect 12434 25100 12440 25112
rect 12492 25100 12498 25152
rect 12526 25100 12532 25152
rect 12584 25140 12590 25152
rect 13081 25143 13139 25149
rect 13081 25140 13093 25143
rect 12584 25112 13093 25140
rect 12584 25100 12590 25112
rect 13081 25109 13093 25112
rect 13127 25109 13139 25143
rect 13630 25140 13636 25152
rect 13591 25112 13636 25140
rect 13081 25103 13139 25109
rect 13630 25100 13636 25112
rect 13688 25100 13694 25152
rect 13814 25100 13820 25152
rect 13872 25140 13878 25152
rect 16224 25140 16252 25171
rect 16298 25168 16304 25220
rect 16356 25208 16362 25220
rect 17221 25211 17279 25217
rect 16356 25180 16401 25208
rect 16356 25168 16362 25180
rect 17221 25177 17233 25211
rect 17267 25208 17279 25211
rect 17494 25208 17500 25220
rect 17267 25180 17500 25208
rect 17267 25177 17279 25180
rect 17221 25171 17279 25177
rect 17494 25168 17500 25180
rect 17552 25168 17558 25220
rect 18708 25208 18736 25236
rect 18064 25180 18736 25208
rect 19306 25208 19334 25248
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25245 23811 25279
rect 23753 25239 23811 25245
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25245 28595 25279
rect 28537 25239 28595 25245
rect 19518 25208 19524 25220
rect 19306 25180 19524 25208
rect 13872 25112 16252 25140
rect 13872 25100 13878 25112
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 18064 25140 18092 25180
rect 19518 25168 19524 25180
rect 19576 25168 19582 25220
rect 19613 25211 19671 25217
rect 19613 25177 19625 25211
rect 19659 25177 19671 25211
rect 19613 25171 19671 25177
rect 22189 25211 22247 25217
rect 22189 25177 22201 25211
rect 22235 25208 22247 25211
rect 22278 25208 22284 25220
rect 22235 25180 22284 25208
rect 22235 25177 22247 25180
rect 22189 25171 22247 25177
rect 16632 25112 18092 25140
rect 18141 25143 18199 25149
rect 16632 25100 16638 25112
rect 18141 25109 18153 25143
rect 18187 25140 18199 25143
rect 18230 25140 18236 25152
rect 18187 25112 18236 25140
rect 18187 25109 18199 25112
rect 18141 25103 18199 25109
rect 18230 25100 18236 25112
rect 18288 25100 18294 25152
rect 18782 25140 18788 25152
rect 18743 25112 18788 25140
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 19334 25100 19340 25152
rect 19392 25140 19398 25152
rect 19621 25140 19649 25171
rect 22278 25168 22284 25180
rect 22336 25168 22342 25220
rect 22462 25168 22468 25220
rect 22520 25208 22526 25220
rect 23768 25208 23796 25239
rect 29086 25236 29092 25288
rect 29144 25276 29150 25288
rect 30101 25279 30159 25285
rect 30101 25276 30113 25279
rect 29144 25248 30113 25276
rect 29144 25236 29150 25248
rect 30101 25245 30113 25248
rect 30147 25245 30159 25279
rect 30101 25239 30159 25245
rect 38013 25279 38071 25285
rect 38013 25245 38025 25279
rect 38059 25245 38071 25279
rect 38013 25239 38071 25245
rect 22520 25180 23796 25208
rect 26329 25211 26387 25217
rect 22520 25168 22526 25180
rect 26329 25177 26341 25211
rect 26375 25208 26387 25211
rect 26694 25208 26700 25220
rect 26375 25180 26700 25208
rect 26375 25177 26387 25180
rect 26329 25171 26387 25177
rect 26694 25168 26700 25180
rect 26752 25168 26758 25220
rect 26881 25211 26939 25217
rect 26881 25177 26893 25211
rect 26927 25177 26939 25211
rect 37642 25208 37648 25220
rect 37603 25180 37648 25208
rect 26881 25171 26939 25177
rect 19392 25112 19649 25140
rect 23845 25143 23903 25149
rect 19392 25100 19398 25112
rect 23845 25109 23857 25143
rect 23891 25140 23903 25143
rect 25038 25140 25044 25152
rect 23891 25112 25044 25140
rect 23891 25109 23903 25112
rect 23845 25103 23903 25109
rect 25038 25100 25044 25112
rect 25096 25100 25102 25152
rect 26050 25100 26056 25152
rect 26108 25140 26114 25152
rect 26896 25140 26924 25171
rect 37642 25168 37648 25180
rect 37700 25208 37706 25220
rect 38028 25208 38056 25239
rect 37700 25180 38056 25208
rect 37700 25168 37706 25180
rect 26108 25112 26924 25140
rect 26108 25100 26114 25112
rect 27062 25100 27068 25152
rect 27120 25140 27126 25152
rect 28629 25143 28687 25149
rect 28629 25140 28641 25143
rect 27120 25112 28641 25140
rect 27120 25100 27126 25112
rect 28629 25109 28641 25112
rect 28675 25109 28687 25143
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 28629 25103 28687 25109
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1946 24896 1952 24948
rect 2004 24936 2010 24948
rect 4430 24936 4436 24948
rect 2004 24908 4436 24936
rect 2004 24896 2010 24908
rect 4430 24896 4436 24908
rect 4488 24896 4494 24948
rect 4706 24896 4712 24948
rect 4764 24936 4770 24948
rect 8202 24936 8208 24948
rect 4764 24908 8208 24936
rect 4764 24896 4770 24908
rect 8202 24896 8208 24908
rect 8260 24896 8266 24948
rect 8294 24896 8300 24948
rect 8352 24936 8358 24948
rect 18782 24936 18788 24948
rect 8352 24908 18788 24936
rect 8352 24896 8358 24908
rect 18782 24896 18788 24908
rect 18840 24896 18846 24948
rect 20254 24936 20260 24948
rect 19168 24908 20260 24936
rect 1762 24828 1768 24880
rect 1820 24868 1826 24880
rect 1857 24871 1915 24877
rect 1857 24868 1869 24871
rect 1820 24840 1869 24868
rect 1820 24828 1826 24840
rect 1857 24837 1869 24840
rect 1903 24837 1915 24871
rect 1857 24831 1915 24837
rect 2314 24828 2320 24880
rect 2372 24868 2378 24880
rect 3418 24868 3424 24880
rect 2372 24840 3424 24868
rect 2372 24828 2378 24840
rect 3418 24828 3424 24840
rect 3476 24828 3482 24880
rect 4249 24871 4307 24877
rect 4249 24837 4261 24871
rect 4295 24868 4307 24871
rect 4614 24868 4620 24880
rect 4295 24840 4620 24868
rect 4295 24837 4307 24840
rect 4249 24831 4307 24837
rect 4614 24828 4620 24840
rect 4672 24828 4678 24880
rect 5169 24871 5227 24877
rect 5169 24837 5181 24871
rect 5215 24868 5227 24871
rect 5258 24868 5264 24880
rect 5215 24840 5264 24868
rect 5215 24837 5227 24840
rect 5169 24831 5227 24837
rect 5258 24828 5264 24840
rect 5316 24828 5322 24880
rect 5994 24828 6000 24880
rect 6052 24868 6058 24880
rect 6733 24871 6791 24877
rect 6733 24868 6745 24871
rect 6052 24840 6745 24868
rect 6052 24828 6058 24840
rect 6733 24837 6745 24840
rect 6779 24837 6791 24871
rect 6733 24831 6791 24837
rect 7282 24828 7288 24880
rect 7340 24868 7346 24880
rect 8665 24871 8723 24877
rect 8665 24868 8677 24871
rect 7340 24840 8677 24868
rect 7340 24828 7346 24840
rect 8665 24837 8677 24840
rect 8711 24837 8723 24871
rect 11238 24868 11244 24880
rect 9890 24840 11244 24868
rect 8665 24831 8723 24837
rect 11238 24828 11244 24840
rect 11296 24828 11302 24880
rect 11698 24828 11704 24880
rect 11756 24868 11762 24880
rect 11977 24871 12035 24877
rect 11977 24868 11989 24871
rect 11756 24840 11989 24868
rect 11756 24828 11762 24840
rect 11977 24837 11989 24840
rect 12023 24837 12035 24871
rect 13722 24868 13728 24880
rect 13202 24840 13728 24868
rect 11977 24831 12035 24837
rect 13722 24828 13728 24840
rect 13780 24828 13786 24880
rect 14090 24868 14096 24880
rect 14051 24840 14096 24868
rect 14090 24828 14096 24840
rect 14148 24828 14154 24880
rect 15746 24868 15752 24880
rect 15707 24840 15752 24868
rect 15746 24828 15752 24840
rect 15804 24828 15810 24880
rect 17034 24868 17040 24880
rect 16995 24840 17040 24868
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 17494 24828 17500 24880
rect 17552 24868 17558 24880
rect 17957 24871 18015 24877
rect 17957 24868 17969 24871
rect 17552 24840 17969 24868
rect 17552 24828 17558 24840
rect 17957 24837 17969 24840
rect 18003 24868 18015 24871
rect 19168 24868 19196 24908
rect 20254 24896 20260 24908
rect 20312 24896 20318 24948
rect 22278 24896 22284 24948
rect 22336 24936 22342 24948
rect 22741 24939 22799 24945
rect 22741 24936 22753 24939
rect 22336 24908 22753 24936
rect 22336 24896 22342 24908
rect 22741 24905 22753 24908
rect 22787 24905 22799 24939
rect 22741 24899 22799 24905
rect 23198 24896 23204 24948
rect 23256 24936 23262 24948
rect 26421 24939 26479 24945
rect 23256 24908 24440 24936
rect 23256 24896 23262 24908
rect 24412 24880 24440 24908
rect 26421 24905 26433 24939
rect 26467 24936 26479 24939
rect 27338 24936 27344 24948
rect 26467 24908 27344 24936
rect 26467 24905 26479 24908
rect 26421 24899 26479 24905
rect 27338 24896 27344 24908
rect 27396 24896 27402 24948
rect 18003 24840 19196 24868
rect 18003 24837 18015 24840
rect 17957 24831 18015 24837
rect 19242 24828 19248 24880
rect 19300 24868 19306 24880
rect 19337 24871 19395 24877
rect 19337 24868 19349 24871
rect 19300 24840 19349 24868
rect 19300 24828 19306 24840
rect 19337 24837 19349 24840
rect 19383 24837 19395 24871
rect 20806 24868 20812 24880
rect 20767 24840 20812 24868
rect 19337 24831 19395 24837
rect 20806 24828 20812 24840
rect 20864 24828 20870 24880
rect 20901 24871 20959 24877
rect 20901 24837 20913 24871
rect 20947 24868 20959 24871
rect 20990 24868 20996 24880
rect 20947 24840 20996 24868
rect 20947 24837 20959 24840
rect 20901 24831 20959 24837
rect 20990 24828 20996 24840
rect 21048 24828 21054 24880
rect 23474 24868 23480 24880
rect 22572 24840 22784 24868
rect 23435 24840 23480 24868
rect 3237 24803 3295 24809
rect 3237 24769 3249 24803
rect 3283 24800 3295 24803
rect 3694 24800 3700 24812
rect 3283 24772 3700 24800
rect 3283 24769 3295 24772
rect 3237 24763 3295 24769
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 7742 24800 7748 24812
rect 7703 24772 7748 24800
rect 7742 24760 7748 24772
rect 7800 24760 7806 24812
rect 10594 24760 10600 24812
rect 10652 24800 10658 24812
rect 10965 24803 11023 24809
rect 10965 24800 10977 24803
rect 10652 24772 10977 24800
rect 10652 24760 10658 24772
rect 10965 24769 10977 24772
rect 11011 24769 11023 24803
rect 10965 24763 11023 24769
rect 14936 24772 15516 24800
rect 1765 24735 1823 24741
rect 1765 24701 1777 24735
rect 1811 24732 1823 24735
rect 1854 24732 1860 24744
rect 1811 24704 1860 24732
rect 1811 24701 1823 24704
rect 1765 24695 1823 24701
rect 1854 24692 1860 24704
rect 1912 24692 1918 24744
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24701 2835 24735
rect 2777 24695 2835 24701
rect 4157 24735 4215 24741
rect 4157 24701 4169 24735
rect 4203 24732 4215 24735
rect 4982 24732 4988 24744
rect 4203 24704 4988 24732
rect 4203 24701 4215 24704
rect 4157 24695 4215 24701
rect 2792 24664 2820 24695
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 5813 24735 5871 24741
rect 5813 24701 5825 24735
rect 5859 24701 5871 24735
rect 5813 24695 5871 24701
rect 4614 24664 4620 24676
rect 2792 24636 4620 24664
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 3418 24596 3424 24608
rect 3379 24568 3424 24596
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 4522 24556 4528 24608
rect 4580 24596 4586 24608
rect 5258 24596 5264 24608
rect 4580 24568 5264 24596
rect 4580 24556 4586 24568
rect 5258 24556 5264 24568
rect 5316 24556 5322 24608
rect 5828 24596 5856 24695
rect 5902 24692 5908 24744
rect 5960 24732 5966 24744
rect 6641 24735 6699 24741
rect 6641 24732 6653 24735
rect 5960 24704 6653 24732
rect 5960 24692 5966 24704
rect 6641 24701 6653 24704
rect 6687 24701 6699 24735
rect 8386 24732 8392 24744
rect 8347 24704 8392 24732
rect 6641 24695 6699 24701
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 9122 24692 9128 24744
rect 9180 24732 9186 24744
rect 9180 24704 9720 24732
rect 9180 24692 9186 24704
rect 7190 24664 7196 24676
rect 7151 24636 7196 24664
rect 7190 24624 7196 24636
rect 7248 24624 7254 24676
rect 9692 24664 9720 24704
rect 11330 24692 11336 24744
rect 11388 24732 11394 24744
rect 11701 24735 11759 24741
rect 11701 24732 11713 24735
rect 11388 24704 11713 24732
rect 11388 24692 11394 24704
rect 11701 24701 11713 24704
rect 11747 24701 11759 24735
rect 13722 24732 13728 24744
rect 11701 24695 11759 24701
rect 11808 24704 13728 24732
rect 10137 24667 10195 24673
rect 10137 24664 10149 24667
rect 7760 24636 8340 24664
rect 9692 24636 10149 24664
rect 7760 24596 7788 24636
rect 5828 24568 7788 24596
rect 7837 24599 7895 24605
rect 7837 24565 7849 24599
rect 7883 24596 7895 24599
rect 8202 24596 8208 24608
rect 7883 24568 8208 24596
rect 7883 24565 7895 24568
rect 7837 24559 7895 24565
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 8312 24596 8340 24636
rect 10137 24633 10149 24636
rect 10183 24633 10195 24667
rect 10137 24627 10195 24633
rect 11057 24667 11115 24673
rect 11057 24633 11069 24667
rect 11103 24664 11115 24667
rect 11808 24664 11836 24704
rect 13722 24692 13728 24704
rect 13780 24692 13786 24744
rect 14001 24735 14059 24741
rect 14001 24701 14013 24735
rect 14047 24732 14059 24735
rect 14936 24732 14964 24772
rect 14047 24704 14964 24732
rect 14047 24701 14059 24704
rect 14001 24695 14059 24701
rect 15010 24692 15016 24744
rect 15068 24732 15074 24744
rect 15068 24704 15113 24732
rect 15068 24692 15074 24704
rect 11103 24636 11836 24664
rect 11103 24633 11115 24636
rect 11057 24627 11115 24633
rect 13262 24624 13268 24676
rect 13320 24664 13326 24676
rect 13449 24667 13507 24673
rect 13449 24664 13461 24667
rect 13320 24636 13461 24664
rect 13320 24624 13326 24636
rect 13449 24633 13461 24636
rect 13495 24664 13507 24667
rect 15194 24664 15200 24676
rect 13495 24636 15200 24664
rect 13495 24633 13507 24636
rect 13449 24627 13507 24633
rect 15194 24624 15200 24636
rect 15252 24624 15258 24676
rect 12986 24596 12992 24608
rect 8312 24568 12992 24596
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 15488 24596 15516 24772
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 18509 24803 18567 24809
rect 18509 24800 18521 24803
rect 17920 24772 18521 24800
rect 17920 24760 17926 24772
rect 18509 24769 18521 24772
rect 18555 24769 18567 24803
rect 18509 24763 18567 24769
rect 20272 24772 20668 24800
rect 15654 24732 15660 24744
rect 15615 24704 15660 24732
rect 15654 24692 15660 24704
rect 15712 24692 15718 24744
rect 16298 24732 16304 24744
rect 16259 24704 16304 24732
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 16945 24735 17003 24741
rect 16945 24701 16957 24735
rect 16991 24732 17003 24735
rect 18046 24732 18052 24744
rect 16991 24704 18052 24732
rect 16991 24701 17003 24704
rect 16945 24695 17003 24701
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 18966 24692 18972 24744
rect 19024 24732 19030 24744
rect 19245 24735 19303 24741
rect 19245 24732 19257 24735
rect 19024 24704 19257 24732
rect 19024 24692 19030 24704
rect 19245 24701 19257 24704
rect 19291 24701 19303 24735
rect 19245 24695 19303 24701
rect 19521 24735 19579 24741
rect 19521 24701 19533 24735
rect 19567 24732 19579 24735
rect 20162 24732 20168 24744
rect 19567 24704 20168 24732
rect 19567 24701 19579 24704
rect 19521 24695 19579 24701
rect 15746 24624 15752 24676
rect 15804 24664 15810 24676
rect 19536 24664 19564 24695
rect 20162 24692 20168 24704
rect 20220 24692 20226 24744
rect 20272 24664 20300 24772
rect 20640 24732 20668 24772
rect 21634 24760 21640 24812
rect 21692 24800 21698 24812
rect 22005 24803 22063 24809
rect 22005 24800 22017 24803
rect 21692 24772 22017 24800
rect 21692 24760 21698 24772
rect 22005 24769 22017 24772
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 20640 24704 21496 24732
rect 21358 24664 21364 24676
rect 15804 24636 19564 24664
rect 19628 24636 20300 24664
rect 21319 24636 21364 24664
rect 15804 24624 15810 24636
rect 17494 24596 17500 24608
rect 15488 24568 17500 24596
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 18322 24556 18328 24608
rect 18380 24596 18386 24608
rect 18601 24599 18659 24605
rect 18601 24596 18613 24599
rect 18380 24568 18613 24596
rect 18380 24556 18386 24568
rect 18601 24565 18613 24568
rect 18647 24565 18659 24599
rect 18601 24559 18659 24565
rect 18690 24556 18696 24608
rect 18748 24596 18754 24608
rect 19628 24596 19656 24636
rect 21358 24624 21364 24636
rect 21416 24624 21422 24676
rect 21468 24664 21496 24704
rect 21542 24692 21548 24744
rect 21600 24732 21606 24744
rect 22572 24732 22600 24840
rect 22649 24803 22707 24809
rect 22649 24769 22661 24803
rect 22695 24769 22707 24803
rect 22649 24763 22707 24769
rect 21600 24704 22600 24732
rect 21600 24692 21606 24704
rect 22664 24664 22692 24763
rect 22756 24732 22784 24840
rect 23474 24828 23480 24840
rect 23532 24828 23538 24880
rect 24394 24868 24400 24880
rect 24355 24840 24400 24868
rect 24394 24828 24400 24840
rect 24452 24828 24458 24880
rect 25038 24868 25044 24880
rect 24999 24840 25044 24868
rect 25038 24828 25044 24840
rect 25096 24828 25102 24880
rect 28258 24868 28264 24880
rect 28219 24840 28264 24868
rect 28258 24828 28264 24840
rect 28316 24828 28322 24880
rect 28813 24871 28871 24877
rect 28813 24837 28825 24871
rect 28859 24868 28871 24871
rect 28902 24868 28908 24880
rect 28859 24840 28908 24868
rect 28859 24837 28871 24840
rect 28813 24831 28871 24837
rect 28902 24828 28908 24840
rect 28960 24828 28966 24880
rect 25593 24803 25651 24809
rect 25593 24769 25605 24803
rect 25639 24800 25651 24803
rect 26050 24800 26056 24812
rect 25639 24772 26056 24800
rect 25639 24769 25651 24772
rect 25593 24763 25651 24769
rect 26050 24760 26056 24772
rect 26108 24760 26114 24812
rect 26329 24803 26387 24809
rect 26329 24769 26341 24803
rect 26375 24800 26387 24803
rect 26602 24800 26608 24812
rect 26375 24772 26608 24800
rect 26375 24769 26387 24772
rect 26329 24763 26387 24769
rect 26602 24760 26608 24772
rect 26660 24760 26666 24812
rect 37550 24800 37556 24812
rect 37511 24772 37556 24800
rect 37550 24760 37556 24772
rect 37608 24760 37614 24812
rect 23382 24732 23388 24744
rect 22756 24704 23388 24732
rect 23382 24692 23388 24704
rect 23440 24692 23446 24744
rect 24949 24735 25007 24741
rect 24949 24701 24961 24735
rect 24995 24732 25007 24735
rect 26970 24732 26976 24744
rect 24995 24704 26976 24732
rect 24995 24701 25007 24704
rect 24949 24695 25007 24701
rect 21468 24636 22692 24664
rect 22738 24624 22744 24676
rect 22796 24664 22802 24676
rect 24964 24664 24992 24695
rect 26970 24692 26976 24704
rect 27028 24732 27034 24744
rect 28169 24735 28227 24741
rect 28169 24732 28181 24735
rect 27028 24704 28181 24732
rect 27028 24692 27034 24704
rect 28169 24701 28181 24704
rect 28215 24701 28227 24735
rect 28169 24695 28227 24701
rect 22796 24636 24992 24664
rect 22796 24624 22802 24636
rect 18748 24568 19656 24596
rect 18748 24556 18754 24568
rect 19978 24556 19984 24608
rect 20036 24596 20042 24608
rect 21082 24596 21088 24608
rect 20036 24568 21088 24596
rect 20036 24556 20042 24568
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 21634 24556 21640 24608
rect 21692 24596 21698 24608
rect 22097 24599 22155 24605
rect 22097 24596 22109 24599
rect 21692 24568 22109 24596
rect 21692 24556 21698 24568
rect 22097 24565 22109 24568
rect 22143 24565 22155 24599
rect 22097 24559 22155 24565
rect 22278 24556 22284 24608
rect 22336 24596 22342 24608
rect 24578 24596 24584 24608
rect 22336 24568 24584 24596
rect 22336 24556 22342 24568
rect 24578 24556 24584 24568
rect 24636 24556 24642 24608
rect 37642 24596 37648 24608
rect 37603 24568 37648 24596
rect 37642 24556 37648 24568
rect 37700 24556 37706 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 4065 24395 4123 24401
rect 4065 24361 4077 24395
rect 4111 24392 4123 24395
rect 4706 24392 4712 24404
rect 4111 24364 4712 24392
rect 4111 24361 4123 24364
rect 4065 24355 4123 24361
rect 4706 24352 4712 24364
rect 4764 24352 4770 24404
rect 4890 24352 4896 24404
rect 4948 24392 4954 24404
rect 5902 24392 5908 24404
rect 4948 24364 5908 24392
rect 4948 24352 4954 24364
rect 5902 24352 5908 24364
rect 5960 24352 5966 24404
rect 5994 24352 6000 24404
rect 6052 24392 6058 24404
rect 7742 24392 7748 24404
rect 6052 24364 7748 24392
rect 6052 24352 6058 24364
rect 7742 24352 7748 24364
rect 7800 24352 7806 24404
rect 8573 24395 8631 24401
rect 8573 24361 8585 24395
rect 8619 24392 8631 24395
rect 8662 24392 8668 24404
rect 8619 24364 8668 24392
rect 8619 24361 8631 24364
rect 8573 24355 8631 24361
rect 8662 24352 8668 24364
rect 8720 24352 8726 24404
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9490 24392 9496 24404
rect 9272 24364 9496 24392
rect 9272 24352 9278 24364
rect 9490 24352 9496 24364
rect 9548 24352 9554 24404
rect 9756 24395 9814 24401
rect 9756 24361 9768 24395
rect 9802 24392 9814 24395
rect 13262 24392 13268 24404
rect 9802 24364 13268 24392
rect 9802 24361 9814 24364
rect 9756 24355 9814 24361
rect 13262 24352 13268 24364
rect 13320 24352 13326 24404
rect 14642 24392 14648 24404
rect 14603 24364 14648 24392
rect 14642 24352 14648 24364
rect 14700 24352 14706 24404
rect 15010 24352 15016 24404
rect 15068 24392 15074 24404
rect 15654 24392 15660 24404
rect 15068 24364 15660 24392
rect 15068 24352 15074 24364
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 16117 24395 16175 24401
rect 16117 24361 16129 24395
rect 16163 24392 16175 24395
rect 17034 24392 17040 24404
rect 16163 24364 17040 24392
rect 16163 24361 16175 24364
rect 16117 24355 16175 24361
rect 17034 24352 17040 24364
rect 17092 24352 17098 24404
rect 17770 24352 17776 24404
rect 17828 24392 17834 24404
rect 19978 24392 19984 24404
rect 17828 24364 19984 24392
rect 17828 24352 17834 24364
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 21174 24392 21180 24404
rect 20180 24364 21180 24392
rect 17218 24324 17224 24336
rect 13740 24296 17224 24324
rect 1581 24259 1639 24265
rect 1581 24225 1593 24259
rect 1627 24256 1639 24259
rect 1854 24256 1860 24268
rect 1627 24228 1860 24256
rect 1627 24225 1639 24228
rect 1581 24219 1639 24225
rect 1854 24216 1860 24228
rect 1912 24256 1918 24268
rect 3234 24256 3240 24268
rect 1912 24228 3240 24256
rect 1912 24216 1918 24228
rect 3234 24216 3240 24228
rect 3292 24216 3298 24268
rect 3418 24216 3424 24268
rect 3476 24256 3482 24268
rect 6178 24256 6184 24268
rect 3476 24228 6184 24256
rect 3476 24216 3482 24228
rect 6178 24216 6184 24228
rect 6236 24216 6242 24268
rect 6365 24259 6423 24265
rect 6365 24225 6377 24259
rect 6411 24256 6423 24259
rect 6730 24256 6736 24268
rect 6411 24228 6736 24256
rect 6411 24225 6423 24228
rect 6365 24219 6423 24225
rect 6730 24216 6736 24228
rect 6788 24216 6794 24268
rect 8386 24256 8392 24268
rect 6840 24228 8392 24256
rect 6840 24200 6868 24228
rect 8386 24216 8392 24228
rect 8444 24216 8450 24268
rect 9493 24259 9551 24265
rect 9493 24225 9505 24259
rect 9539 24256 9551 24259
rect 10962 24256 10968 24268
rect 9539 24228 10968 24256
rect 9539 24225 9551 24228
rect 9493 24219 9551 24225
rect 10962 24216 10968 24228
rect 11020 24256 11026 24268
rect 11330 24256 11336 24268
rect 11020 24228 11336 24256
rect 11020 24216 11026 24228
rect 11330 24216 11336 24228
rect 11388 24256 11394 24268
rect 11701 24259 11759 24265
rect 11701 24256 11713 24259
rect 11388 24228 11713 24256
rect 11388 24216 11394 24228
rect 11701 24225 11713 24228
rect 11747 24225 11759 24259
rect 11701 24219 11759 24225
rect 3694 24148 3700 24200
rect 3752 24188 3758 24200
rect 3973 24191 4031 24197
rect 3973 24188 3985 24191
rect 3752 24160 3985 24188
rect 3752 24148 3758 24160
rect 3973 24157 3985 24160
rect 4019 24188 4031 24191
rect 4062 24188 4068 24200
rect 4019 24160 4068 24188
rect 4019 24157 4031 24160
rect 3973 24151 4031 24157
rect 4062 24148 4068 24160
rect 4120 24148 4126 24200
rect 4614 24188 4620 24200
rect 4575 24160 4620 24188
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 6822 24188 6828 24200
rect 6026 24160 6316 24188
rect 6783 24160 6828 24188
rect 1578 24080 1584 24132
rect 1636 24120 1642 24132
rect 1857 24123 1915 24129
rect 1857 24120 1869 24123
rect 1636 24092 1869 24120
rect 1636 24080 1642 24092
rect 1857 24089 1869 24092
rect 1903 24120 1915 24123
rect 3142 24120 3148 24132
rect 1903 24092 2084 24120
rect 3082 24092 3148 24120
rect 1903 24089 1915 24092
rect 1857 24083 1915 24089
rect 2056 24064 2084 24092
rect 3142 24080 3148 24092
rect 3200 24080 3206 24132
rect 4798 24080 4804 24132
rect 4856 24120 4862 24132
rect 4893 24123 4951 24129
rect 4893 24120 4905 24123
rect 4856 24092 4905 24120
rect 4856 24080 4862 24092
rect 4893 24089 4905 24092
rect 4939 24089 4951 24123
rect 4893 24083 4951 24089
rect 2038 24012 2044 24064
rect 2096 24012 2102 24064
rect 2130 24012 2136 24064
rect 2188 24052 2194 24064
rect 3329 24055 3387 24061
rect 3329 24052 3341 24055
rect 2188 24024 3341 24052
rect 2188 24012 2194 24024
rect 3329 24021 3341 24024
rect 3375 24052 3387 24055
rect 5902 24052 5908 24064
rect 3375 24024 5908 24052
rect 3375 24021 3387 24024
rect 3329 24015 3387 24021
rect 5902 24012 5908 24024
rect 5960 24012 5966 24064
rect 6288 24052 6316 24160
rect 6822 24148 6828 24160
rect 6880 24148 6886 24200
rect 13740 24188 13768 24296
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 18874 24284 18880 24336
rect 18932 24324 18938 24336
rect 19242 24324 19248 24336
rect 18932 24296 19248 24324
rect 18932 24284 18938 24296
rect 19242 24284 19248 24296
rect 19300 24284 19306 24336
rect 19702 24324 19708 24336
rect 19663 24296 19708 24324
rect 19702 24284 19708 24296
rect 19760 24284 19766 24336
rect 13814 24216 13820 24268
rect 13872 24256 13878 24268
rect 15473 24259 15531 24265
rect 15473 24256 15485 24259
rect 13872 24228 15485 24256
rect 13872 24216 13878 24228
rect 15473 24225 15485 24228
rect 15519 24225 15531 24259
rect 20180 24256 20208 24364
rect 21174 24352 21180 24364
rect 21232 24352 21238 24404
rect 21266 24352 21272 24404
rect 21324 24392 21330 24404
rect 23198 24392 23204 24404
rect 21324 24364 23204 24392
rect 21324 24352 21330 24364
rect 23198 24352 23204 24364
rect 23256 24352 23262 24404
rect 28169 24395 28227 24401
rect 28169 24361 28181 24395
rect 28215 24392 28227 24395
rect 28258 24392 28264 24404
rect 28215 24364 28264 24392
rect 28215 24361 28227 24364
rect 28169 24355 28227 24361
rect 28258 24352 28264 24364
rect 28316 24352 28322 24404
rect 20530 24324 20536 24336
rect 20272 24296 20536 24324
rect 20272 24265 20300 24296
rect 20530 24284 20536 24296
rect 20588 24324 20594 24336
rect 20990 24324 20996 24336
rect 20588 24296 20996 24324
rect 20588 24284 20594 24296
rect 20990 24284 20996 24296
rect 21048 24284 21054 24336
rect 21542 24284 21548 24336
rect 21600 24324 21606 24336
rect 21910 24324 21916 24336
rect 21600 24296 21916 24324
rect 21600 24284 21606 24296
rect 21910 24284 21916 24296
rect 21968 24284 21974 24336
rect 22370 24284 22376 24336
rect 22428 24324 22434 24336
rect 23753 24327 23811 24333
rect 23753 24324 23765 24327
rect 22428 24296 23765 24324
rect 22428 24284 22434 24296
rect 23753 24293 23765 24296
rect 23799 24293 23811 24327
rect 23753 24287 23811 24293
rect 25866 24284 25872 24336
rect 25924 24324 25930 24336
rect 25924 24296 31754 24324
rect 25924 24284 25930 24296
rect 15473 24219 15531 24225
rect 16040 24228 20208 24256
rect 20257 24259 20315 24265
rect 16040 24197 16068 24228
rect 20257 24225 20269 24259
rect 20303 24225 20315 24259
rect 20714 24256 20720 24268
rect 20675 24228 20720 24256
rect 20257 24219 20315 24225
rect 20714 24216 20720 24228
rect 20772 24216 20778 24268
rect 23382 24216 23388 24268
rect 23440 24256 23446 24268
rect 24673 24259 24731 24265
rect 24673 24256 24685 24259
rect 23440 24228 24685 24256
rect 23440 24216 23446 24228
rect 24673 24225 24685 24228
rect 24719 24225 24731 24259
rect 24673 24219 24731 24225
rect 25317 24259 25375 24265
rect 25317 24225 25329 24259
rect 25363 24256 25375 24259
rect 28902 24256 28908 24268
rect 25363 24228 28908 24256
rect 25363 24225 25375 24228
rect 25317 24219 25375 24225
rect 28902 24216 28908 24228
rect 28960 24216 28966 24268
rect 31726 24256 31754 24296
rect 38378 24256 38384 24268
rect 31726 24228 38384 24256
rect 38378 24216 38384 24228
rect 38436 24216 38442 24268
rect 13110 24160 13768 24188
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24157 15439 24191
rect 15381 24151 15439 24157
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24157 16083 24191
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 16025 24151 16083 24157
rect 7098 24080 7104 24132
rect 7156 24120 7162 24132
rect 10042 24120 10048 24132
rect 7156 24092 7201 24120
rect 8326 24092 10048 24120
rect 7156 24080 7162 24092
rect 10042 24080 10048 24092
rect 10100 24080 10106 24132
rect 10994 24092 11652 24120
rect 7466 24052 7472 24064
rect 6288 24024 7472 24052
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 8754 24012 8760 24064
rect 8812 24052 8818 24064
rect 11054 24052 11060 24064
rect 8812 24024 11060 24052
rect 8812 24012 8818 24024
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 11238 24052 11244 24064
rect 11199 24024 11244 24052
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 11624 24052 11652 24092
rect 11698 24080 11704 24132
rect 11756 24120 11762 24132
rect 11977 24123 12035 24129
rect 11977 24120 11989 24123
rect 11756 24092 11989 24120
rect 11756 24080 11762 24092
rect 11977 24089 11989 24092
rect 12023 24089 12035 24123
rect 11977 24083 12035 24089
rect 12066 24080 12072 24132
rect 12124 24120 12130 24132
rect 12250 24120 12256 24132
rect 12124 24092 12256 24120
rect 12124 24080 12130 24092
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 13262 24080 13268 24132
rect 13320 24120 13326 24132
rect 13725 24123 13783 24129
rect 13725 24120 13737 24123
rect 13320 24092 13737 24120
rect 13320 24080 13326 24092
rect 13725 24089 13737 24092
rect 13771 24089 13783 24123
rect 13998 24120 14004 24132
rect 13725 24083 13783 24089
rect 13825 24092 14004 24120
rect 13825 24052 13853 24092
rect 13998 24080 14004 24092
rect 14056 24080 14062 24132
rect 14553 24123 14611 24129
rect 14553 24089 14565 24123
rect 14599 24120 14611 24123
rect 15102 24120 15108 24132
rect 14599 24092 15108 24120
rect 14599 24089 14611 24092
rect 14553 24083 14611 24089
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 11624 24024 13853 24052
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 15010 24052 15016 24064
rect 13964 24024 15016 24052
rect 13964 24012 13970 24024
rect 15010 24012 15016 24024
rect 15068 24012 15074 24064
rect 15396 24052 15424 24151
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 18785 24191 18843 24197
rect 18785 24157 18797 24191
rect 18831 24188 18843 24191
rect 21818 24188 21824 24200
rect 18831 24160 19656 24188
rect 21779 24160 21824 24188
rect 18831 24157 18843 24160
rect 18785 24151 18843 24157
rect 16758 24120 16764 24132
rect 16719 24092 16764 24120
rect 16758 24080 16764 24092
rect 16816 24080 16822 24132
rect 16853 24123 16911 24129
rect 16853 24089 16865 24123
rect 16899 24120 16911 24123
rect 17586 24120 17592 24132
rect 16899 24092 17592 24120
rect 16899 24089 16911 24092
rect 16853 24083 16911 24089
rect 17586 24080 17592 24092
rect 17644 24080 17650 24132
rect 17770 24120 17776 24132
rect 17731 24092 17776 24120
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 19521 24123 19579 24129
rect 19521 24089 19533 24123
rect 19567 24089 19579 24123
rect 19628 24120 19656 24160
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22094 24148 22100 24200
rect 22152 24188 22158 24200
rect 22370 24188 22376 24200
rect 22152 24160 22376 24188
rect 22152 24148 22158 24160
rect 22370 24148 22376 24160
rect 22428 24148 22434 24200
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24157 22523 24191
rect 22465 24151 22523 24157
rect 26421 24191 26479 24197
rect 26421 24157 26433 24191
rect 26467 24188 26479 24191
rect 28077 24191 28135 24197
rect 28077 24188 28089 24191
rect 26467 24160 28089 24188
rect 26467 24157 26479 24160
rect 26421 24151 26479 24157
rect 28077 24157 28089 24160
rect 28123 24188 28135 24191
rect 28166 24188 28172 24200
rect 28123 24160 28172 24188
rect 28123 24157 28135 24160
rect 28077 24151 28135 24157
rect 20349 24123 20407 24129
rect 20349 24120 20361 24123
rect 19628 24092 20361 24120
rect 19521 24083 19579 24089
rect 20349 24089 20361 24092
rect 20395 24089 20407 24123
rect 20349 24083 20407 24089
rect 17034 24052 17040 24064
rect 15396 24024 17040 24052
rect 17034 24012 17040 24024
rect 17092 24052 17098 24064
rect 17954 24052 17960 24064
rect 17092 24024 17960 24052
rect 17092 24012 17098 24024
rect 17954 24012 17960 24024
rect 18012 24012 18018 24064
rect 18046 24012 18052 24064
rect 18104 24052 18110 24064
rect 19536 24052 19564 24083
rect 20530 24080 20536 24132
rect 20588 24120 20594 24132
rect 22480 24120 22508 24151
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24188 30067 24191
rect 33778 24188 33784 24200
rect 30055 24160 33784 24188
rect 30055 24157 30067 24160
rect 30009 24151 30067 24157
rect 33778 24148 33784 24160
rect 33836 24148 33842 24200
rect 37458 24188 37464 24200
rect 37419 24160 37464 24188
rect 37458 24148 37464 24160
rect 37516 24148 37522 24200
rect 37734 24188 37740 24200
rect 37695 24160 37740 24188
rect 37734 24148 37740 24160
rect 37792 24148 37798 24200
rect 20588 24092 22508 24120
rect 23201 24123 23259 24129
rect 20588 24080 20594 24092
rect 23201 24089 23213 24123
rect 23247 24089 23259 24123
rect 23201 24083 23259 24089
rect 23293 24123 23351 24129
rect 23293 24089 23305 24123
rect 23339 24120 23351 24123
rect 23658 24120 23664 24132
rect 23339 24092 23664 24120
rect 23339 24089 23351 24092
rect 23293 24083 23351 24089
rect 21910 24052 21916 24064
rect 18104 24024 19564 24052
rect 21871 24024 21916 24052
rect 18104 24012 18110 24024
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 22554 24052 22560 24064
rect 22515 24024 22560 24052
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 23216 24052 23244 24083
rect 23658 24080 23664 24092
rect 23716 24080 23722 24132
rect 24765 24123 24823 24129
rect 24765 24089 24777 24123
rect 24811 24120 24823 24123
rect 24946 24120 24952 24132
rect 24811 24092 24952 24120
rect 24811 24089 24823 24092
rect 24765 24083 24823 24089
rect 24946 24080 24952 24092
rect 25004 24080 25010 24132
rect 29270 24120 29276 24132
rect 26436 24092 29276 24120
rect 24670 24052 24676 24064
rect 23216 24024 24676 24052
rect 24670 24012 24676 24024
rect 24728 24052 24734 24064
rect 26436 24052 26464 24092
rect 29270 24080 29276 24092
rect 29328 24120 29334 24132
rect 29328 24092 30144 24120
rect 29328 24080 29334 24092
rect 24728 24024 26464 24052
rect 26513 24055 26571 24061
rect 24728 24012 24734 24024
rect 26513 24021 26525 24055
rect 26559 24052 26571 24055
rect 27338 24052 27344 24064
rect 26559 24024 27344 24052
rect 26559 24021 26571 24024
rect 26513 24015 26571 24021
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 30116 24061 30144 24092
rect 30101 24055 30159 24061
rect 30101 24021 30113 24055
rect 30147 24021 30159 24055
rect 30101 24015 30159 24021
rect 30558 24012 30564 24064
rect 30616 24052 30622 24064
rect 30653 24055 30711 24061
rect 30653 24052 30665 24055
rect 30616 24024 30665 24052
rect 30616 24012 30622 24024
rect 30653 24021 30665 24024
rect 30699 24021 30711 24055
rect 30653 24015 30711 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 2958 23808 2964 23860
rect 3016 23848 3022 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 3016 23820 3617 23848
rect 3016 23808 3022 23820
rect 3605 23817 3617 23820
rect 3651 23848 3663 23851
rect 4062 23848 4068 23860
rect 3651 23820 4068 23848
rect 3651 23817 3663 23820
rect 3605 23811 3663 23817
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 4614 23848 4620 23860
rect 4356 23820 4620 23848
rect 2866 23740 2872 23792
rect 2924 23740 2930 23792
rect 4356 23780 4384 23820
rect 4614 23808 4620 23820
rect 4672 23848 4678 23860
rect 6270 23848 6276 23860
rect 4672 23820 6276 23848
rect 4672 23808 4678 23820
rect 6270 23808 6276 23820
rect 6328 23848 6334 23860
rect 10226 23848 10232 23860
rect 6328 23820 7328 23848
rect 6328 23808 6334 23820
rect 6914 23780 6920 23792
rect 4264 23752 4384 23780
rect 5750 23752 6920 23780
rect 4264 23721 4292 23752
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 7300 23789 7328 23820
rect 7392 23820 10232 23848
rect 7285 23783 7343 23789
rect 7285 23749 7297 23783
rect 7331 23749 7343 23783
rect 7285 23743 7343 23749
rect 4249 23715 4307 23721
rect 4249 23681 4261 23715
rect 4295 23681 4307 23715
rect 4249 23675 4307 23681
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23712 6607 23715
rect 7392 23712 7420 23820
rect 10226 23808 10232 23820
rect 10284 23808 10290 23860
rect 11698 23808 11704 23860
rect 11756 23848 11762 23860
rect 14182 23848 14188 23860
rect 11756 23820 14188 23848
rect 11756 23808 11762 23820
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14366 23808 14372 23860
rect 14424 23848 14430 23860
rect 15194 23848 15200 23860
rect 14424 23820 15200 23848
rect 14424 23808 14430 23820
rect 15194 23808 15200 23820
rect 15252 23808 15258 23860
rect 15286 23808 15292 23860
rect 15344 23848 15350 23860
rect 21818 23848 21824 23860
rect 15344 23820 21824 23848
rect 15344 23808 15350 23820
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 23658 23848 23664 23860
rect 21928 23820 23336 23848
rect 23619 23820 23664 23848
rect 8021 23783 8079 23789
rect 8021 23749 8033 23783
rect 8067 23780 8079 23783
rect 8938 23780 8944 23792
rect 8067 23752 8944 23780
rect 8067 23749 8079 23752
rect 8021 23743 8079 23749
rect 8938 23740 8944 23752
rect 8996 23740 9002 23792
rect 10686 23780 10692 23792
rect 10074 23752 10692 23780
rect 10686 23740 10692 23752
rect 10744 23740 10750 23792
rect 12066 23780 12072 23792
rect 11072 23752 12072 23780
rect 11072 23724 11100 23752
rect 12066 23740 12072 23752
rect 12124 23740 12130 23792
rect 13446 23740 13452 23792
rect 13504 23780 13510 23792
rect 14461 23783 14519 23789
rect 14461 23780 14473 23783
rect 13504 23752 14473 23780
rect 13504 23740 13510 23752
rect 14461 23749 14473 23752
rect 14507 23749 14519 23783
rect 14461 23743 14519 23749
rect 16209 23783 16267 23789
rect 16209 23749 16221 23783
rect 16255 23780 16267 23783
rect 17313 23783 17371 23789
rect 17313 23780 17325 23783
rect 16255 23752 17325 23780
rect 16255 23749 16267 23752
rect 16209 23743 16267 23749
rect 17313 23749 17325 23752
rect 17359 23749 17371 23783
rect 17313 23743 17371 23749
rect 17862 23740 17868 23792
rect 17920 23780 17926 23792
rect 18785 23783 18843 23789
rect 18785 23780 18797 23783
rect 17920 23752 18797 23780
rect 17920 23740 17926 23752
rect 18785 23749 18797 23752
rect 18831 23749 18843 23783
rect 18785 23743 18843 23749
rect 18877 23783 18935 23789
rect 18877 23749 18889 23783
rect 18923 23780 18935 23783
rect 19242 23780 19248 23792
rect 18923 23752 19248 23780
rect 18923 23749 18935 23752
rect 18877 23743 18935 23749
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 19426 23740 19432 23792
rect 19484 23780 19490 23792
rect 19794 23780 19800 23792
rect 19484 23752 19800 23780
rect 19484 23740 19490 23752
rect 19794 23740 19800 23752
rect 19852 23740 19858 23792
rect 19886 23740 19892 23792
rect 19944 23780 19950 23792
rect 20441 23783 20499 23789
rect 20441 23780 20453 23783
rect 19944 23752 20453 23780
rect 19944 23740 19950 23752
rect 20441 23749 20453 23752
rect 20487 23749 20499 23783
rect 20441 23743 20499 23749
rect 20533 23783 20591 23789
rect 20533 23749 20545 23783
rect 20579 23780 20591 23783
rect 21634 23780 21640 23792
rect 20579 23752 21640 23780
rect 20579 23749 20591 23752
rect 20533 23743 20591 23749
rect 21634 23740 21640 23752
rect 21692 23740 21698 23792
rect 6595 23684 7420 23712
rect 6595 23681 6607 23684
rect 6549 23675 6607 23681
rect 1854 23644 1860 23656
rect 1815 23616 1860 23644
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 2133 23647 2191 23653
rect 2133 23613 2145 23647
rect 2179 23644 2191 23647
rect 3418 23644 3424 23656
rect 2179 23616 3424 23644
rect 2179 23613 2191 23616
rect 2133 23607 2191 23613
rect 3418 23604 3424 23616
rect 3476 23604 3482 23656
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23644 4583 23647
rect 5074 23644 5080 23656
rect 4571 23616 5080 23644
rect 4571 23613 4583 23616
rect 4525 23607 4583 23613
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 5258 23604 5264 23656
rect 5316 23644 5322 23656
rect 6564 23644 6592 23675
rect 7926 23672 7932 23724
rect 7984 23712 7990 23724
rect 10597 23715 10655 23721
rect 7984 23684 8029 23712
rect 7984 23672 7990 23684
rect 10597 23681 10609 23715
rect 10643 23712 10655 23715
rect 11054 23712 11060 23724
rect 10643 23684 11060 23712
rect 10643 23681 10655 23684
rect 10597 23675 10655 23681
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 14182 23712 14188 23724
rect 13202 23684 14188 23712
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 16117 23715 16175 23721
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 19720 23684 20300 23712
rect 5316 23616 6592 23644
rect 5316 23604 5322 23616
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 8294 23644 8300 23656
rect 6972 23616 8300 23644
rect 6972 23604 6978 23616
rect 8294 23604 8300 23616
rect 8352 23604 8358 23656
rect 8386 23604 8392 23656
rect 8444 23644 8450 23656
rect 8573 23647 8631 23653
rect 8573 23644 8585 23647
rect 8444 23616 8585 23644
rect 8444 23604 8450 23616
rect 8573 23613 8585 23616
rect 8619 23613 8631 23647
rect 8846 23644 8852 23656
rect 8807 23616 8852 23644
rect 8573 23607 8631 23613
rect 8846 23604 8852 23616
rect 8904 23604 8910 23656
rect 8938 23604 8944 23656
rect 8996 23644 9002 23656
rect 8996 23616 10548 23644
rect 8996 23604 9002 23616
rect 5997 23579 6055 23585
rect 5997 23545 6009 23579
rect 6043 23576 6055 23579
rect 7282 23576 7288 23588
rect 6043 23548 7288 23576
rect 6043 23545 6055 23548
rect 5997 23539 6055 23545
rect 7282 23536 7288 23548
rect 7340 23536 7346 23588
rect 7650 23536 7656 23588
rect 7708 23576 7714 23588
rect 8110 23576 8116 23588
rect 7708 23548 8116 23576
rect 7708 23536 7714 23548
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 10520 23576 10548 23616
rect 10962 23604 10968 23656
rect 11020 23644 11026 23656
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11020 23616 11805 23644
rect 11020 23604 11026 23616
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 12069 23647 12127 23653
rect 12069 23644 12081 23647
rect 11793 23607 11851 23613
rect 11900 23616 12081 23644
rect 11422 23576 11428 23588
rect 10520 23548 11428 23576
rect 11422 23536 11428 23548
rect 11480 23536 11486 23588
rect 11514 23536 11520 23588
rect 11572 23576 11578 23588
rect 11900 23576 11928 23616
rect 12069 23613 12081 23616
rect 12115 23644 12127 23647
rect 12158 23644 12164 23656
rect 12115 23616 12164 23644
rect 12115 23613 12127 23616
rect 12069 23607 12127 23613
rect 12158 23604 12164 23616
rect 12216 23604 12222 23656
rect 12618 23604 12624 23656
rect 12676 23644 12682 23656
rect 13814 23644 13820 23656
rect 12676 23616 13124 23644
rect 13775 23616 13820 23644
rect 12676 23604 12682 23616
rect 11572 23548 11928 23576
rect 13096 23576 13124 23616
rect 13814 23604 13820 23616
rect 13872 23604 13878 23656
rect 14366 23644 14372 23656
rect 14327 23616 14372 23644
rect 14366 23604 14372 23616
rect 14424 23604 14430 23656
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 14645 23647 14703 23653
rect 14645 23644 14657 23647
rect 14608 23616 14657 23644
rect 14608 23604 14614 23616
rect 14645 23613 14657 23616
rect 14691 23613 14703 23647
rect 14645 23607 14703 23613
rect 13446 23576 13452 23588
rect 13096 23548 13452 23576
rect 11572 23536 11578 23548
rect 13446 23536 13452 23548
rect 13504 23576 13510 23588
rect 16022 23576 16028 23588
rect 13504 23548 16028 23576
rect 13504 23536 13510 23548
rect 16022 23536 16028 23548
rect 16080 23536 16086 23588
rect 2222 23468 2228 23520
rect 2280 23508 2286 23520
rect 5626 23508 5632 23520
rect 2280 23480 5632 23508
rect 2280 23468 2286 23480
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 6730 23468 6736 23520
rect 6788 23508 6794 23520
rect 7098 23508 7104 23520
rect 6788 23480 7104 23508
rect 6788 23468 6794 23480
rect 7098 23468 7104 23480
rect 7156 23468 7162 23520
rect 7190 23468 7196 23520
rect 7248 23508 7254 23520
rect 7742 23508 7748 23520
rect 7248 23480 7748 23508
rect 7248 23468 7254 23480
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 9490 23468 9496 23520
rect 9548 23508 9554 23520
rect 16132 23508 16160 23675
rect 17218 23644 17224 23656
rect 17179 23616 17224 23644
rect 17218 23604 17224 23616
rect 17276 23604 17282 23656
rect 17494 23644 17500 23656
rect 17455 23616 17500 23644
rect 17494 23604 17500 23616
rect 17552 23644 17558 23656
rect 19720 23644 19748 23684
rect 17552 23616 19748 23644
rect 17552 23604 17558 23616
rect 19794 23604 19800 23656
rect 19852 23644 19858 23656
rect 20272 23644 20300 23684
rect 20898 23644 20904 23656
rect 19852 23616 20208 23644
rect 20272 23616 20904 23644
rect 19852 23604 19858 23616
rect 16758 23536 16764 23588
rect 16816 23576 16822 23588
rect 17862 23576 17868 23588
rect 16816 23548 17868 23576
rect 16816 23536 16822 23548
rect 17862 23536 17868 23548
rect 17920 23536 17926 23588
rect 17954 23536 17960 23588
rect 18012 23576 18018 23588
rect 19426 23576 19432 23588
rect 18012 23548 19432 23576
rect 18012 23536 18018 23548
rect 19426 23536 19432 23548
rect 19484 23536 19490 23588
rect 20180 23576 20208 23616
rect 20898 23604 20904 23616
rect 20956 23604 20962 23656
rect 21082 23644 21088 23656
rect 21043 23616 21088 23644
rect 21082 23604 21088 23616
rect 21140 23644 21146 23656
rect 21928 23644 21956 23820
rect 22189 23783 22247 23789
rect 22189 23749 22201 23783
rect 22235 23780 22247 23783
rect 22278 23780 22284 23792
rect 22235 23752 22284 23780
rect 22235 23749 22247 23752
rect 22189 23743 22247 23749
rect 22278 23740 22284 23752
rect 22336 23740 22342 23792
rect 23109 23783 23167 23789
rect 23109 23749 23121 23783
rect 23155 23780 23167 23783
rect 23198 23780 23204 23792
rect 23155 23752 23204 23780
rect 23155 23749 23167 23752
rect 23109 23743 23167 23749
rect 23198 23740 23204 23752
rect 23256 23740 23262 23792
rect 23308 23780 23336 23820
rect 23658 23808 23664 23820
rect 23716 23808 23722 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 25280 23820 29868 23848
rect 25280 23808 25286 23820
rect 23934 23780 23940 23792
rect 23308 23752 23940 23780
rect 23934 23740 23940 23752
rect 23992 23740 23998 23792
rect 27338 23780 27344 23792
rect 24228 23752 25084 23780
rect 27299 23752 27344 23780
rect 23566 23712 23572 23724
rect 23527 23684 23572 23712
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 24228 23721 24256 23752
rect 25056 23724 25084 23752
rect 27338 23740 27344 23752
rect 27396 23740 27402 23792
rect 28626 23780 28632 23792
rect 28587 23752 28632 23780
rect 28626 23740 28632 23752
rect 28684 23740 28690 23792
rect 24213 23715 24271 23721
rect 24213 23681 24225 23715
rect 24259 23681 24271 23715
rect 24213 23675 24271 23681
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 24857 23715 24915 23721
rect 24857 23712 24869 23715
rect 24544 23684 24869 23712
rect 24544 23672 24550 23684
rect 24857 23681 24869 23684
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 21140 23616 21956 23644
rect 22097 23647 22155 23653
rect 21140 23604 21146 23616
rect 22097 23613 22109 23647
rect 22143 23644 22155 23647
rect 22738 23644 22744 23656
rect 22143 23616 22744 23644
rect 22143 23613 22155 23616
rect 22097 23607 22155 23613
rect 22738 23604 22744 23616
rect 22796 23604 22802 23656
rect 22370 23576 22376 23588
rect 20180 23548 22376 23576
rect 22370 23536 22376 23548
rect 22428 23536 22434 23588
rect 24872 23576 24900 23675
rect 25038 23672 25044 23724
rect 25096 23712 25102 23724
rect 25501 23715 25559 23721
rect 25501 23712 25513 23715
rect 25096 23684 25513 23712
rect 25096 23672 25102 23684
rect 25501 23681 25513 23684
rect 25547 23681 25559 23715
rect 25501 23675 25559 23681
rect 26145 23715 26203 23721
rect 26145 23681 26157 23715
rect 26191 23712 26203 23715
rect 26602 23712 26608 23724
rect 26191 23684 26608 23712
rect 26191 23681 26203 23684
rect 26145 23675 26203 23681
rect 26602 23672 26608 23684
rect 26660 23672 26666 23724
rect 29840 23721 29868 23820
rect 30558 23780 30564 23792
rect 30519 23752 30564 23780
rect 30558 23740 30564 23752
rect 30616 23740 30622 23792
rect 30653 23783 30711 23789
rect 30653 23749 30665 23783
rect 30699 23780 30711 23783
rect 30742 23780 30748 23792
rect 30699 23752 30748 23780
rect 30699 23749 30711 23752
rect 30653 23743 30711 23749
rect 30742 23740 30748 23752
rect 30800 23740 30806 23792
rect 29825 23715 29883 23721
rect 29825 23681 29837 23715
rect 29871 23681 29883 23715
rect 29825 23675 29883 23681
rect 26510 23604 26516 23656
rect 26568 23644 26574 23656
rect 27246 23644 27252 23656
rect 26568 23616 27252 23644
rect 26568 23604 26574 23616
rect 27246 23604 27252 23616
rect 27304 23604 27310 23656
rect 27890 23644 27896 23656
rect 27851 23616 27896 23644
rect 27890 23604 27896 23616
rect 27948 23604 27954 23656
rect 28537 23647 28595 23653
rect 28537 23613 28549 23647
rect 28583 23644 28595 23647
rect 28902 23644 28908 23656
rect 28583 23616 28908 23644
rect 28583 23613 28595 23616
rect 28537 23607 28595 23613
rect 28902 23604 28908 23616
rect 28960 23604 28966 23656
rect 29181 23647 29239 23653
rect 29181 23613 29193 23647
rect 29227 23644 29239 23647
rect 30650 23644 30656 23656
rect 29227 23616 30656 23644
rect 29227 23613 29239 23616
rect 29181 23607 29239 23613
rect 30650 23604 30656 23616
rect 30708 23644 30714 23656
rect 30834 23644 30840 23656
rect 30708 23616 30840 23644
rect 30708 23604 30714 23616
rect 30834 23604 30840 23616
rect 30892 23604 30898 23656
rect 29730 23576 29736 23588
rect 24872 23548 29736 23576
rect 29730 23536 29736 23548
rect 29788 23536 29794 23588
rect 9548 23480 16160 23508
rect 9548 23468 9554 23480
rect 16390 23468 16396 23520
rect 16448 23508 16454 23520
rect 21266 23508 21272 23520
rect 16448 23480 21272 23508
rect 16448 23468 16454 23480
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 23658 23468 23664 23520
rect 23716 23508 23722 23520
rect 24305 23511 24363 23517
rect 24305 23508 24317 23511
rect 23716 23480 24317 23508
rect 23716 23468 23722 23480
rect 24305 23477 24317 23480
rect 24351 23477 24363 23511
rect 24305 23471 24363 23477
rect 24946 23468 24952 23520
rect 25004 23508 25010 23520
rect 25593 23511 25651 23517
rect 25593 23508 25605 23511
rect 25004 23480 25605 23508
rect 25004 23468 25010 23480
rect 25593 23477 25605 23480
rect 25639 23477 25651 23511
rect 26234 23508 26240 23520
rect 26195 23480 26240 23508
rect 25593 23471 25651 23477
rect 26234 23468 26240 23480
rect 26292 23468 26298 23520
rect 29641 23511 29699 23517
rect 29641 23477 29653 23511
rect 29687 23508 29699 23511
rect 36078 23508 36084 23520
rect 29687 23480 36084 23508
rect 29687 23477 29699 23480
rect 29641 23471 29699 23477
rect 36078 23468 36084 23480
rect 36136 23468 36142 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 2222 23264 2228 23316
rect 2280 23304 2286 23316
rect 2406 23304 2412 23316
rect 2280 23276 2412 23304
rect 2280 23264 2286 23276
rect 2406 23264 2412 23276
rect 2464 23264 2470 23316
rect 5721 23307 5779 23313
rect 5721 23304 5733 23307
rect 3896 23276 5733 23304
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 1854 23168 1860 23180
rect 1627 23140 1860 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 1854 23128 1860 23140
rect 1912 23128 1918 23180
rect 1946 23128 1952 23180
rect 2004 23168 2010 23180
rect 2406 23168 2412 23180
rect 2004 23140 2412 23168
rect 2004 23128 2010 23140
rect 2406 23128 2412 23140
rect 2464 23168 2470 23180
rect 3896 23168 3924 23276
rect 5721 23273 5733 23276
rect 5767 23273 5779 23307
rect 5721 23267 5779 23273
rect 5810 23264 5816 23316
rect 5868 23304 5874 23316
rect 20806 23304 20812 23316
rect 5868 23276 10640 23304
rect 5868 23264 5874 23276
rect 8570 23236 8576 23248
rect 7944 23208 8576 23236
rect 2464 23140 3924 23168
rect 3973 23171 4031 23177
rect 2464 23128 2470 23140
rect 3973 23137 3985 23171
rect 4019 23168 4031 23171
rect 4246 23168 4252 23180
rect 4019 23140 4252 23168
rect 4019 23137 4031 23140
rect 3973 23131 4031 23137
rect 4246 23128 4252 23140
rect 4304 23168 4310 23180
rect 4614 23168 4620 23180
rect 4304 23140 4620 23168
rect 4304 23128 4310 23140
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 5442 23168 5448 23180
rect 5368 23140 5448 23168
rect 5368 23086 5396 23140
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 6825 23171 6883 23177
rect 6825 23137 6837 23171
rect 6871 23168 6883 23171
rect 7944 23168 7972 23208
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 8662 23196 8668 23248
rect 8720 23236 8726 23248
rect 8938 23236 8944 23248
rect 8720 23208 8944 23236
rect 8720 23196 8726 23208
rect 8938 23196 8944 23208
rect 8996 23196 9002 23248
rect 10612 23236 10640 23276
rect 11716 23276 20812 23304
rect 11716 23236 11744 23276
rect 10612 23208 11744 23236
rect 6871 23140 7972 23168
rect 6871 23137 6883 23140
rect 6825 23131 6883 23137
rect 8018 23128 8024 23180
rect 8076 23128 8082 23180
rect 8386 23128 8392 23180
rect 8444 23128 8450 23180
rect 9585 23171 9643 23177
rect 9585 23137 9597 23171
rect 9631 23168 9643 23171
rect 11238 23168 11244 23180
rect 9631 23140 11244 23168
rect 9631 23137 9643 23140
rect 9585 23131 9643 23137
rect 11238 23128 11244 23140
rect 11296 23128 11302 23180
rect 11330 23128 11336 23180
rect 11388 23168 11394 23180
rect 11974 23168 11980 23180
rect 11388 23140 11980 23168
rect 11388 23128 11394 23140
rect 11974 23128 11980 23140
rect 12032 23128 12038 23180
rect 12066 23128 12072 23180
rect 12124 23168 12130 23180
rect 13262 23168 13268 23180
rect 12124 23140 13268 23168
rect 12124 23128 12130 23140
rect 13262 23128 13268 23140
rect 13320 23128 13326 23180
rect 13740 23177 13768 23276
rect 20806 23264 20812 23276
rect 20864 23304 20870 23316
rect 23382 23304 23388 23316
rect 20864 23276 23388 23304
rect 20864 23264 20870 23276
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 23477 23307 23535 23313
rect 23477 23273 23489 23307
rect 23523 23304 23535 23307
rect 30558 23304 30564 23316
rect 23523 23276 30564 23304
rect 23523 23273 23535 23276
rect 23477 23267 23535 23273
rect 30558 23264 30564 23276
rect 30616 23264 30622 23316
rect 14366 23196 14372 23248
rect 14424 23236 14430 23248
rect 14826 23236 14832 23248
rect 14424 23208 14832 23236
rect 14424 23196 14430 23208
rect 14826 23196 14832 23208
rect 14884 23196 14890 23248
rect 15470 23196 15476 23248
rect 15528 23236 15534 23248
rect 15933 23239 15991 23245
rect 15933 23236 15945 23239
rect 15528 23208 15945 23236
rect 15528 23196 15534 23208
rect 15933 23205 15945 23208
rect 15979 23205 15991 23239
rect 15933 23199 15991 23205
rect 16850 23196 16856 23248
rect 16908 23236 16914 23248
rect 21450 23236 21456 23248
rect 16908 23208 17448 23236
rect 16908 23196 16914 23208
rect 17420 23180 17448 23208
rect 18064 23208 21456 23236
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23137 13783 23171
rect 17218 23168 17224 23180
rect 13725 23131 13783 23137
rect 14200 23140 17224 23168
rect 6549 23103 6607 23109
rect 6549 23069 6561 23103
rect 6595 23069 6607 23103
rect 8036 23100 8064 23128
rect 7958 23072 8064 23100
rect 8404 23100 8432 23128
rect 9306 23100 9312 23112
rect 8404 23072 9312 23100
rect 6549 23063 6607 23069
rect 1762 22992 1768 23044
rect 1820 23032 1826 23044
rect 1857 23035 1915 23041
rect 1857 23032 1869 23035
rect 1820 23004 1869 23032
rect 1820 22992 1826 23004
rect 1857 23001 1869 23004
rect 1903 23001 1915 23035
rect 3602 23032 3608 23044
rect 3082 23004 3608 23032
rect 1857 22995 1915 23001
rect 3602 22992 3608 23004
rect 3660 22992 3666 23044
rect 4249 23035 4307 23041
rect 4249 23001 4261 23035
rect 4295 23001 4307 23035
rect 6564 23032 6592 23063
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 10962 23060 10968 23112
rect 11020 23100 11026 23112
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 11020 23072 11713 23100
rect 11020 23060 11026 23072
rect 11701 23069 11713 23072
rect 11747 23069 11759 23103
rect 13280 23100 13308 23128
rect 14200 23100 14228 23140
rect 17218 23128 17224 23140
rect 17276 23128 17282 23180
rect 17402 23168 17408 23180
rect 17363 23140 17408 23168
rect 17402 23128 17408 23140
rect 17460 23128 17466 23180
rect 15841 23103 15899 23109
rect 15841 23100 15853 23103
rect 13280 23072 14228 23100
rect 15212 23072 15853 23100
rect 11701 23063 11759 23069
rect 6914 23032 6920 23044
rect 6564 23004 6920 23032
rect 4249 22995 4307 23001
rect 3326 22964 3332 22976
rect 3287 22936 3332 22964
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 4264 22964 4292 22995
rect 6914 22992 6920 23004
rect 6972 22992 6978 23044
rect 8386 22992 8392 23044
rect 8444 23032 8450 23044
rect 8573 23035 8631 23041
rect 8573 23032 8585 23035
rect 8444 23004 8585 23032
rect 8444 22992 8450 23004
rect 8573 23001 8585 23004
rect 8619 23032 8631 23035
rect 11238 23032 11244 23044
rect 8619 23004 9812 23032
rect 10810 23004 11244 23032
rect 8619 23001 8631 23004
rect 8573 22995 8631 23001
rect 9784 22976 9812 23004
rect 11238 22992 11244 23004
rect 11296 22992 11302 23044
rect 11977 23035 12035 23041
rect 11977 23001 11989 23035
rect 12023 23032 12035 23035
rect 12250 23032 12256 23044
rect 12023 23004 12256 23032
rect 12023 23001 12035 23004
rect 11977 22995 12035 23001
rect 12250 22992 12256 23004
rect 12308 22992 12314 23044
rect 13630 23032 13636 23044
rect 13202 23004 13636 23032
rect 13630 22992 13636 23004
rect 13688 22992 13694 23044
rect 14090 22992 14096 23044
rect 14148 23032 14154 23044
rect 14369 23035 14427 23041
rect 14369 23032 14381 23035
rect 14148 23004 14381 23032
rect 14148 22992 14154 23004
rect 14369 23001 14381 23004
rect 14415 23001 14427 23035
rect 14369 22995 14427 23001
rect 14458 22992 14464 23044
rect 14516 23032 14522 23044
rect 14516 23004 14561 23032
rect 14516 22992 14522 23004
rect 15010 22992 15016 23044
rect 15068 23032 15074 23044
rect 15212 23032 15240 23072
rect 15841 23069 15853 23072
rect 15887 23100 15899 23103
rect 15887 23072 16436 23100
rect 15887 23069 15899 23072
rect 15841 23063 15899 23069
rect 15068 23004 15240 23032
rect 15381 23035 15439 23041
rect 15068 22992 15074 23004
rect 15381 23001 15393 23035
rect 15427 23032 15439 23035
rect 16206 23032 16212 23044
rect 15427 23004 16212 23032
rect 15427 23001 15439 23004
rect 15381 22995 15439 23001
rect 16206 22992 16212 23004
rect 16264 22992 16270 23044
rect 16408 23032 16436 23072
rect 16577 23035 16635 23041
rect 16408 23004 16528 23032
rect 16500 22976 16528 23004
rect 16577 23001 16589 23035
rect 16623 23001 16635 23035
rect 16577 22995 16635 23001
rect 6546 22964 6552 22976
rect 4264 22936 6552 22964
rect 6546 22924 6552 22936
rect 6604 22924 6610 22976
rect 9766 22924 9772 22976
rect 9824 22924 9830 22976
rect 11057 22967 11115 22973
rect 11057 22933 11069 22967
rect 11103 22964 11115 22967
rect 11606 22964 11612 22976
rect 11103 22936 11612 22964
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 11606 22924 11612 22936
rect 11664 22964 11670 22976
rect 15194 22964 15200 22976
rect 11664 22936 15200 22964
rect 11664 22924 11670 22936
rect 15194 22924 15200 22936
rect 15252 22924 15258 22976
rect 16482 22924 16488 22976
rect 16540 22924 16546 22976
rect 16592 22964 16620 22995
rect 16666 22992 16672 23044
rect 16724 23032 16730 23044
rect 16724 23004 16769 23032
rect 16724 22992 16730 23004
rect 18064 22964 18092 23208
rect 21450 23196 21456 23208
rect 21508 23196 21514 23248
rect 21542 23196 21548 23248
rect 21600 23236 21606 23248
rect 28534 23236 28540 23248
rect 21600 23208 24992 23236
rect 21600 23196 21606 23208
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23168 18291 23171
rect 19886 23168 19892 23180
rect 18279 23140 19892 23168
rect 18279 23137 18291 23140
rect 18233 23131 18291 23137
rect 19886 23128 19892 23140
rect 19944 23168 19950 23180
rect 20346 23168 20352 23180
rect 19944 23140 20352 23168
rect 19944 23128 19950 23140
rect 20346 23128 20352 23140
rect 20404 23128 20410 23180
rect 22002 23128 22008 23180
rect 22060 23168 22066 23180
rect 24670 23168 24676 23180
rect 22060 23140 23428 23168
rect 24631 23140 24676 23168
rect 22060 23128 22066 23140
rect 23400 23109 23428 23140
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 24964 23177 24992 23208
rect 27816 23208 28540 23236
rect 24949 23171 25007 23177
rect 24949 23137 24961 23171
rect 24995 23137 25007 23171
rect 24949 23131 25007 23137
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 27816 23168 27844 23208
rect 28534 23196 28540 23208
rect 28592 23196 28598 23248
rect 26835 23140 27844 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 27890 23128 27896 23180
rect 27948 23168 27954 23180
rect 28626 23168 28632 23180
rect 27948 23140 28632 23168
rect 27948 23128 27954 23140
rect 28626 23128 28632 23140
rect 28684 23128 28690 23180
rect 23385 23103 23443 23109
rect 23385 23069 23397 23103
rect 23431 23069 23443 23103
rect 29730 23100 29736 23112
rect 29691 23072 29736 23100
rect 23385 23063 23443 23069
rect 29730 23060 29736 23072
rect 29788 23100 29794 23112
rect 30282 23100 30288 23112
rect 29788 23072 30288 23100
rect 29788 23060 29794 23072
rect 30282 23060 30288 23072
rect 30340 23060 30346 23112
rect 18322 22992 18328 23044
rect 18380 23032 18386 23044
rect 18874 23032 18880 23044
rect 18380 23004 18425 23032
rect 18835 23004 18880 23032
rect 18380 22992 18386 23004
rect 18874 22992 18880 23004
rect 18932 22992 18938 23044
rect 19981 23035 20039 23041
rect 19981 23001 19993 23035
rect 20027 23001 20039 23035
rect 20898 23032 20904 23044
rect 20859 23004 20904 23032
rect 19981 22995 20039 23001
rect 16592 22936 18092 22964
rect 19996 22964 20024 22995
rect 20898 22992 20904 23004
rect 20956 23032 20962 23044
rect 21542 23032 21548 23044
rect 20956 23004 21548 23032
rect 20956 22992 20962 23004
rect 21542 22992 21548 23004
rect 21600 22992 21606 23044
rect 21910 23032 21916 23044
rect 21871 23004 21916 23032
rect 21910 22992 21916 23004
rect 21968 22992 21974 23044
rect 22005 23035 22063 23041
rect 22005 23001 22017 23035
rect 22051 23032 22063 23035
rect 22554 23032 22560 23044
rect 22051 23004 22560 23032
rect 22051 23001 22063 23004
rect 22005 22995 22063 23001
rect 22554 22992 22560 23004
rect 22612 22992 22618 23044
rect 22738 22992 22744 23044
rect 22796 23032 22802 23044
rect 22925 23035 22983 23041
rect 22925 23032 22937 23035
rect 22796 23004 22937 23032
rect 22796 22992 22802 23004
rect 22925 23001 22937 23004
rect 22971 23001 22983 23035
rect 23566 23032 23572 23044
rect 22925 22995 22983 23001
rect 23032 23004 23572 23032
rect 23032 22964 23060 23004
rect 23566 22992 23572 23004
rect 23624 22992 23630 23044
rect 24765 23035 24823 23041
rect 24765 23001 24777 23035
rect 24811 23032 24823 23035
rect 24946 23032 24952 23044
rect 24811 23004 24952 23032
rect 24811 23001 24823 23004
rect 24765 22995 24823 23001
rect 24946 22992 24952 23004
rect 25004 22992 25010 23044
rect 25498 22992 25504 23044
rect 25556 23032 25562 23044
rect 26881 23035 26939 23041
rect 26881 23032 26893 23035
rect 25556 23004 26893 23032
rect 25556 22992 25562 23004
rect 26881 23001 26893 23004
rect 26927 23001 26939 23035
rect 26881 22995 26939 23001
rect 27801 23035 27859 23041
rect 27801 23001 27813 23035
rect 27847 23032 27859 23035
rect 27982 23032 27988 23044
rect 27847 23004 27988 23032
rect 27847 23001 27859 23004
rect 27801 22995 27859 23001
rect 27982 22992 27988 23004
rect 28040 22992 28046 23044
rect 28350 23032 28356 23044
rect 28311 23004 28356 23032
rect 28350 22992 28356 23004
rect 28408 22992 28414 23044
rect 28445 23035 28503 23041
rect 28445 23001 28457 23035
rect 28491 23001 28503 23035
rect 28445 22995 28503 23001
rect 19996 22936 23060 22964
rect 28460 22964 28488 22995
rect 29825 22967 29883 22973
rect 29825 22964 29837 22967
rect 28460 22936 29837 22964
rect 29825 22933 29837 22936
rect 29871 22933 29883 22967
rect 29825 22927 29883 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1670 22720 1676 22772
rect 1728 22760 1734 22772
rect 4154 22760 4160 22772
rect 1728 22732 4160 22760
rect 1728 22720 1734 22732
rect 4154 22720 4160 22732
rect 4212 22720 4218 22772
rect 5718 22720 5724 22772
rect 5776 22760 5782 22772
rect 5905 22763 5963 22769
rect 5905 22760 5917 22763
rect 5776 22732 5917 22760
rect 5776 22720 5782 22732
rect 5905 22729 5917 22732
rect 5951 22760 5963 22763
rect 6454 22760 6460 22772
rect 5951 22732 6460 22760
rect 5951 22729 5963 22732
rect 5905 22723 5963 22729
rect 6454 22720 6460 22732
rect 6512 22720 6518 22772
rect 10962 22760 10968 22772
rect 7668 22732 10968 22760
rect 1302 22652 1308 22704
rect 1360 22692 1366 22704
rect 1360 22664 2622 22692
rect 1360 22652 1366 22664
rect 3510 22652 3516 22704
rect 3568 22692 3574 22704
rect 4433 22695 4491 22701
rect 4433 22692 4445 22695
rect 3568 22664 4445 22692
rect 3568 22652 3574 22664
rect 4433 22661 4445 22664
rect 4479 22692 4491 22695
rect 4522 22692 4528 22704
rect 4479 22664 4528 22692
rect 4479 22661 4491 22664
rect 4433 22655 4491 22661
rect 4522 22652 4528 22664
rect 4580 22652 4586 22704
rect 6638 22652 6644 22704
rect 6696 22692 6702 22704
rect 6733 22695 6791 22701
rect 6733 22692 6745 22695
rect 6696 22664 6745 22692
rect 6696 22652 6702 22664
rect 6733 22661 6745 22664
rect 6779 22661 6791 22695
rect 6733 22655 6791 22661
rect 4154 22624 4160 22636
rect 4115 22596 4160 22624
rect 4154 22584 4160 22596
rect 4212 22584 4218 22636
rect 5534 22584 5540 22636
rect 5592 22584 5598 22636
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 7668 22624 7696 22732
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 11238 22720 11244 22772
rect 11296 22760 11302 22772
rect 12434 22760 12440 22772
rect 11296 22732 12440 22760
rect 11296 22720 11302 22732
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 12802 22720 12808 22772
rect 12860 22760 12866 22772
rect 13998 22760 14004 22772
rect 12860 22732 14004 22760
rect 12860 22720 12866 22732
rect 13998 22720 14004 22732
rect 14056 22720 14062 22772
rect 17678 22760 17684 22772
rect 14108 22732 17684 22760
rect 9582 22692 9588 22704
rect 9246 22664 9588 22692
rect 9582 22652 9588 22664
rect 9640 22652 9646 22704
rect 9766 22652 9772 22704
rect 9824 22692 9830 22704
rect 10042 22692 10048 22704
rect 9824 22664 10048 22692
rect 9824 22652 9830 22664
rect 10042 22652 10048 22664
rect 10100 22652 10106 22704
rect 12161 22695 12219 22701
rect 12161 22661 12173 22695
rect 12207 22692 12219 22695
rect 12250 22692 12256 22704
rect 12207 22664 12256 22692
rect 12207 22661 12219 22664
rect 12161 22655 12219 22661
rect 12250 22652 12256 22664
rect 12308 22652 12314 22704
rect 12618 22652 12624 22704
rect 12676 22652 12682 22704
rect 13538 22652 13544 22704
rect 13596 22692 13602 22704
rect 14108 22692 14136 22732
rect 17678 22720 17684 22732
rect 17736 22720 17742 22772
rect 18874 22760 18880 22772
rect 17788 22732 18880 22760
rect 14274 22692 14280 22704
rect 13596 22664 14136 22692
rect 14235 22664 14280 22692
rect 13596 22652 13602 22664
rect 14274 22652 14280 22664
rect 14332 22652 14338 22704
rect 14642 22652 14648 22704
rect 14700 22692 14706 22704
rect 15930 22692 15936 22704
rect 14700 22664 15936 22692
rect 14700 22652 14706 22664
rect 15930 22652 15936 22664
rect 15988 22652 15994 22704
rect 16209 22695 16267 22701
rect 16209 22661 16221 22695
rect 16255 22692 16267 22695
rect 17037 22695 17095 22701
rect 17037 22692 17049 22695
rect 16255 22664 17049 22692
rect 16255 22661 16267 22664
rect 16209 22655 16267 22661
rect 17037 22661 17049 22664
rect 17083 22661 17095 22695
rect 17037 22655 17095 22661
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 7340 22596 7385 22624
rect 7668 22596 7757 22624
rect 7340 22584 7346 22596
rect 7745 22593 7757 22596
rect 7791 22593 7803 22627
rect 7745 22587 7803 22593
rect 9306 22584 9312 22636
rect 9364 22624 9370 22636
rect 9950 22624 9956 22636
rect 9364 22596 9956 22624
rect 9364 22584 9370 22596
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 10226 22624 10232 22636
rect 10187 22596 10232 22624
rect 10226 22584 10232 22596
rect 10284 22584 10290 22636
rect 15286 22584 15292 22636
rect 15344 22624 15350 22636
rect 15746 22624 15752 22636
rect 15344 22596 15752 22624
rect 15344 22584 15350 22596
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 16117 22627 16175 22633
rect 16117 22593 16129 22627
rect 16163 22624 16175 22627
rect 16666 22624 16672 22636
rect 16163 22596 16672 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 16758 22584 16764 22636
rect 16816 22584 16822 22636
rect 1670 22516 1676 22568
rect 1728 22556 1734 22568
rect 1857 22559 1915 22565
rect 1857 22556 1869 22559
rect 1728 22528 1869 22556
rect 1728 22516 1734 22528
rect 1857 22525 1869 22528
rect 1903 22525 1915 22559
rect 2130 22556 2136 22568
rect 2091 22528 2136 22556
rect 1857 22519 1915 22525
rect 2130 22516 2136 22528
rect 2188 22516 2194 22568
rect 2774 22516 2780 22568
rect 2832 22556 2838 22568
rect 6641 22559 6699 22565
rect 2832 22528 3280 22556
rect 2832 22516 2838 22528
rect 3252 22500 3280 22528
rect 6641 22525 6653 22559
rect 6687 22556 6699 22559
rect 7374 22556 7380 22568
rect 6687 22528 7380 22556
rect 6687 22525 6699 22528
rect 6641 22519 6699 22525
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 8018 22556 8024 22568
rect 7979 22528 8024 22556
rect 8018 22516 8024 22528
rect 8076 22516 8082 22568
rect 8570 22516 8576 22568
rect 8628 22556 8634 22568
rect 9214 22556 9220 22568
rect 8628 22528 9220 22556
rect 8628 22516 8634 22528
rect 9214 22516 9220 22528
rect 9272 22556 9278 22568
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9272 22528 9781 22556
rect 9272 22516 9278 22528
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 10962 22556 10968 22568
rect 10923 22528 10968 22556
rect 9769 22519 9827 22525
rect 10962 22516 10968 22528
rect 11020 22556 11026 22568
rect 11885 22559 11943 22565
rect 11885 22556 11897 22559
rect 11020 22528 11897 22556
rect 11020 22516 11026 22528
rect 11885 22525 11897 22528
rect 11931 22525 11943 22559
rect 13170 22556 13176 22568
rect 11885 22519 11943 22525
rect 11992 22528 13176 22556
rect 3234 22448 3240 22500
rect 3292 22488 3298 22500
rect 3605 22491 3663 22497
rect 3605 22488 3617 22491
rect 3292 22460 3617 22488
rect 3292 22448 3298 22460
rect 3605 22457 3617 22460
rect 3651 22457 3663 22491
rect 3605 22451 3663 22457
rect 5534 22448 5540 22500
rect 5592 22488 5598 22500
rect 7466 22488 7472 22500
rect 5592 22460 7472 22488
rect 5592 22448 5598 22460
rect 7466 22448 7472 22460
rect 7524 22448 7530 22500
rect 9122 22448 9128 22500
rect 9180 22488 9186 22500
rect 11992 22488 12020 22528
rect 13170 22516 13176 22528
rect 13228 22516 13234 22568
rect 13538 22516 13544 22568
rect 13596 22556 13602 22568
rect 13633 22559 13691 22565
rect 13633 22556 13645 22559
rect 13596 22528 13645 22556
rect 13596 22516 13602 22528
rect 13633 22525 13645 22528
rect 13679 22556 13691 22559
rect 13906 22556 13912 22568
rect 13679 22528 13912 22556
rect 13679 22525 13691 22528
rect 13633 22519 13691 22525
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 14185 22559 14243 22565
rect 14185 22525 14197 22559
rect 14231 22525 14243 22559
rect 14550 22556 14556 22568
rect 14511 22528 14556 22556
rect 14185 22519 14243 22525
rect 9180 22460 12020 22488
rect 9180 22448 9186 22460
rect 1946 22380 1952 22432
rect 2004 22420 2010 22432
rect 5552 22420 5580 22448
rect 2004 22392 5580 22420
rect 2004 22380 2010 22392
rect 7282 22380 7288 22432
rect 7340 22420 7346 22432
rect 14090 22420 14096 22432
rect 7340 22392 14096 22420
rect 7340 22380 7346 22392
rect 14090 22380 14096 22392
rect 14148 22380 14154 22432
rect 14200 22420 14228 22519
rect 14550 22516 14556 22528
rect 14608 22516 14614 22568
rect 16776 22556 16804 22584
rect 16945 22559 17003 22565
rect 16945 22556 16957 22559
rect 15764 22528 16957 22556
rect 14458 22448 14464 22500
rect 14516 22488 14522 22500
rect 15764 22488 15792 22528
rect 16945 22525 16957 22528
rect 16991 22525 17003 22559
rect 17221 22559 17279 22565
rect 17221 22556 17233 22559
rect 16945 22519 17003 22525
rect 17052 22528 17233 22556
rect 14516 22460 15792 22488
rect 14516 22448 14522 22460
rect 16850 22448 16856 22500
rect 16908 22488 16914 22500
rect 17052 22488 17080 22528
rect 17221 22525 17233 22528
rect 17267 22556 17279 22559
rect 17788 22556 17816 22732
rect 18874 22720 18880 22732
rect 18932 22760 18938 22772
rect 22094 22760 22100 22772
rect 18932 22732 22100 22760
rect 18932 22720 18938 22732
rect 22094 22720 22100 22732
rect 22152 22720 22158 22772
rect 24780 22732 26648 22760
rect 18322 22652 18328 22704
rect 18380 22692 18386 22704
rect 18509 22695 18567 22701
rect 18509 22692 18521 22695
rect 18380 22664 18521 22692
rect 18380 22652 18386 22664
rect 18509 22661 18521 22664
rect 18555 22661 18567 22695
rect 18509 22655 18567 22661
rect 18601 22695 18659 22701
rect 18601 22661 18613 22695
rect 18647 22692 18659 22695
rect 18690 22692 18696 22704
rect 18647 22664 18696 22692
rect 18647 22661 18659 22664
rect 18601 22655 18659 22661
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 20806 22692 20812 22704
rect 20464 22664 20812 22692
rect 20346 22624 20352 22636
rect 19536 22596 20352 22624
rect 17267 22528 17816 22556
rect 17267 22525 17279 22528
rect 17221 22519 17279 22525
rect 18690 22516 18696 22568
rect 18748 22556 18754 22568
rect 18785 22559 18843 22565
rect 18785 22556 18797 22559
rect 18748 22528 18797 22556
rect 18748 22516 18754 22528
rect 18785 22525 18797 22528
rect 18831 22556 18843 22559
rect 19536 22556 19564 22596
rect 20346 22584 20352 22596
rect 20404 22584 20410 22636
rect 20464 22633 20492 22664
rect 20806 22652 20812 22664
rect 20864 22652 20870 22704
rect 22373 22695 22431 22701
rect 22373 22661 22385 22695
rect 22419 22692 22431 22695
rect 23658 22692 23664 22704
rect 22419 22664 23664 22692
rect 22419 22661 22431 22664
rect 22373 22655 22431 22661
rect 23658 22652 23664 22664
rect 23716 22652 23722 22704
rect 23934 22692 23940 22704
rect 23895 22664 23940 22692
rect 23934 22652 23940 22664
rect 23992 22652 23998 22704
rect 20441 22627 20499 22633
rect 20441 22593 20453 22627
rect 20487 22593 20499 22627
rect 20441 22587 20499 22593
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21100 22556 21128 22587
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 18831 22528 19564 22556
rect 19628 22528 21128 22556
rect 22204 22528 22293 22556
rect 18831 22525 18843 22528
rect 18785 22519 18843 22525
rect 16908 22460 17080 22488
rect 16908 22448 16914 22460
rect 17126 22448 17132 22500
rect 17184 22488 17190 22500
rect 17586 22488 17592 22500
rect 17184 22460 17592 22488
rect 17184 22448 17190 22460
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 14642 22420 14648 22432
rect 14200 22392 14648 22420
rect 14642 22380 14648 22392
rect 14700 22380 14706 22432
rect 14826 22380 14832 22432
rect 14884 22420 14890 22432
rect 16298 22420 16304 22432
rect 14884 22392 16304 22420
rect 14884 22380 14890 22392
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 19628 22420 19656 22528
rect 22204 22500 22232 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 22281 22519 22339 22525
rect 22370 22516 22376 22568
rect 22428 22556 22434 22568
rect 22554 22556 22560 22568
rect 22428 22528 22560 22556
rect 22428 22516 22434 22528
rect 22554 22516 22560 22528
rect 22612 22516 22618 22568
rect 23845 22559 23903 22565
rect 23845 22525 23857 22559
rect 23891 22556 23903 22559
rect 24780 22556 24808 22732
rect 25958 22692 25964 22704
rect 25919 22664 25964 22692
rect 25958 22652 25964 22664
rect 26016 22652 26022 22704
rect 26053 22695 26111 22701
rect 26053 22661 26065 22695
rect 26099 22692 26111 22695
rect 26234 22692 26240 22704
rect 26099 22664 26240 22692
rect 26099 22661 26111 22664
rect 26053 22655 26111 22661
rect 26234 22652 26240 22664
rect 26292 22652 26298 22704
rect 26620 22692 26648 22732
rect 26694 22720 26700 22772
rect 26752 22760 26758 22772
rect 27249 22763 27307 22769
rect 27249 22760 27261 22763
rect 26752 22732 27261 22760
rect 26752 22720 26758 22732
rect 27249 22729 27261 22732
rect 27295 22729 27307 22763
rect 28074 22760 28080 22772
rect 28035 22732 28080 22760
rect 27249 22723 27307 22729
rect 28074 22720 28080 22732
rect 28132 22720 28138 22772
rect 28350 22692 28356 22704
rect 26620 22664 28356 22692
rect 28350 22652 28356 22664
rect 28408 22652 28414 22704
rect 29362 22692 29368 22704
rect 29323 22664 29368 22692
rect 29362 22652 29368 22664
rect 29420 22652 29426 22704
rect 27062 22584 27068 22636
rect 27120 22624 27126 22636
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 27120 22596 27169 22624
rect 27120 22584 27126 22596
rect 27157 22593 27169 22596
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 27985 22627 28043 22633
rect 27985 22593 27997 22627
rect 28031 22624 28043 22627
rect 28994 22624 29000 22636
rect 28031 22596 29000 22624
rect 28031 22593 28043 22596
rect 27985 22587 28043 22593
rect 28994 22584 29000 22596
rect 29052 22584 29058 22636
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22624 30803 22627
rect 37550 22624 37556 22636
rect 30791 22596 37556 22624
rect 30791 22593 30803 22596
rect 30745 22587 30803 22593
rect 37550 22584 37556 22596
rect 37608 22584 37614 22636
rect 38010 22624 38016 22636
rect 37971 22596 38016 22624
rect 38010 22584 38016 22596
rect 38068 22584 38074 22636
rect 23891 22528 24808 22556
rect 23891 22525 23903 22528
rect 23845 22519 23903 22525
rect 24854 22516 24860 22568
rect 24912 22556 24918 22568
rect 29270 22556 29276 22568
rect 24912 22528 24957 22556
rect 26206 22528 28994 22556
rect 29231 22528 29276 22556
rect 24912 22516 24918 22528
rect 20806 22448 20812 22500
rect 20864 22488 20870 22500
rect 21910 22488 21916 22500
rect 20864 22460 21916 22488
rect 20864 22448 20870 22460
rect 21910 22448 21916 22460
rect 21968 22448 21974 22500
rect 22186 22448 22192 22500
rect 22244 22448 22250 22500
rect 26206 22488 26234 22528
rect 26510 22488 26516 22500
rect 22296 22460 26234 22488
rect 26471 22460 26516 22488
rect 16632 22392 19656 22420
rect 20533 22423 20591 22429
rect 16632 22380 16638 22392
rect 20533 22389 20545 22423
rect 20579 22420 20591 22423
rect 20622 22420 20628 22432
rect 20579 22392 20628 22420
rect 20579 22389 20591 22392
rect 20533 22383 20591 22389
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 21177 22423 21235 22429
rect 21177 22389 21189 22423
rect 21223 22420 21235 22423
rect 21266 22420 21272 22432
rect 21223 22392 21272 22420
rect 21223 22389 21235 22392
rect 21177 22383 21235 22389
rect 21266 22380 21272 22392
rect 21324 22380 21330 22432
rect 21450 22380 21456 22432
rect 21508 22420 21514 22432
rect 22296 22420 22324 22460
rect 26510 22448 26516 22460
rect 26568 22448 26574 22500
rect 28966 22488 28994 22528
rect 29270 22516 29276 22528
rect 29328 22516 29334 22568
rect 29546 22556 29552 22568
rect 29507 22528 29552 22556
rect 29546 22516 29552 22528
rect 29604 22516 29610 22568
rect 30837 22491 30895 22497
rect 30837 22488 30849 22491
rect 28966 22460 30849 22488
rect 30837 22457 30849 22460
rect 30883 22457 30895 22491
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 30837 22451 30895 22457
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 21508 22392 22324 22420
rect 21508 22380 21514 22392
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 26602 22420 26608 22432
rect 23440 22392 26608 22420
rect 23440 22380 23446 22392
rect 26602 22380 26608 22392
rect 26660 22380 26666 22432
rect 29178 22380 29184 22432
rect 29236 22420 29242 22432
rect 29546 22420 29552 22432
rect 29236 22392 29552 22420
rect 29236 22380 29242 22392
rect 29546 22380 29552 22392
rect 29604 22380 29610 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 2406 22176 2412 22228
rect 2464 22216 2470 22228
rect 4322 22219 4380 22225
rect 4322 22216 4334 22219
rect 2464 22188 4334 22216
rect 2464 22176 2470 22188
rect 4322 22185 4334 22188
rect 4368 22185 4380 22219
rect 4322 22179 4380 22185
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6536 22219 6594 22225
rect 6536 22216 6548 22219
rect 6236 22188 6548 22216
rect 6236 22176 6242 22188
rect 6536 22185 6548 22188
rect 6582 22216 6594 22219
rect 9122 22216 9128 22228
rect 6582 22188 7972 22216
rect 6582 22185 6594 22188
rect 6536 22179 6594 22185
rect 5626 22108 5632 22160
rect 5684 22148 5690 22160
rect 7944 22148 7972 22188
rect 8588 22188 9128 22216
rect 8588 22148 8616 22188
rect 9122 22176 9128 22188
rect 9180 22176 9186 22228
rect 9214 22176 9220 22228
rect 9272 22216 9278 22228
rect 11146 22216 11152 22228
rect 9272 22188 11152 22216
rect 9272 22176 9278 22188
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 14458 22216 14464 22228
rect 11440 22188 14464 22216
rect 5684 22120 6132 22148
rect 7944 22120 8616 22148
rect 9140 22120 10088 22148
rect 5684 22108 5690 22120
rect 1670 22080 1676 22092
rect 1631 22052 1676 22080
rect 1670 22040 1676 22052
rect 1728 22040 1734 22092
rect 1946 22080 1952 22092
rect 1907 22052 1952 22080
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 3421 22083 3479 22089
rect 3421 22049 3433 22083
rect 3467 22080 3479 22083
rect 3510 22080 3516 22092
rect 3467 22052 3516 22080
rect 3467 22049 3479 22052
rect 3421 22043 3479 22049
rect 3510 22040 3516 22052
rect 3568 22040 3574 22092
rect 3970 22054 3976 22106
rect 4028 22094 4034 22106
rect 4028 22080 4200 22094
rect 5902 22080 5908 22092
rect 4028 22066 5488 22080
rect 4028 22054 4034 22066
rect 4172 22052 5488 22066
rect 4062 22012 4068 22024
rect 4023 21984 4068 22012
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 5460 21998 5488 22052
rect 5644 22052 5908 22080
rect 5644 22024 5672 22052
rect 5902 22040 5908 22052
rect 5960 22040 5966 22092
rect 5626 21972 5632 22024
rect 5684 21972 5690 22024
rect 4430 21944 4436 21956
rect 3174 21916 4436 21944
rect 4430 21904 4436 21916
rect 4488 21904 4494 21956
rect 6104 21944 6132 22120
rect 6270 22080 6276 22092
rect 6231 22052 6276 22080
rect 6270 22040 6276 22052
rect 6328 22040 6334 22092
rect 7006 22040 7012 22092
rect 7064 22080 7070 22092
rect 7064 22052 7604 22080
rect 7064 22040 7070 22052
rect 7576 22024 7604 22052
rect 8662 22040 8668 22092
rect 8720 22080 8726 22092
rect 9140 22080 9168 22120
rect 10060 22092 10088 22120
rect 10502 22108 10508 22160
rect 10560 22108 10566 22160
rect 11440 22148 11468 22188
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 16758 22216 16764 22228
rect 15120 22188 16764 22216
rect 10612 22120 11468 22148
rect 8720 22052 9168 22080
rect 9217 22083 9275 22089
rect 8720 22040 8726 22052
rect 9217 22049 9229 22083
rect 9263 22080 9275 22083
rect 9674 22080 9680 22092
rect 9263 22052 9680 22080
rect 9263 22049 9275 22052
rect 9217 22043 9275 22049
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 10042 22080 10048 22092
rect 10003 22052 10048 22080
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 10520 22080 10548 22108
rect 10612 22089 10640 22120
rect 10428 22052 10548 22080
rect 10597 22083 10655 22089
rect 7558 21972 7564 22024
rect 7616 21972 7622 22024
rect 6270 21944 6276 21956
rect 6104 21916 6276 21944
rect 6270 21904 6276 21916
rect 6328 21904 6334 21956
rect 8202 21944 8208 21956
rect 7774 21916 8208 21944
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 9309 21947 9367 21953
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 9398 21944 9404 21956
rect 9355 21916 9404 21944
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 10428 21944 10456 22052
rect 10597 22049 10609 22083
rect 10643 22049 10655 22083
rect 11606 22080 11612 22092
rect 11519 22052 11612 22080
rect 10597 22043 10655 22049
rect 11606 22040 11612 22052
rect 11664 22080 11670 22092
rect 11664 22052 13124 22080
rect 11664 22040 11670 22052
rect 10502 21972 10508 22024
rect 10560 22012 10566 22024
rect 10560 21984 10605 22012
rect 10560 21972 10566 21984
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11333 22015 11391 22021
rect 11333 22012 11345 22015
rect 11020 21984 11345 22012
rect 11020 21972 11026 21984
rect 11333 21981 11345 21984
rect 11379 21981 11391 22015
rect 11333 21975 11391 21981
rect 12710 21972 12716 22024
rect 12768 21972 12774 22024
rect 13096 22012 13124 22052
rect 13170 22040 13176 22092
rect 13228 22080 13234 22092
rect 13357 22083 13415 22089
rect 13357 22080 13369 22083
rect 13228 22052 13369 22080
rect 13228 22040 13234 22052
rect 13357 22049 13369 22052
rect 13403 22049 13415 22083
rect 13357 22043 13415 22049
rect 14182 22040 14188 22092
rect 14240 22080 14246 22092
rect 14645 22083 14703 22089
rect 14645 22080 14657 22083
rect 14240 22052 14657 22080
rect 14240 22040 14246 22052
rect 14645 22049 14657 22052
rect 14691 22049 14703 22083
rect 14645 22043 14703 22049
rect 13814 22012 13820 22024
rect 13096 21984 13820 22012
rect 13814 21972 13820 21984
rect 13872 21972 13878 22024
rect 14553 22015 14611 22021
rect 14553 21981 14565 22015
rect 14599 22012 14611 22015
rect 15010 22012 15016 22024
rect 14599 21984 15016 22012
rect 14599 21981 14611 21984
rect 14553 21975 14611 21981
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 9876 21916 10456 21944
rect 11057 21947 11115 21953
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 5810 21876 5816 21888
rect 3292 21848 5816 21876
rect 3292 21836 3298 21848
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 7190 21836 7196 21888
rect 7248 21876 7254 21888
rect 8021 21879 8079 21885
rect 8021 21876 8033 21879
rect 7248 21848 8033 21876
rect 7248 21836 7254 21848
rect 8021 21845 8033 21848
rect 8067 21845 8079 21879
rect 8021 21839 8079 21845
rect 8662 21836 8668 21888
rect 8720 21876 8726 21888
rect 9876 21876 9904 21916
rect 11057 21913 11069 21947
rect 11103 21944 11115 21947
rect 11606 21944 11612 21956
rect 11103 21916 11612 21944
rect 11103 21913 11115 21916
rect 11057 21907 11115 21913
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 15120 21944 15148 22188
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 17494 22216 17500 22228
rect 16868 22188 17500 22216
rect 15194 22108 15200 22160
rect 15252 22148 15258 22160
rect 15252 22120 16160 22148
rect 15252 22108 15258 22120
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 16022 22080 16028 22092
rect 15335 22052 16028 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 16022 22040 16028 22052
rect 16080 22040 16086 22092
rect 16132 22080 16160 22120
rect 16482 22108 16488 22160
rect 16540 22148 16546 22160
rect 16868 22148 16896 22188
rect 17494 22176 17500 22188
rect 17552 22176 17558 22228
rect 18141 22219 18199 22225
rect 18141 22185 18153 22219
rect 18187 22216 18199 22219
rect 18598 22216 18604 22228
rect 18187 22188 18604 22216
rect 18187 22185 18199 22188
rect 18141 22179 18199 22185
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 20070 22216 20076 22228
rect 20031 22188 20076 22216
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 22922 22216 22928 22228
rect 20496 22188 22928 22216
rect 20496 22176 20502 22188
rect 22922 22176 22928 22188
rect 22980 22176 22986 22228
rect 23934 22176 23940 22228
rect 23992 22216 23998 22228
rect 24673 22219 24731 22225
rect 24673 22216 24685 22219
rect 23992 22188 24685 22216
rect 23992 22176 23998 22188
rect 24673 22185 24685 22188
rect 24719 22185 24731 22219
rect 24673 22179 24731 22185
rect 16540 22120 16896 22148
rect 16540 22108 16546 22120
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 26418 22148 26424 22160
rect 17276 22120 26424 22148
rect 17276 22108 17282 22120
rect 26418 22108 26424 22120
rect 26476 22148 26482 22160
rect 27062 22148 27068 22160
rect 26476 22120 27068 22148
rect 26476 22108 26482 22120
rect 27062 22108 27068 22120
rect 27120 22108 27126 22160
rect 28905 22151 28963 22157
rect 28905 22117 28917 22151
rect 28951 22148 28963 22151
rect 30650 22148 30656 22160
rect 28951 22120 30656 22148
rect 28951 22117 28963 22120
rect 28905 22111 28963 22117
rect 30650 22108 30656 22120
rect 30708 22108 30714 22160
rect 16132 22052 18644 22080
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 17218 22012 17224 22024
rect 17175 21984 17224 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 17954 21972 17960 22024
rect 18012 22012 18018 22024
rect 18049 22015 18107 22021
rect 18049 22012 18061 22015
rect 18012 21984 18061 22012
rect 18012 21972 18018 21984
rect 18049 21981 18061 21984
rect 18095 21981 18107 22015
rect 18616 22014 18644 22052
rect 19426 22040 19432 22092
rect 19484 22080 19490 22092
rect 20717 22083 20775 22089
rect 20717 22080 20729 22083
rect 19484 22052 20729 22080
rect 19484 22040 19490 22052
rect 20717 22049 20729 22052
rect 20763 22049 20775 22083
rect 21358 22080 21364 22092
rect 21319 22052 21364 22080
rect 20717 22043 20775 22049
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 22278 22080 22284 22092
rect 22239 22052 22284 22080
rect 22278 22040 22284 22052
rect 22336 22040 22342 22092
rect 23566 22040 23572 22092
rect 23624 22080 23630 22092
rect 23750 22080 23756 22092
rect 23624 22052 23756 22080
rect 23624 22040 23630 22052
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 24029 22083 24087 22089
rect 24029 22049 24041 22083
rect 24075 22080 24087 22083
rect 26510 22080 26516 22092
rect 24075 22052 26516 22080
rect 24075 22049 24087 22052
rect 24029 22043 24087 22049
rect 26510 22040 26516 22052
rect 26568 22040 26574 22092
rect 26970 22080 26976 22092
rect 26931 22052 26976 22080
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 28626 22080 28632 22092
rect 28184 22052 28632 22080
rect 18693 22015 18751 22021
rect 18693 22014 18705 22015
rect 18616 21986 18705 22014
rect 18049 21975 18107 21981
rect 18693 21981 18705 21986
rect 18739 21981 18751 22015
rect 19981 22015 20039 22021
rect 19981 22012 19993 22015
rect 18693 21975 18751 21981
rect 19904 21984 19993 22012
rect 15378 21953 15384 21956
rect 13096 21916 15148 21944
rect 15358 21947 15384 21953
rect 8720 21848 9904 21876
rect 8720 21836 8726 21848
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 13096 21876 13124 21916
rect 15358 21913 15370 21947
rect 15358 21907 15384 21913
rect 15378 21904 15384 21907
rect 15436 21904 15442 21956
rect 15930 21944 15936 21956
rect 15891 21916 15936 21944
rect 15930 21904 15936 21916
rect 15988 21904 15994 21956
rect 16482 21944 16488 21956
rect 16443 21916 16488 21944
rect 16482 21904 16488 21916
rect 16540 21904 16546 21956
rect 16574 21904 16580 21956
rect 16632 21944 16638 21956
rect 16632 21916 16677 21944
rect 16632 21904 16638 21916
rect 16758 21904 16764 21956
rect 16816 21944 16822 21956
rect 19904 21944 19932 21984
rect 19981 21981 19993 21984
rect 20027 21981 20039 22015
rect 22186 22012 22192 22024
rect 22147 21984 22192 22012
rect 19981 21975 20039 21981
rect 22186 21972 22192 21984
rect 22244 21972 22250 22024
rect 24486 21972 24492 22024
rect 24544 22012 24550 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 24544 21984 24593 22012
rect 24544 21972 24550 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 16816 21916 19932 21944
rect 20809 21947 20867 21953
rect 16816 21904 16822 21916
rect 20809 21913 20821 21947
rect 20855 21944 20867 21947
rect 21266 21944 21272 21956
rect 20855 21916 21272 21944
rect 20855 21913 20867 21916
rect 20809 21907 20867 21913
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 22094 21904 22100 21956
rect 22152 21944 22158 21956
rect 23198 21944 23204 21956
rect 22152 21916 23204 21944
rect 22152 21904 22158 21916
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 23382 21944 23388 21956
rect 23343 21916 23388 21944
rect 23382 21904 23388 21916
rect 23440 21904 23446 21956
rect 23477 21947 23535 21953
rect 23477 21913 23489 21947
rect 23523 21944 23535 21947
rect 24210 21944 24216 21956
rect 23523 21916 24216 21944
rect 23523 21913 23535 21916
rect 23477 21907 23535 21913
rect 24210 21904 24216 21916
rect 24268 21904 24274 21956
rect 26528 21944 26556 22040
rect 26878 22012 26884 22024
rect 26839 21984 26884 22012
rect 26878 21972 26884 21984
rect 26936 21972 26942 22024
rect 28184 21944 28212 22052
rect 28626 22040 28632 22052
rect 28684 22040 28690 22092
rect 33778 21972 33784 22024
rect 33836 22012 33842 22024
rect 34149 22015 34207 22021
rect 34149 22012 34161 22015
rect 33836 21984 34161 22012
rect 33836 21972 33842 21984
rect 34149 21981 34161 21984
rect 34195 21981 34207 22015
rect 38286 22012 38292 22024
rect 38247 21984 38292 22012
rect 34149 21975 34207 21981
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 28353 21947 28411 21953
rect 28353 21944 28365 21947
rect 26528 21916 28365 21944
rect 28353 21913 28365 21916
rect 28399 21913 28411 21947
rect 28353 21907 28411 21913
rect 28445 21947 28503 21953
rect 28445 21913 28457 21947
rect 28491 21913 28503 21947
rect 28445 21907 28503 21913
rect 12492 21848 13124 21876
rect 12492 21836 12498 21848
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 15654 21876 15660 21888
rect 13228 21848 15660 21876
rect 13228 21836 13234 21848
rect 15654 21836 15660 21848
rect 15712 21836 15718 21888
rect 15838 21836 15844 21888
rect 15896 21876 15902 21888
rect 16942 21876 16948 21888
rect 15896 21848 16948 21876
rect 15896 21836 15902 21848
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17402 21876 17408 21888
rect 17092 21848 17408 21876
rect 17092 21836 17098 21848
rect 17402 21836 17408 21848
rect 17460 21836 17466 21888
rect 18782 21876 18788 21888
rect 18743 21848 18788 21876
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 22646 21836 22652 21888
rect 22704 21876 22710 21888
rect 28460 21876 28488 21907
rect 32674 21904 32680 21956
rect 32732 21944 32738 21956
rect 32732 21916 35894 21944
rect 32732 21904 32738 21916
rect 22704 21848 28488 21876
rect 22704 21836 22710 21848
rect 33594 21836 33600 21888
rect 33652 21876 33658 21888
rect 33965 21879 34023 21885
rect 33965 21876 33977 21879
rect 33652 21848 33977 21876
rect 33652 21836 33658 21848
rect 33965 21845 33977 21848
rect 34011 21845 34023 21879
rect 35866 21876 35894 21916
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 35866 21848 38117 21876
rect 33965 21839 34023 21845
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2498 21632 2504 21684
rect 2556 21672 2562 21684
rect 3234 21672 3240 21684
rect 2556 21644 3240 21672
rect 2556 21632 2562 21644
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 3326 21632 3332 21684
rect 3384 21632 3390 21684
rect 4617 21675 4675 21681
rect 4617 21641 4629 21675
rect 4663 21672 4675 21675
rect 5074 21672 5080 21684
rect 4663 21644 5080 21672
rect 4663 21641 4675 21644
rect 4617 21635 4675 21641
rect 5074 21632 5080 21644
rect 5132 21632 5138 21684
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 6454 21672 6460 21684
rect 5408 21644 6460 21672
rect 5408 21632 5414 21644
rect 6454 21632 6460 21644
rect 6512 21632 6518 21684
rect 9214 21672 9220 21684
rect 7852 21644 9220 21672
rect 1854 21564 1860 21616
rect 1912 21604 1918 21616
rect 3145 21607 3203 21613
rect 1912 21576 2728 21604
rect 1912 21564 1918 21576
rect 1578 21536 1584 21548
rect 1539 21508 1584 21536
rect 1578 21496 1584 21508
rect 1636 21496 1642 21548
rect 2700 21536 2728 21576
rect 3145 21573 3157 21607
rect 3191 21604 3203 21607
rect 3344 21604 3372 21632
rect 5166 21604 5172 21616
rect 3191 21576 3372 21604
rect 4370 21576 5172 21604
rect 3191 21573 3203 21576
rect 3145 21567 3203 21573
rect 5166 21564 5172 21576
rect 5224 21564 5230 21616
rect 5445 21607 5503 21613
rect 5445 21573 5457 21607
rect 5491 21604 5503 21607
rect 6638 21604 6644 21616
rect 5491 21576 6644 21604
rect 5491 21573 5503 21576
rect 5445 21567 5503 21573
rect 6638 21564 6644 21576
rect 6696 21564 6702 21616
rect 7006 21564 7012 21616
rect 7064 21604 7070 21616
rect 7852 21613 7880 21644
rect 9214 21632 9220 21644
rect 9272 21632 9278 21684
rect 11238 21672 11244 21684
rect 9876 21644 11244 21672
rect 7837 21607 7895 21613
rect 7064 21576 7604 21604
rect 7064 21564 7070 21576
rect 2869 21539 2927 21545
rect 2869 21536 2881 21539
rect 2700 21508 2881 21536
rect 2869 21505 2881 21508
rect 2915 21505 2927 21539
rect 2869 21499 2927 21505
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21536 6975 21539
rect 7190 21536 7196 21548
rect 6963 21508 7196 21536
rect 6963 21505 6975 21508
rect 6917 21499 6975 21505
rect 7190 21496 7196 21508
rect 7248 21496 7254 21548
rect 7576 21545 7604 21576
rect 7837 21573 7849 21607
rect 7883 21573 7895 21607
rect 7837 21567 7895 21573
rect 8846 21564 8852 21616
rect 8904 21564 8910 21616
rect 9585 21607 9643 21613
rect 9585 21573 9597 21607
rect 9631 21604 9643 21607
rect 9876 21604 9904 21644
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 11333 21675 11391 21681
rect 11333 21641 11345 21675
rect 11379 21672 11391 21675
rect 11606 21672 11612 21684
rect 11379 21644 11612 21672
rect 11379 21641 11391 21644
rect 11333 21635 11391 21641
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 15378 21672 15384 21684
rect 11716 21644 15384 21672
rect 9631 21576 9904 21604
rect 9631 21573 9643 21576
rect 9585 21567 9643 21573
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21505 7619 21539
rect 7561 21499 7619 21505
rect 1857 21471 1915 21477
rect 1857 21437 1869 21471
rect 1903 21468 1915 21471
rect 1946 21468 1952 21480
rect 1903 21440 1952 21468
rect 1903 21437 1915 21440
rect 1857 21431 1915 21437
rect 1946 21428 1952 21440
rect 2004 21468 2010 21480
rect 2498 21468 2504 21480
rect 2004 21440 2504 21468
rect 2004 21428 2010 21440
rect 2498 21428 2504 21440
rect 2556 21428 2562 21480
rect 4522 21428 4528 21480
rect 4580 21468 4586 21480
rect 4706 21468 4712 21480
rect 4580 21440 4712 21468
rect 4580 21428 4586 21440
rect 4706 21428 4712 21440
rect 4764 21428 4770 21480
rect 5166 21428 5172 21480
rect 5224 21468 5230 21480
rect 5353 21471 5411 21477
rect 5353 21468 5365 21471
rect 5224 21440 5365 21468
rect 5224 21428 5230 21440
rect 5353 21437 5365 21440
rect 5399 21437 5411 21471
rect 7466 21468 7472 21480
rect 5353 21431 5411 21437
rect 5828 21440 7472 21468
rect 4430 21360 4436 21412
rect 4488 21400 4494 21412
rect 5828 21400 5856 21440
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 8386 21468 8392 21480
rect 7668 21440 8392 21468
rect 4488 21372 5856 21400
rect 5905 21403 5963 21409
rect 4488 21360 4494 21372
rect 5905 21369 5917 21403
rect 5951 21400 5963 21403
rect 6822 21400 6828 21412
rect 5951 21372 6828 21400
rect 5951 21369 5963 21372
rect 5905 21363 5963 21369
rect 6822 21360 6828 21372
rect 6880 21360 6886 21412
rect 7668 21400 7696 21440
rect 8386 21428 8392 21440
rect 8444 21428 8450 21480
rect 6932 21372 7696 21400
rect 9876 21400 9904 21576
rect 9950 21564 9956 21616
rect 10008 21604 10014 21616
rect 10781 21607 10839 21613
rect 10781 21604 10793 21607
rect 10008 21576 10793 21604
rect 10008 21564 10014 21576
rect 10781 21573 10793 21576
rect 10827 21573 10839 21607
rect 11716 21604 11744 21644
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 18690 21672 18696 21684
rect 15488 21644 18696 21672
rect 10781 21567 10839 21573
rect 10888 21576 11744 21604
rect 11885 21607 11943 21613
rect 10045 21539 10103 21545
rect 10045 21536 10057 21539
rect 9968 21508 10057 21536
rect 9968 21480 9996 21508
rect 10045 21505 10057 21508
rect 10091 21536 10103 21539
rect 10226 21536 10232 21548
rect 10091 21508 10232 21536
rect 10091 21505 10103 21508
rect 10045 21499 10103 21505
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 10594 21496 10600 21548
rect 10652 21536 10658 21548
rect 10888 21536 10916 21576
rect 11885 21573 11897 21607
rect 11931 21604 11943 21607
rect 11974 21604 11980 21616
rect 11931 21576 11980 21604
rect 11931 21573 11943 21576
rect 11885 21567 11943 21573
rect 11974 21564 11980 21576
rect 12032 21564 12038 21616
rect 12250 21564 12256 21616
rect 12308 21604 12314 21616
rect 13725 21607 13783 21613
rect 13725 21604 13737 21607
rect 12308 21576 13737 21604
rect 12308 21564 12314 21576
rect 13725 21573 13737 21576
rect 13771 21573 13783 21607
rect 13725 21567 13783 21573
rect 14090 21564 14096 21616
rect 14148 21604 14154 21616
rect 14277 21607 14335 21613
rect 14277 21604 14289 21607
rect 14148 21576 14289 21604
rect 14148 21564 14154 21576
rect 14277 21573 14289 21576
rect 14323 21604 14335 21607
rect 15488 21604 15516 21644
rect 18690 21632 18696 21644
rect 18748 21632 18754 21684
rect 18782 21632 18788 21684
rect 18840 21672 18846 21684
rect 21266 21672 21272 21684
rect 18840 21644 20492 21672
rect 21227 21644 21272 21672
rect 18840 21632 18846 21644
rect 14323 21576 15516 21604
rect 15749 21607 15807 21613
rect 14323 21573 14335 21576
rect 14277 21567 14335 21573
rect 15749 21573 15761 21607
rect 15795 21604 15807 21607
rect 15838 21604 15844 21616
rect 15795 21576 15844 21604
rect 15795 21573 15807 21576
rect 15749 21567 15807 21573
rect 15838 21564 15844 21576
rect 15896 21564 15902 21616
rect 18138 21604 18144 21616
rect 17604 21576 18144 21604
rect 10652 21508 10916 21536
rect 14921 21539 14979 21545
rect 10652 21496 10658 21508
rect 14921 21505 14933 21539
rect 14967 21536 14979 21539
rect 15010 21536 15016 21548
rect 14967 21508 15016 21536
rect 14967 21505 14979 21508
rect 14921 21499 14979 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 17126 21536 17132 21548
rect 16356 21508 16401 21536
rect 17087 21508 17132 21536
rect 16356 21496 16362 21508
rect 17126 21496 17132 21508
rect 17184 21496 17190 21548
rect 9950 21428 9956 21480
rect 10008 21428 10014 21480
rect 11790 21468 11796 21480
rect 11751 21440 11796 21468
rect 11790 21428 11796 21440
rect 11848 21428 11854 21480
rect 12805 21471 12863 21477
rect 12805 21437 12817 21471
rect 12851 21468 12863 21471
rect 12894 21468 12900 21480
rect 12851 21440 12900 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 12986 21428 12992 21480
rect 13044 21468 13050 21480
rect 13633 21471 13691 21477
rect 13633 21468 13645 21471
rect 13044 21440 13645 21468
rect 13044 21428 13050 21440
rect 13633 21437 13645 21440
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 14826 21468 14832 21480
rect 14148 21440 14832 21468
rect 14148 21428 14154 21440
rect 14826 21428 14832 21440
rect 14884 21428 14890 21480
rect 15657 21471 15715 21477
rect 15657 21437 15669 21471
rect 15703 21468 15715 21471
rect 15838 21468 15844 21480
rect 15703 21440 15844 21468
rect 15703 21437 15715 21440
rect 15657 21431 15715 21437
rect 15838 21428 15844 21440
rect 15896 21428 15902 21480
rect 16022 21428 16028 21480
rect 16080 21468 16086 21480
rect 17604 21468 17632 21576
rect 18138 21564 18144 21576
rect 18196 21564 18202 21616
rect 18506 21604 18512 21616
rect 18467 21576 18512 21604
rect 18506 21564 18512 21576
rect 18564 21564 18570 21616
rect 18601 21607 18659 21613
rect 18601 21573 18613 21607
rect 18647 21604 18659 21607
rect 19797 21607 19855 21613
rect 18647 21576 19334 21604
rect 18647 21573 18659 21576
rect 18601 21567 18659 21573
rect 17770 21536 17776 21548
rect 17731 21508 17776 21536
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 19306 21536 19334 21576
rect 19797 21573 19809 21607
rect 19843 21604 19855 21607
rect 20162 21604 20168 21616
rect 19843 21576 20168 21604
rect 19843 21573 19855 21576
rect 19797 21567 19855 21573
rect 20162 21564 20168 21576
rect 20220 21564 20226 21616
rect 20464 21604 20492 21644
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 23474 21632 23480 21684
rect 23532 21672 23538 21684
rect 23569 21675 23627 21681
rect 23569 21672 23581 21675
rect 23532 21644 23581 21672
rect 23532 21632 23538 21644
rect 23569 21641 23581 21644
rect 23615 21641 23627 21675
rect 24210 21672 24216 21684
rect 24171 21644 24216 21672
rect 23569 21635 23627 21641
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 24854 21632 24860 21684
rect 24912 21672 24918 21684
rect 30742 21672 30748 21684
rect 24912 21644 30748 21672
rect 24912 21632 24918 21644
rect 30742 21632 30748 21644
rect 30800 21632 30806 21684
rect 38194 21672 38200 21684
rect 38155 21644 38200 21672
rect 38194 21632 38200 21644
rect 38252 21632 38258 21684
rect 21910 21604 21916 21616
rect 20464 21576 21916 21604
rect 21910 21564 21916 21576
rect 21968 21564 21974 21616
rect 26513 21607 26571 21613
rect 22020 21576 25452 21604
rect 22020 21548 22048 21576
rect 21174 21536 21180 21548
rect 19306 21508 19472 21536
rect 21135 21508 21180 21536
rect 16080 21440 17632 21468
rect 17865 21471 17923 21477
rect 16080 21428 16086 21440
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 19334 21468 19340 21480
rect 17911 21440 19340 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 19334 21428 19340 21440
rect 19392 21428 19398 21480
rect 10502 21400 10508 21412
rect 9876 21372 10508 21400
rect 5626 21292 5632 21344
rect 5684 21332 5690 21344
rect 6932 21332 6960 21372
rect 10502 21360 10508 21372
rect 10560 21360 10566 21412
rect 13906 21400 13912 21412
rect 10704 21372 13912 21400
rect 5684 21304 6960 21332
rect 7009 21335 7067 21341
rect 5684 21292 5690 21304
rect 7009 21301 7021 21335
rect 7055 21332 7067 21335
rect 10704 21332 10732 21372
rect 13906 21360 13912 21372
rect 13964 21360 13970 21412
rect 17221 21403 17279 21409
rect 17221 21400 17233 21403
rect 14292 21372 17233 21400
rect 7055 21304 10732 21332
rect 7055 21301 7067 21304
rect 7009 21295 7067 21301
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 12434 21332 12440 21344
rect 11848 21304 12440 21332
rect 11848 21292 11854 21304
rect 12434 21292 12440 21304
rect 12492 21292 12498 21344
rect 12526 21292 12532 21344
rect 12584 21332 12590 21344
rect 14292 21332 14320 21372
rect 17221 21369 17233 21372
rect 17267 21369 17279 21403
rect 18782 21400 18788 21412
rect 17221 21363 17279 21369
rect 17788 21372 18788 21400
rect 12584 21304 14320 21332
rect 15013 21335 15071 21341
rect 12584 21292 12590 21304
rect 15013 21301 15025 21335
rect 15059 21332 15071 21335
rect 17788 21332 17816 21372
rect 18782 21360 18788 21372
rect 18840 21360 18846 21412
rect 19061 21403 19119 21409
rect 19061 21369 19073 21403
rect 19107 21369 19119 21403
rect 19061 21363 19119 21369
rect 15059 21304 17816 21332
rect 15059 21301 15071 21304
rect 15013 21295 15071 21301
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 19076 21332 19104 21363
rect 18196 21304 19104 21332
rect 19444 21332 19472 21508
rect 21174 21496 21180 21508
rect 21232 21536 21238 21548
rect 21542 21536 21548 21548
rect 21232 21508 21548 21536
rect 21232 21496 21238 21508
rect 21542 21496 21548 21508
rect 21600 21496 21606 21548
rect 22002 21536 22008 21548
rect 21963 21508 22008 21536
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 23014 21536 23020 21548
rect 22879 21508 23020 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 23474 21536 23480 21548
rect 23435 21508 23480 21536
rect 23474 21496 23480 21508
rect 23532 21536 23538 21548
rect 23842 21536 23848 21548
rect 23532 21508 23848 21536
rect 23532 21496 23538 21508
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 24118 21536 24124 21548
rect 24079 21508 24124 21536
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24210 21496 24216 21548
rect 24268 21536 24274 21548
rect 25424 21545 25452 21576
rect 26513 21573 26525 21607
rect 26559 21604 26571 21607
rect 27341 21607 27399 21613
rect 27341 21604 27353 21607
rect 26559 21576 27353 21604
rect 26559 21573 26571 21576
rect 26513 21567 26571 21573
rect 27341 21573 27353 21576
rect 27387 21573 27399 21607
rect 28902 21604 28908 21616
rect 28863 21576 28908 21604
rect 27341 21567 27399 21573
rect 28902 21564 28908 21576
rect 28960 21564 28966 21616
rect 28994 21564 29000 21616
rect 29052 21604 29058 21616
rect 29052 21576 29960 21604
rect 29052 21564 29058 21576
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24268 21508 24777 21536
rect 24268 21496 24274 21508
rect 24765 21505 24777 21508
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 25409 21539 25467 21545
rect 25409 21505 25421 21539
rect 25455 21505 25467 21539
rect 26418 21536 26424 21548
rect 26379 21508 26424 21536
rect 25409 21499 25467 21505
rect 26418 21496 26424 21508
rect 26476 21496 26482 21548
rect 29932 21545 29960 21576
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21536 29975 21539
rect 37550 21536 37556 21548
rect 29963 21508 37556 21536
rect 29963 21505 29975 21508
rect 29917 21499 29975 21505
rect 37550 21496 37556 21508
rect 37608 21496 37614 21548
rect 38102 21536 38108 21548
rect 38063 21508 38108 21536
rect 38102 21496 38108 21508
rect 38160 21496 38166 21548
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21437 19763 21471
rect 20254 21468 20260 21480
rect 20215 21440 20260 21468
rect 19705 21431 19763 21437
rect 19720 21400 19748 21431
rect 20254 21428 20260 21440
rect 20312 21468 20318 21480
rect 20714 21468 20720 21480
rect 20312 21440 20720 21468
rect 20312 21428 20318 21440
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 22094 21468 22100 21480
rect 21928 21440 22100 21468
rect 21928 21400 21956 21440
rect 22094 21428 22100 21440
rect 22152 21428 22158 21480
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 25501 21471 25559 21477
rect 25501 21468 25513 21471
rect 22244 21440 25513 21468
rect 22244 21428 22250 21440
rect 25501 21437 25513 21440
rect 25547 21437 25559 21471
rect 25501 21431 25559 21437
rect 27249 21471 27307 21477
rect 27249 21437 27261 21471
rect 27295 21437 27307 21471
rect 27249 21431 27307 21437
rect 19720 21372 21956 21400
rect 21082 21332 21088 21344
rect 19444 21304 21088 21332
rect 18196 21292 18202 21304
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 22097 21335 22155 21341
rect 22097 21301 22109 21335
rect 22143 21332 22155 21335
rect 22186 21332 22192 21344
rect 22143 21304 22192 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 22925 21335 22983 21341
rect 22925 21332 22937 21335
rect 22520 21304 22937 21332
rect 22520 21292 22526 21304
rect 22925 21301 22937 21304
rect 22971 21301 22983 21335
rect 22925 21295 22983 21301
rect 24857 21335 24915 21341
rect 24857 21301 24869 21335
rect 24903 21332 24915 21335
rect 25314 21332 25320 21344
rect 24903 21304 25320 21332
rect 24903 21301 24915 21304
rect 24857 21295 24915 21301
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 27264 21332 27292 21431
rect 27430 21428 27436 21480
rect 27488 21468 27494 21480
rect 27525 21471 27583 21477
rect 27525 21468 27537 21471
rect 27488 21440 27537 21468
rect 27488 21428 27494 21440
rect 27525 21437 27537 21440
rect 27571 21437 27583 21471
rect 27525 21431 27583 21437
rect 28350 21428 28356 21480
rect 28408 21468 28414 21480
rect 28813 21471 28871 21477
rect 28813 21468 28825 21471
rect 28408 21440 28825 21468
rect 28408 21428 28414 21440
rect 28813 21437 28825 21440
rect 28859 21468 28871 21471
rect 30009 21471 30067 21477
rect 30009 21468 30021 21471
rect 28859 21440 30021 21468
rect 28859 21437 28871 21440
rect 28813 21431 28871 21437
rect 30009 21437 30021 21440
rect 30055 21437 30067 21471
rect 30009 21431 30067 21437
rect 29270 21400 29276 21412
rect 28736 21372 29276 21400
rect 28736 21332 28764 21372
rect 29270 21360 29276 21372
rect 29328 21360 29334 21412
rect 29365 21403 29423 21409
rect 29365 21369 29377 21403
rect 29411 21369 29423 21403
rect 29365 21363 29423 21369
rect 27264 21304 28764 21332
rect 28810 21292 28816 21344
rect 28868 21332 28874 21344
rect 29380 21332 29408 21363
rect 28868 21304 29408 21332
rect 28868 21292 28874 21304
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1118 21088 1124 21140
rect 1176 21128 1182 21140
rect 1176 21100 4016 21128
rect 1176 21088 1182 21100
rect 3326 21060 3332 21072
rect 3287 21032 3332 21060
rect 3326 21020 3332 21032
rect 3384 21020 3390 21072
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 1854 20992 1860 21004
rect 1627 20964 1860 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 3988 20933 4016 21100
rect 5350 21088 5356 21140
rect 5408 21128 5414 21140
rect 5408 21100 8340 21128
rect 5408 21088 5414 21100
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 4893 20995 4951 21001
rect 4893 20992 4905 20995
rect 4120 20964 4905 20992
rect 4120 20952 4126 20964
rect 4893 20961 4905 20964
rect 4939 20961 4951 20995
rect 4893 20955 4951 20961
rect 6362 20952 6368 21004
rect 6420 20952 6426 21004
rect 6454 20952 6460 21004
rect 6512 20992 6518 21004
rect 7561 20995 7619 21001
rect 7561 20992 7573 20995
rect 6512 20964 7573 20992
rect 6512 20952 6518 20964
rect 7561 20961 7573 20964
rect 7607 20992 7619 20995
rect 8202 20992 8208 21004
rect 7607 20964 8208 20992
rect 7607 20961 7619 20964
rect 7561 20955 7619 20961
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 8312 20992 8340 21100
rect 8386 21088 8392 21140
rect 8444 21128 8450 21140
rect 8444 21100 12388 21128
rect 8444 21088 8450 21100
rect 9122 21020 9128 21072
rect 9180 21060 9186 21072
rect 10410 21060 10416 21072
rect 9180 21032 10416 21060
rect 9180 21020 9186 21032
rect 10410 21020 10416 21032
rect 10468 21020 10474 21072
rect 12360 21060 12388 21100
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 12713 21131 12771 21137
rect 12713 21128 12725 21131
rect 12492 21100 12725 21128
rect 12492 21088 12498 21100
rect 12713 21097 12725 21100
rect 12759 21128 12771 21131
rect 16298 21128 16304 21140
rect 12759 21100 16304 21128
rect 12759 21097 12771 21100
rect 12713 21091 12771 21097
rect 16298 21088 16304 21100
rect 16356 21088 16362 21140
rect 16393 21131 16451 21137
rect 16393 21097 16405 21131
rect 16439 21128 16451 21131
rect 16574 21128 16580 21140
rect 16439 21100 16580 21128
rect 16439 21097 16451 21100
rect 16393 21091 16451 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 16684 21100 20208 21128
rect 12360 21032 12848 21060
rect 10229 20995 10287 21001
rect 8312 20964 10088 20992
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20893 4031 20927
rect 6380 20924 6408 20952
rect 8662 20924 8668 20936
rect 6302 20896 6408 20924
rect 8496 20896 8668 20924
rect 3973 20887 4031 20893
rect 1857 20859 1915 20865
rect 1857 20825 1869 20859
rect 1903 20825 1915 20859
rect 3786 20856 3792 20868
rect 3082 20828 3792 20856
rect 1857 20819 1915 20825
rect 1872 20788 1900 20819
rect 3786 20816 3792 20828
rect 3844 20816 3850 20868
rect 5074 20816 5080 20868
rect 5132 20856 5138 20868
rect 5169 20859 5227 20865
rect 5169 20856 5181 20859
rect 5132 20828 5181 20856
rect 5132 20816 5138 20828
rect 5169 20825 5181 20828
rect 5215 20825 5227 20859
rect 5169 20819 5227 20825
rect 6546 20816 6552 20868
rect 6604 20856 6610 20868
rect 6917 20859 6975 20865
rect 6917 20856 6929 20859
rect 6604 20828 6929 20856
rect 6604 20816 6610 20828
rect 6917 20825 6929 20828
rect 6963 20856 6975 20859
rect 7006 20856 7012 20868
rect 6963 20828 7012 20856
rect 6963 20825 6975 20828
rect 6917 20819 6975 20825
rect 7006 20816 7012 20828
rect 7064 20816 7070 20868
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 7653 20859 7711 20865
rect 7653 20856 7665 20859
rect 7616 20828 7665 20856
rect 7616 20816 7622 20828
rect 7653 20825 7665 20828
rect 7699 20825 7711 20859
rect 8496 20856 8524 20896
rect 8662 20884 8668 20896
rect 8720 20884 8726 20936
rect 10060 20924 10088 20964
rect 10229 20961 10241 20995
rect 10275 20992 10287 20995
rect 10318 20992 10324 21004
rect 10275 20964 10324 20992
rect 10275 20961 10287 20964
rect 10229 20955 10287 20961
rect 10318 20952 10324 20964
rect 10376 20952 10382 21004
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20992 11299 20995
rect 11287 20964 12572 20992
rect 11287 20961 11299 20964
rect 11241 20955 11299 20961
rect 12544 20936 12572 20964
rect 10594 20924 10600 20936
rect 10060 20896 10600 20924
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10962 20924 10968 20936
rect 10923 20896 10968 20924
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 12526 20884 12532 20936
rect 12584 20884 12590 20936
rect 12820 20924 12848 21032
rect 13722 21020 13728 21072
rect 13780 21060 13786 21072
rect 16684 21060 16712 21100
rect 17126 21060 17132 21072
rect 13780 21032 16712 21060
rect 16776 21032 17132 21060
rect 13780 21020 13786 21032
rect 13630 20952 13636 21004
rect 13688 20992 13694 21004
rect 16776 20992 16804 21032
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 18690 21020 18696 21072
rect 18748 21020 18754 21072
rect 18785 21063 18843 21069
rect 18785 21029 18797 21063
rect 18831 21060 18843 21063
rect 19334 21060 19340 21072
rect 18831 21032 19340 21060
rect 18831 21029 18843 21032
rect 18785 21023 18843 21029
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 19426 21020 19432 21072
rect 19484 21060 19490 21072
rect 20180 21060 20208 21100
rect 20530 21088 20536 21140
rect 20588 21128 20594 21140
rect 21450 21128 21456 21140
rect 20588 21100 21456 21128
rect 20588 21088 20594 21100
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 25498 21128 25504 21140
rect 22244 21100 25504 21128
rect 22244 21088 22250 21100
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 28810 21128 28816 21140
rect 25792 21100 28816 21128
rect 25792 21072 25820 21100
rect 28810 21088 28816 21100
rect 28868 21088 28874 21140
rect 29362 21088 29368 21140
rect 29420 21128 29426 21140
rect 29825 21131 29883 21137
rect 29825 21128 29837 21131
rect 29420 21100 29837 21128
rect 29420 21088 29426 21100
rect 29825 21097 29837 21100
rect 29871 21097 29883 21131
rect 29825 21091 29883 21097
rect 19484 21032 20116 21060
rect 20180 21032 23520 21060
rect 19484 21020 19490 21032
rect 18506 20992 18512 21004
rect 13688 20964 16804 20992
rect 16868 20964 18512 20992
rect 13688 20952 13694 20964
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 12820 20896 13553 20924
rect 13541 20893 13553 20896
rect 13587 20924 13599 20927
rect 13722 20924 13728 20936
rect 13587 20896 13728 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 15470 20884 15476 20936
rect 15528 20924 15534 20936
rect 16114 20924 16120 20936
rect 15528 20896 16120 20924
rect 15528 20884 15534 20896
rect 16114 20884 16120 20896
rect 16172 20924 16178 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 16172 20896 16313 20924
rect 16172 20884 16178 20896
rect 16301 20893 16313 20896
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 16390 20884 16396 20936
rect 16448 20924 16454 20936
rect 16868 20924 16896 20964
rect 18506 20952 18512 20964
rect 18564 20952 18570 21004
rect 18708 20992 18736 21020
rect 19521 20995 19579 21001
rect 18708 20964 18828 20992
rect 16448 20896 16896 20924
rect 16448 20884 16454 20896
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18012 20896 18705 20924
rect 18012 20884 18018 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 7653 20819 7711 20825
rect 8036 20828 8524 20856
rect 8573 20859 8631 20865
rect 2774 20788 2780 20800
rect 1872 20760 2780 20788
rect 2774 20748 2780 20760
rect 2832 20748 2838 20800
rect 3970 20748 3976 20800
rect 4028 20788 4034 20800
rect 4157 20791 4215 20797
rect 4157 20788 4169 20791
rect 4028 20760 4169 20788
rect 4028 20748 4034 20760
rect 4157 20757 4169 20760
rect 4203 20757 4215 20791
rect 7024 20788 7052 20816
rect 8036 20788 8064 20828
rect 8573 20825 8585 20859
rect 8619 20856 8631 20859
rect 8846 20856 8852 20868
rect 8619 20828 8852 20856
rect 8619 20825 8631 20828
rect 8573 20819 8631 20825
rect 8846 20816 8852 20828
rect 8904 20856 8910 20868
rect 9030 20856 9036 20868
rect 8904 20828 9036 20856
rect 8904 20816 8910 20828
rect 9030 20816 9036 20828
rect 9088 20816 9094 20868
rect 9214 20856 9220 20868
rect 9175 20828 9220 20856
rect 9214 20816 9220 20828
rect 9272 20816 9278 20868
rect 9309 20859 9367 20865
rect 9309 20825 9321 20859
rect 9355 20825 9367 20859
rect 9309 20819 9367 20825
rect 7024 20760 8064 20788
rect 4157 20751 4215 20757
rect 8110 20748 8116 20800
rect 8168 20788 8174 20800
rect 9324 20788 9352 20819
rect 10318 20816 10324 20868
rect 10376 20856 10382 20868
rect 11146 20856 11152 20868
rect 10376 20828 11152 20856
rect 10376 20816 10382 20828
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 11698 20816 11704 20868
rect 11756 20816 11762 20868
rect 12710 20816 12716 20868
rect 12768 20856 12774 20868
rect 12768 20828 14136 20856
rect 12768 20816 12774 20828
rect 8168 20760 9352 20788
rect 8168 20748 8174 20760
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 9950 20788 9956 20800
rect 9824 20760 9956 20788
rect 9824 20748 9830 20760
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 10870 20788 10876 20800
rect 10100 20760 10876 20788
rect 10100 20748 10106 20760
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 11422 20748 11428 20800
rect 11480 20788 11486 20800
rect 12526 20788 12532 20800
rect 11480 20760 12532 20788
rect 11480 20748 11486 20760
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 13633 20791 13691 20797
rect 13633 20788 13645 20791
rect 13136 20760 13645 20788
rect 13136 20748 13142 20760
rect 13633 20757 13645 20760
rect 13679 20757 13691 20791
rect 14108 20788 14136 20828
rect 14182 20816 14188 20868
rect 14240 20856 14246 20868
rect 14369 20859 14427 20865
rect 14369 20856 14381 20859
rect 14240 20828 14381 20856
rect 14240 20816 14246 20828
rect 14369 20825 14381 20828
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 14458 20816 14464 20868
rect 14516 20856 14522 20868
rect 15286 20856 15292 20868
rect 14516 20828 14561 20856
rect 14752 20828 15292 20856
rect 14516 20816 14522 20828
rect 14752 20788 14780 20828
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 15378 20816 15384 20868
rect 15436 20856 15442 20868
rect 15436 20828 15481 20856
rect 15436 20816 15442 20828
rect 16850 20816 16856 20868
rect 16908 20856 16914 20868
rect 17037 20859 17095 20865
rect 17037 20856 17049 20859
rect 16908 20828 17049 20856
rect 16908 20816 16914 20828
rect 17037 20825 17049 20828
rect 17083 20825 17095 20859
rect 17037 20819 17095 20825
rect 17126 20816 17132 20868
rect 17184 20856 17190 20868
rect 17184 20828 17229 20856
rect 17184 20816 17190 20828
rect 17862 20816 17868 20868
rect 17920 20856 17926 20868
rect 18049 20859 18107 20865
rect 18049 20856 18061 20859
rect 17920 20828 18061 20856
rect 17920 20816 17926 20828
rect 18049 20825 18061 20828
rect 18095 20825 18107 20859
rect 18800 20856 18828 20964
rect 19521 20961 19533 20995
rect 19567 20992 19579 20995
rect 19794 20992 19800 21004
rect 19567 20964 19800 20992
rect 19567 20961 19579 20964
rect 19521 20955 19579 20961
rect 19794 20952 19800 20964
rect 19852 20952 19858 21004
rect 20088 20992 20116 21032
rect 20533 20995 20591 21001
rect 20088 20964 20492 20992
rect 20464 20924 20492 20964
rect 20533 20961 20545 20995
rect 20579 20992 20591 20995
rect 20714 20992 20720 21004
rect 20579 20964 20720 20992
rect 20579 20961 20591 20964
rect 20533 20955 20591 20961
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 21910 20992 21916 21004
rect 21468 20964 21916 20992
rect 21468 20924 21496 20964
rect 21910 20952 21916 20964
rect 21968 20952 21974 21004
rect 22281 20995 22339 21001
rect 22281 20961 22293 20995
rect 22327 20992 22339 20995
rect 22922 20992 22928 21004
rect 22327 20964 22928 20992
rect 22327 20961 22339 20964
rect 22281 20955 22339 20961
rect 22922 20952 22928 20964
rect 22980 20952 22986 21004
rect 20464 20896 21496 20924
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 22094 20924 22100 20936
rect 21591 20896 22100 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 22094 20884 22100 20896
rect 22152 20884 22158 20936
rect 22189 20927 22247 20933
rect 22189 20893 22201 20927
rect 22235 20924 22247 20927
rect 22554 20924 22560 20936
rect 22235 20896 22560 20924
rect 22235 20893 22247 20896
rect 22189 20887 22247 20893
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 22830 20924 22836 20936
rect 22791 20896 22836 20924
rect 22830 20884 22836 20896
rect 22888 20884 22894 20936
rect 23492 20933 23520 21032
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 24486 21060 24492 21072
rect 23900 21032 24492 21060
rect 23900 21020 23906 21032
rect 24486 21020 24492 21032
rect 24544 21020 24550 21072
rect 25774 21060 25780 21072
rect 25687 21032 25780 21060
rect 25774 21020 25780 21032
rect 25832 21020 25838 21072
rect 25958 21020 25964 21072
rect 26016 21060 26022 21072
rect 26016 21032 28580 21060
rect 26016 21020 26022 21032
rect 25225 20995 25283 21001
rect 25225 20961 25237 20995
rect 25271 20992 25283 20995
rect 27246 20992 27252 21004
rect 25271 20964 27252 20992
rect 25271 20961 25283 20964
rect 25225 20955 25283 20961
rect 27246 20952 27252 20964
rect 27304 20952 27310 21004
rect 28552 21001 28580 21032
rect 28537 20995 28595 21001
rect 28537 20961 28549 20995
rect 28583 20961 28595 20995
rect 28537 20955 28595 20961
rect 28626 20952 28632 21004
rect 28684 20992 28690 21004
rect 29638 20992 29644 21004
rect 28684 20964 29644 20992
rect 28684 20952 28690 20964
rect 29638 20952 29644 20964
rect 29696 20952 29702 21004
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 26234 20884 26240 20936
rect 26292 20924 26298 20936
rect 26329 20927 26387 20933
rect 26329 20924 26341 20927
rect 26292 20896 26341 20924
rect 26292 20884 26298 20896
rect 26329 20893 26341 20896
rect 26375 20893 26387 20927
rect 27798 20924 27804 20936
rect 27759 20896 27804 20924
rect 26329 20887 26387 20893
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 29730 20924 29736 20936
rect 29691 20896 29736 20924
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 18800 20828 19288 20856
rect 18049 20819 18107 20825
rect 14108 20760 14780 20788
rect 13633 20751 13691 20757
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 19150 20788 19156 20800
rect 14884 20760 19156 20788
rect 14884 20748 14890 20760
rect 19150 20748 19156 20760
rect 19208 20748 19214 20800
rect 19260 20788 19288 20828
rect 19518 20816 19524 20868
rect 19576 20856 19582 20868
rect 19613 20859 19671 20865
rect 19613 20856 19625 20859
rect 19576 20828 19625 20856
rect 19576 20816 19582 20828
rect 19613 20825 19625 20828
rect 19659 20825 19671 20859
rect 19613 20819 19671 20825
rect 19794 20816 19800 20868
rect 19852 20856 19858 20868
rect 20346 20856 20352 20868
rect 19852 20828 20352 20856
rect 19852 20816 19858 20828
rect 20346 20816 20352 20828
rect 20404 20816 20410 20868
rect 23014 20816 23020 20868
rect 23072 20856 23078 20868
rect 24854 20856 24860 20868
rect 23072 20828 24860 20856
rect 23072 20816 23078 20828
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 25314 20816 25320 20868
rect 25372 20856 25378 20868
rect 25372 20828 25417 20856
rect 25372 20816 25378 20828
rect 25958 20816 25964 20868
rect 26016 20856 26022 20868
rect 26421 20859 26479 20865
rect 26421 20856 26433 20859
rect 26016 20828 26433 20856
rect 26016 20816 26022 20828
rect 26421 20825 26433 20828
rect 26467 20825 26479 20859
rect 26421 20819 26479 20825
rect 28629 20859 28687 20865
rect 28629 20825 28641 20859
rect 28675 20825 28687 20859
rect 28629 20819 28687 20825
rect 29181 20859 29239 20865
rect 29181 20825 29193 20859
rect 29227 20856 29239 20859
rect 30374 20856 30380 20868
rect 29227 20828 30380 20856
rect 29227 20825 29239 20828
rect 29181 20819 29239 20825
rect 21450 20788 21456 20800
rect 19260 20760 21456 20788
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 21637 20791 21695 20797
rect 21637 20757 21649 20791
rect 21683 20788 21695 20791
rect 22186 20788 22192 20800
rect 21683 20760 22192 20788
rect 21683 20757 21695 20760
rect 21637 20751 21695 20757
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 22370 20748 22376 20800
rect 22428 20788 22434 20800
rect 22925 20791 22983 20797
rect 22925 20788 22937 20791
rect 22428 20760 22937 20788
rect 22428 20748 22434 20760
rect 22925 20757 22937 20760
rect 22971 20757 22983 20791
rect 22925 20751 22983 20757
rect 23569 20791 23627 20797
rect 23569 20757 23581 20791
rect 23615 20788 23627 20791
rect 24762 20788 24768 20800
rect 23615 20760 24768 20788
rect 23615 20757 23627 20760
rect 23569 20751 23627 20757
rect 24762 20748 24768 20760
rect 24820 20748 24826 20800
rect 27893 20791 27951 20797
rect 27893 20757 27905 20791
rect 27939 20788 27951 20791
rect 28644 20788 28672 20819
rect 30374 20816 30380 20828
rect 30432 20816 30438 20868
rect 27939 20760 28672 20788
rect 27939 20757 27951 20760
rect 27893 20751 27951 20757
rect 29270 20748 29276 20800
rect 29328 20788 29334 20800
rect 29546 20788 29552 20800
rect 29328 20760 29552 20788
rect 29328 20748 29334 20760
rect 29546 20748 29552 20760
rect 29604 20748 29610 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1210 20544 1216 20596
rect 1268 20584 1274 20596
rect 1268 20556 4016 20584
rect 1268 20544 1274 20556
rect 3878 20516 3884 20528
rect 3358 20488 3884 20516
rect 3878 20476 3884 20488
rect 3936 20476 3942 20528
rect 1854 20448 1860 20460
rect 1815 20420 1860 20448
rect 1854 20408 1860 20420
rect 1912 20408 1918 20460
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20380 2191 20383
rect 3326 20380 3332 20392
rect 2179 20352 3332 20380
rect 2179 20349 2191 20352
rect 2133 20343 2191 20349
rect 3326 20340 3332 20352
rect 3384 20340 3390 20392
rect 3878 20380 3884 20392
rect 3839 20352 3884 20380
rect 3878 20340 3884 20352
rect 3936 20340 3942 20392
rect 3988 20380 4016 20556
rect 4062 20544 4068 20596
rect 4120 20584 4126 20596
rect 4120 20556 6684 20584
rect 4120 20544 4126 20556
rect 4982 20516 4988 20528
rect 4943 20488 4988 20516
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 5077 20519 5135 20525
rect 5077 20485 5089 20519
rect 5123 20516 5135 20519
rect 5442 20516 5448 20528
rect 5123 20488 5448 20516
rect 5123 20485 5135 20488
rect 5077 20479 5135 20485
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 6656 20525 6684 20556
rect 6748 20556 9996 20584
rect 6641 20519 6699 20525
rect 6641 20485 6653 20519
rect 6687 20485 6699 20519
rect 6641 20479 6699 20485
rect 6748 20448 6776 20556
rect 7190 20476 7196 20528
rect 7248 20516 7254 20528
rect 7653 20519 7711 20525
rect 7653 20516 7665 20519
rect 7248 20488 7665 20516
rect 7248 20476 7254 20488
rect 7653 20485 7665 20488
rect 7699 20485 7711 20519
rect 9398 20516 9404 20528
rect 8878 20488 9404 20516
rect 7653 20479 7711 20485
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 9968 20525 9996 20556
rect 10226 20544 10232 20596
rect 10284 20584 10290 20596
rect 12894 20584 12900 20596
rect 10284 20556 12900 20584
rect 10284 20544 10290 20556
rect 12894 20544 12900 20556
rect 12952 20544 12958 20596
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 14826 20584 14832 20596
rect 14691 20556 14832 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15344 20556 15516 20584
rect 15344 20544 15350 20556
rect 9953 20519 10011 20525
rect 9953 20485 9965 20519
rect 9999 20485 10011 20519
rect 9953 20479 10011 20485
rect 10778 20476 10784 20528
rect 10836 20516 10842 20528
rect 10873 20519 10931 20525
rect 10873 20516 10885 20519
rect 10836 20488 10885 20516
rect 10836 20476 10842 20488
rect 10873 20485 10885 20488
rect 10919 20516 10931 20519
rect 11974 20516 11980 20528
rect 10919 20488 11980 20516
rect 10919 20485 10931 20488
rect 10873 20479 10931 20485
rect 11974 20476 11980 20488
rect 12032 20476 12038 20528
rect 13354 20516 13360 20528
rect 13202 20488 13360 20516
rect 13354 20476 13360 20488
rect 13412 20476 13418 20528
rect 13446 20476 13452 20528
rect 13504 20516 13510 20528
rect 13725 20519 13783 20525
rect 13725 20516 13737 20519
rect 13504 20488 13737 20516
rect 13504 20476 13510 20488
rect 13725 20485 13737 20488
rect 13771 20485 13783 20519
rect 13725 20479 13783 20485
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 15381 20519 15439 20525
rect 15381 20516 15393 20519
rect 13964 20488 15393 20516
rect 13964 20476 13970 20488
rect 15381 20485 15393 20488
rect 15427 20485 15439 20519
rect 15488 20516 15516 20556
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 17126 20584 17132 20596
rect 16632 20556 17132 20584
rect 16632 20544 16638 20556
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 17405 20587 17463 20593
rect 17405 20553 17417 20587
rect 17451 20553 17463 20587
rect 17405 20547 17463 20553
rect 17420 20516 17448 20547
rect 18690 20544 18696 20596
rect 18748 20584 18754 20596
rect 19242 20584 19248 20596
rect 18748 20556 19248 20584
rect 18748 20544 18754 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19886 20584 19892 20596
rect 19484 20556 19892 20584
rect 19484 20544 19490 20556
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 25041 20587 25099 20593
rect 25041 20584 25053 20587
rect 20180 20556 25053 20584
rect 18782 20516 18788 20528
rect 15488 20488 17448 20516
rect 18743 20488 18788 20516
rect 15381 20479 15439 20485
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 19705 20519 19763 20525
rect 19705 20485 19717 20519
rect 19751 20516 19763 20519
rect 20070 20516 20076 20528
rect 19751 20488 20076 20516
rect 19751 20485 19763 20488
rect 19705 20479 19763 20485
rect 20070 20476 20076 20488
rect 20128 20476 20134 20528
rect 5828 20420 6776 20448
rect 5828 20380 5856 20420
rect 6914 20408 6920 20460
rect 6972 20448 6978 20460
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 6972 20420 7389 20448
rect 6972 20408 6978 20420
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 9214 20448 9220 20460
rect 7377 20411 7435 20417
rect 8864 20420 9220 20448
rect 3988 20352 5856 20380
rect 5997 20383 6055 20389
rect 5997 20349 6009 20383
rect 6043 20380 6055 20383
rect 7282 20380 7288 20392
rect 6043 20352 7288 20380
rect 6043 20349 6055 20352
rect 5997 20343 6055 20349
rect 7282 20340 7288 20352
rect 7340 20340 7346 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 8864 20380 8892 20420
rect 9214 20408 9220 20420
rect 9272 20408 9278 20460
rect 9493 20451 9551 20457
rect 9493 20417 9505 20451
rect 9539 20448 9551 20451
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 9539 20420 9720 20448
rect 9539 20417 9551 20420
rect 9493 20411 9551 20417
rect 8352 20352 8892 20380
rect 9125 20383 9183 20389
rect 8352 20340 8358 20352
rect 9125 20349 9137 20383
rect 9171 20380 9183 20383
rect 9692 20380 9720 20420
rect 13188 20420 14565 20448
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9171 20352 9628 20380
rect 9692 20352 9873 20380
rect 9171 20349 9183 20352
rect 9125 20343 9183 20349
rect 3510 20272 3516 20324
rect 3568 20312 3574 20324
rect 9600 20312 9628 20352
rect 9861 20349 9873 20352
rect 9907 20380 9919 20383
rect 9950 20380 9956 20392
rect 9907 20352 9956 20380
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 9950 20340 9956 20352
rect 10008 20340 10014 20392
rect 10962 20340 10968 20392
rect 11020 20380 11026 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 11020 20352 11713 20380
rect 11020 20340 11026 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 11964 20383 12022 20389
rect 11964 20349 11976 20383
rect 12010 20380 12022 20383
rect 12066 20380 12072 20392
rect 12010 20352 12072 20380
rect 12010 20349 12022 20352
rect 11964 20343 12022 20349
rect 12066 20340 12072 20352
rect 12124 20340 12130 20392
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 13188 20380 13216 20420
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17954 20448 17960 20460
rect 17915 20420 17960 20448
rect 17313 20411 17371 20417
rect 12584 20352 13216 20380
rect 12584 20340 12590 20352
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14642 20380 14648 20392
rect 13872 20352 14648 20380
rect 13872 20340 13878 20352
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 15286 20380 15292 20392
rect 15247 20352 15292 20380
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 16114 20380 16120 20392
rect 15488 20340 15769 20368
rect 16075 20352 16120 20380
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 17218 20380 17224 20392
rect 16356 20352 17224 20380
rect 16356 20340 16362 20352
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 17336 20380 17364 20411
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 20180 20448 20208 20556
rect 25041 20553 25053 20556
rect 25087 20553 25099 20587
rect 25041 20547 25099 20553
rect 26237 20587 26295 20593
rect 26237 20553 26249 20587
rect 26283 20584 26295 20587
rect 26326 20584 26332 20596
rect 26283 20556 26332 20584
rect 26283 20553 26295 20556
rect 26237 20547 26295 20553
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 28445 20587 28503 20593
rect 28445 20553 28457 20587
rect 28491 20584 28503 20587
rect 28902 20584 28908 20596
rect 28491 20556 28908 20584
rect 28491 20553 28503 20556
rect 28445 20547 28503 20553
rect 28902 20544 28908 20556
rect 28960 20544 28966 20596
rect 20257 20519 20315 20525
rect 20257 20485 20269 20519
rect 20303 20516 20315 20519
rect 20438 20516 20444 20528
rect 20303 20488 20444 20516
rect 20303 20485 20315 20488
rect 20257 20479 20315 20485
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 22370 20516 22376 20528
rect 22331 20488 22376 20516
rect 22370 20476 22376 20488
rect 22428 20476 22434 20528
rect 22462 20476 22468 20528
rect 22520 20516 22526 20528
rect 22520 20488 24900 20516
rect 22520 20476 22526 20488
rect 20901 20451 20959 20457
rect 19668 20420 20208 20448
rect 19668 20408 19674 20420
rect 20346 20398 20352 20450
rect 20404 20438 20410 20450
rect 20640 20438 20760 20448
rect 20404 20420 20760 20438
rect 20404 20410 20668 20420
rect 20404 20398 20410 20410
rect 17494 20380 17500 20392
rect 17336 20352 17500 20380
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 18690 20380 18696 20392
rect 18651 20352 18696 20380
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 18782 20340 18788 20392
rect 18840 20380 18846 20392
rect 20732 20380 20760 20420
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 21726 20448 21732 20460
rect 20947 20420 21732 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 21726 20408 21732 20420
rect 21784 20408 21790 20460
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 23385 20451 23443 20457
rect 23385 20448 23397 20451
rect 23072 20420 23397 20448
rect 23072 20408 23078 20420
rect 23385 20417 23397 20420
rect 23431 20448 23443 20451
rect 23474 20448 23480 20460
rect 23431 20420 23480 20448
rect 23431 20417 23443 20420
rect 23385 20411 23443 20417
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 24118 20448 24124 20460
rect 23768 20420 24124 20448
rect 21174 20380 21180 20392
rect 18840 20352 20208 20380
rect 20732 20352 21180 20380
rect 18840 20340 18846 20352
rect 11606 20312 11612 20324
rect 3568 20284 4016 20312
rect 9600 20284 11612 20312
rect 3568 20272 3574 20284
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 3878 20244 3884 20256
rect 1820 20216 3884 20244
rect 1820 20204 1826 20216
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 3988 20244 4016 20284
rect 11606 20272 11612 20284
rect 11664 20272 11670 20324
rect 5994 20244 6000 20256
rect 3988 20216 6000 20244
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6733 20247 6791 20253
rect 6733 20213 6745 20247
rect 6779 20244 6791 20247
rect 15488 20244 15516 20340
rect 15741 20312 15769 20340
rect 19978 20312 19984 20324
rect 15741 20284 19984 20312
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 20180 20312 20208 20352
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 21818 20340 21824 20392
rect 21876 20380 21882 20392
rect 22002 20380 22008 20392
rect 21876 20352 22008 20380
rect 21876 20340 21882 20352
rect 22002 20340 22008 20352
rect 22060 20340 22066 20392
rect 22278 20380 22284 20392
rect 22239 20352 22284 20380
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 23768 20380 23796 20420
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 24872 20448 24900 20488
rect 26142 20476 26148 20528
rect 26200 20516 26206 20528
rect 27798 20516 27804 20528
rect 26200 20488 27804 20516
rect 26200 20476 26206 20488
rect 27798 20476 27804 20488
rect 27856 20476 27862 20528
rect 27890 20476 27896 20528
rect 27948 20516 27954 20528
rect 29454 20516 29460 20528
rect 27948 20488 29460 20516
rect 27948 20476 27954 20488
rect 29454 20476 29460 20488
rect 29512 20476 29518 20528
rect 24949 20451 25007 20457
rect 24949 20448 24961 20451
rect 24872 20420 24961 20448
rect 24949 20417 24961 20420
rect 24995 20417 25007 20451
rect 24949 20411 25007 20417
rect 25593 20451 25651 20457
rect 25593 20417 25605 20451
rect 25639 20417 25651 20451
rect 25593 20411 25651 20417
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20417 26479 20451
rect 26421 20411 26479 20417
rect 22388 20352 23796 20380
rect 22388 20312 22416 20352
rect 23842 20340 23848 20392
rect 23900 20380 23906 20392
rect 25608 20380 25636 20411
rect 23900 20352 25636 20380
rect 23900 20340 23906 20352
rect 25682 20340 25688 20392
rect 25740 20380 25746 20392
rect 25740 20352 25785 20380
rect 25740 20340 25746 20352
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26436 20380 26464 20411
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 27120 20420 27169 20448
rect 27120 20408 27126 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27816 20448 27844 20476
rect 28353 20451 28411 20457
rect 28353 20448 28365 20451
rect 27816 20420 28365 20448
rect 27157 20411 27215 20417
rect 28353 20417 28365 20420
rect 28399 20417 28411 20451
rect 28994 20448 29000 20460
rect 28955 20420 29000 20448
rect 28353 20411 28411 20417
rect 28994 20408 29000 20420
rect 29052 20448 29058 20460
rect 29641 20451 29699 20457
rect 29641 20448 29653 20451
rect 29052 20420 29653 20448
rect 29052 20408 29058 20420
rect 29641 20417 29653 20420
rect 29687 20448 29699 20451
rect 29730 20448 29736 20460
rect 29687 20420 29736 20448
rect 29687 20417 29699 20420
rect 29641 20411 29699 20417
rect 29730 20408 29736 20420
rect 29788 20408 29794 20460
rect 28442 20380 28448 20392
rect 26016 20352 28448 20380
rect 26016 20340 26022 20352
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 22830 20312 22836 20324
rect 20180 20284 22416 20312
rect 22791 20284 22836 20312
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 22922 20272 22928 20324
rect 22980 20312 22986 20324
rect 25774 20312 25780 20324
rect 22980 20284 25780 20312
rect 22980 20272 22986 20284
rect 25774 20272 25780 20284
rect 25832 20272 25838 20324
rect 27249 20315 27307 20321
rect 27249 20281 27261 20315
rect 27295 20312 27307 20315
rect 30006 20312 30012 20324
rect 27295 20284 30012 20312
rect 27295 20281 27307 20284
rect 27249 20275 27307 20281
rect 30006 20272 30012 20284
rect 30064 20272 30070 20324
rect 6779 20216 15516 20244
rect 6779 20213 6791 20216
rect 6733 20207 6791 20213
rect 15838 20204 15844 20256
rect 15896 20244 15902 20256
rect 17862 20244 17868 20256
rect 15896 20216 17868 20244
rect 15896 20204 15902 20216
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 18012 20216 18061 20244
rect 18012 20204 18018 20216
rect 18049 20213 18061 20216
rect 18095 20213 18107 20247
rect 18049 20207 18107 20213
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 19058 20244 19064 20256
rect 18564 20216 19064 20244
rect 18564 20204 18570 20216
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19242 20204 19248 20256
rect 19300 20244 19306 20256
rect 20349 20247 20407 20253
rect 20349 20244 20361 20247
rect 19300 20216 20361 20244
rect 19300 20204 19306 20216
rect 20349 20213 20361 20216
rect 20395 20213 20407 20247
rect 20349 20207 20407 20213
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 20993 20247 21051 20253
rect 20993 20244 21005 20247
rect 20772 20216 21005 20244
rect 20772 20204 20778 20216
rect 20993 20213 21005 20216
rect 21039 20213 21051 20247
rect 20993 20207 21051 20213
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 23014 20244 23020 20256
rect 21324 20216 23020 20244
rect 21324 20204 21330 20216
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 23474 20244 23480 20256
rect 23435 20216 23480 20244
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 24397 20247 24455 20253
rect 24397 20244 24409 20247
rect 24360 20216 24409 20244
rect 24360 20204 24366 20216
rect 24397 20213 24409 20216
rect 24443 20213 24455 20247
rect 24397 20207 24455 20213
rect 24486 20204 24492 20256
rect 24544 20244 24550 20256
rect 27062 20244 27068 20256
rect 24544 20216 27068 20244
rect 24544 20204 24550 20216
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 27338 20204 27344 20256
rect 27396 20244 27402 20256
rect 29089 20247 29147 20253
rect 29089 20244 29101 20247
rect 27396 20216 29101 20244
rect 27396 20204 27402 20216
rect 29089 20213 29101 20216
rect 29135 20213 29147 20247
rect 29730 20244 29736 20256
rect 29691 20216 29736 20244
rect 29089 20207 29147 20213
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1844 20043 1902 20049
rect 1844 20009 1856 20043
rect 1890 20040 1902 20043
rect 2958 20040 2964 20052
rect 1890 20012 2964 20040
rect 1890 20009 1902 20012
rect 1844 20003 1902 20009
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 3329 20043 3387 20049
rect 3329 20009 3341 20043
rect 3375 20040 3387 20043
rect 3694 20040 3700 20052
rect 3375 20012 3700 20040
rect 3375 20009 3387 20012
rect 3329 20003 3387 20009
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 8481 20043 8539 20049
rect 3936 20012 7236 20040
rect 3936 20000 3942 20012
rect 7208 19972 7236 20012
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 11698 20040 11704 20052
rect 8527 20012 11704 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 11698 20000 11704 20012
rect 11756 20000 11762 20052
rect 12894 20040 12900 20052
rect 12268 20012 12900 20040
rect 12268 19972 12296 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13630 20040 13636 20052
rect 13591 20012 13636 20040
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 16758 20040 16764 20052
rect 13964 20012 16764 20040
rect 13964 20000 13970 20012
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 18782 20040 18788 20052
rect 17000 20012 18788 20040
rect 17000 20000 17006 20012
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 19610 20040 19616 20052
rect 18932 20012 19616 20040
rect 18932 20000 18938 20012
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 21082 20040 21088 20052
rect 19713 20012 20953 20040
rect 21043 20012 21088 20040
rect 12434 19972 12440 19984
rect 7208 19944 11008 19972
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19904 1639 19907
rect 1854 19904 1860 19916
rect 1627 19876 1860 19904
rect 1627 19873 1639 19876
rect 1581 19867 1639 19873
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 2866 19864 2872 19916
rect 2924 19904 2930 19916
rect 3418 19904 3424 19916
rect 2924 19876 3424 19904
rect 2924 19864 2930 19876
rect 3418 19864 3424 19876
rect 3476 19904 3482 19916
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3476 19876 4077 19904
rect 3476 19864 3482 19876
rect 4065 19873 4077 19876
rect 4111 19904 4123 19907
rect 5350 19904 5356 19916
rect 4111 19876 5356 19904
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 5350 19864 5356 19876
rect 5408 19864 5414 19916
rect 5905 19907 5963 19913
rect 5905 19873 5917 19907
rect 5951 19904 5963 19907
rect 6914 19904 6920 19916
rect 5951 19876 6920 19904
rect 5951 19873 5963 19876
rect 5905 19867 5963 19873
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 10226 19904 10232 19916
rect 9272 19876 10088 19904
rect 10187 19876 10232 19904
rect 9272 19864 9278 19876
rect 8386 19836 8392 19848
rect 8347 19808 8392 19836
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 10060 19836 10088 19876
rect 10226 19864 10232 19876
rect 10284 19864 10290 19916
rect 10870 19904 10876 19916
rect 10831 19876 10876 19904
rect 10870 19864 10876 19876
rect 10928 19864 10934 19916
rect 10980 19904 11008 19944
rect 12177 19944 12296 19972
rect 12360 19944 12440 19972
rect 12177 19904 12205 19944
rect 12360 19904 12388 19944
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 12526 19932 12532 19984
rect 12584 19972 12590 19984
rect 18141 19975 18199 19981
rect 18141 19972 18153 19975
rect 12584 19944 18153 19972
rect 12584 19932 12590 19944
rect 18141 19941 18153 19944
rect 18187 19941 18199 19975
rect 19426 19972 19432 19984
rect 18141 19935 18199 19941
rect 18524 19944 19432 19972
rect 10980 19876 12205 19904
rect 12268 19876 12388 19904
rect 10594 19836 10600 19848
rect 10060 19808 10600 19836
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 12268 19822 12296 19876
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 16942 19904 16948 19916
rect 12768 19876 16948 19904
rect 12768 19864 12774 19876
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17037 19907 17095 19913
rect 17037 19873 17049 19907
rect 17083 19904 17095 19907
rect 17310 19904 17316 19916
rect 17083 19876 17316 19904
rect 17083 19873 17095 19876
rect 17037 19867 17095 19873
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 18524 19904 18552 19944
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 19713 19972 19741 20012
rect 19536 19944 19741 19972
rect 19536 19913 19564 19944
rect 19886 19932 19892 19984
rect 19944 19972 19950 19984
rect 20346 19972 20352 19984
rect 19944 19944 20352 19972
rect 19944 19932 19950 19944
rect 20346 19932 20352 19944
rect 20404 19972 20410 19984
rect 20806 19972 20812 19984
rect 20404 19944 20812 19972
rect 20404 19932 20410 19944
rect 20806 19932 20812 19944
rect 20864 19932 20870 19984
rect 20925 19972 20953 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 23382 20040 23388 20052
rect 22520 20012 23388 20040
rect 22520 20000 22526 20012
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 23716 20012 23761 20040
rect 23716 20000 23722 20012
rect 24302 19972 24308 19984
rect 20925 19944 24308 19972
rect 24302 19932 24308 19944
rect 24360 19972 24366 19984
rect 25590 19972 25596 19984
rect 24360 19944 25596 19972
rect 24360 19932 24366 19944
rect 25590 19932 25596 19944
rect 25648 19932 25654 19984
rect 27706 19972 27712 19984
rect 27667 19944 27712 19972
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 17420 19876 18552 19904
rect 19521 19907 19579 19913
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 13722 19836 13728 19848
rect 13596 19808 13728 19836
rect 13596 19796 13602 19808
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 17420 19836 17448 19876
rect 19521 19873 19533 19907
rect 19567 19873 19579 19907
rect 19521 19867 19579 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19797 19907 19855 19913
rect 19797 19904 19809 19907
rect 19668 19876 19809 19904
rect 19668 19864 19674 19876
rect 19797 19873 19809 19876
rect 19843 19904 19855 19907
rect 20070 19904 20076 19916
rect 19843 19876 20076 19904
rect 19843 19873 19855 19876
rect 19797 19867 19855 19873
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 25682 19904 25688 19916
rect 20464 19876 25688 19904
rect 17336 19808 17448 19836
rect 2590 19728 2596 19780
rect 2648 19728 2654 19780
rect 4157 19771 4215 19777
rect 3252 19740 3464 19768
rect 2682 19660 2688 19712
rect 2740 19700 2746 19712
rect 3252 19700 3280 19740
rect 2740 19672 3280 19700
rect 3436 19700 3464 19740
rect 4157 19737 4169 19771
rect 4203 19737 4215 19771
rect 4157 19731 4215 19737
rect 4172 19700 4200 19731
rect 4614 19728 4620 19780
rect 4672 19768 4678 19780
rect 5077 19771 5135 19777
rect 5077 19768 5089 19771
rect 4672 19740 5089 19768
rect 4672 19728 4678 19740
rect 5077 19737 5089 19740
rect 5123 19768 5135 19771
rect 5442 19768 5448 19780
rect 5123 19740 5448 19768
rect 5123 19737 5135 19740
rect 5077 19731 5135 19737
rect 5442 19728 5448 19740
rect 5500 19728 5506 19780
rect 5810 19728 5816 19780
rect 5868 19768 5874 19780
rect 6181 19771 6239 19777
rect 6181 19768 6193 19771
rect 5868 19740 6193 19768
rect 5868 19728 5874 19740
rect 6181 19737 6193 19740
rect 6227 19737 6239 19771
rect 7834 19768 7840 19780
rect 7406 19740 7840 19768
rect 6181 19731 6239 19737
rect 7834 19728 7840 19740
rect 7892 19728 7898 19780
rect 9030 19728 9036 19780
rect 9088 19768 9094 19780
rect 9206 19771 9264 19777
rect 9206 19768 9218 19771
rect 9088 19740 9218 19768
rect 9088 19728 9094 19740
rect 9206 19737 9218 19740
rect 9252 19737 9264 19771
rect 9206 19731 9264 19737
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19737 9367 19771
rect 9309 19731 9367 19737
rect 3436 19672 4200 19700
rect 2740 19660 2746 19672
rect 4706 19660 4712 19712
rect 4764 19700 4770 19712
rect 7653 19703 7711 19709
rect 7653 19700 7665 19703
rect 4764 19672 7665 19700
rect 4764 19660 4770 19672
rect 7653 19669 7665 19672
rect 7699 19669 7711 19703
rect 7653 19663 7711 19669
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 9324 19700 9352 19731
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 10870 19768 10876 19780
rect 9456 19740 10876 19768
rect 9456 19728 9462 19740
rect 10870 19728 10876 19740
rect 10928 19728 10934 19780
rect 11149 19771 11207 19777
rect 11149 19737 11161 19771
rect 11195 19768 11207 19771
rect 11238 19768 11244 19780
rect 11195 19740 11244 19768
rect 11195 19737 11207 19740
rect 11149 19731 11207 19737
rect 11238 19728 11244 19740
rect 11296 19728 11302 19780
rect 12710 19768 12716 19780
rect 12452 19740 12716 19768
rect 8720 19672 9352 19700
rect 8720 19660 8726 19672
rect 9490 19660 9496 19712
rect 9548 19700 9554 19712
rect 12452 19700 12480 19740
rect 12710 19728 12716 19740
rect 12768 19728 12774 19780
rect 12897 19771 12955 19777
rect 12897 19737 12909 19771
rect 12943 19768 12955 19771
rect 13354 19768 13360 19780
rect 12943 19740 13360 19768
rect 12943 19737 12955 19740
rect 12897 19731 12955 19737
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 13446 19728 13452 19780
rect 13504 19768 13510 19780
rect 13906 19768 13912 19780
rect 13504 19740 13912 19768
rect 13504 19728 13510 19740
rect 13906 19728 13912 19740
rect 13964 19728 13970 19780
rect 14090 19728 14096 19780
rect 14148 19768 14154 19780
rect 14369 19771 14427 19777
rect 14369 19768 14381 19771
rect 14148 19740 14381 19768
rect 14148 19728 14154 19740
rect 14369 19737 14381 19740
rect 14415 19737 14427 19771
rect 14369 19731 14427 19737
rect 14461 19771 14519 19777
rect 14461 19737 14473 19771
rect 14507 19768 14519 19771
rect 14918 19768 14924 19780
rect 14507 19740 14924 19768
rect 14507 19737 14519 19740
rect 14461 19731 14519 19737
rect 14918 19728 14924 19740
rect 14976 19728 14982 19780
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 15562 19768 15568 19780
rect 15427 19740 15568 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 15562 19728 15568 19740
rect 15620 19728 15626 19780
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 16025 19771 16083 19777
rect 16025 19768 16037 19771
rect 15896 19740 16037 19768
rect 15896 19728 15902 19740
rect 16025 19737 16037 19740
rect 16071 19737 16083 19771
rect 16025 19731 16083 19737
rect 16117 19771 16175 19777
rect 16117 19737 16129 19771
rect 16163 19768 16175 19771
rect 17336 19768 17364 19808
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18472 19808 18705 19836
rect 18472 19796 18478 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 17586 19768 17592 19780
rect 16163 19740 17364 19768
rect 17547 19740 17592 19768
rect 16163 19737 16175 19740
rect 16117 19731 16175 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 17736 19740 17781 19768
rect 17880 19740 18920 19768
rect 17736 19728 17742 19740
rect 9548 19672 12480 19700
rect 9548 19660 9554 19672
rect 12526 19660 12532 19712
rect 12584 19700 12590 19712
rect 13630 19700 13636 19712
rect 12584 19672 13636 19700
rect 12584 19660 12590 19672
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 13722 19660 13728 19712
rect 13780 19700 13786 19712
rect 17880 19700 17908 19740
rect 18782 19700 18788 19712
rect 13780 19672 17908 19700
rect 18743 19672 18788 19700
rect 13780 19660 13786 19672
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 18892 19700 18920 19740
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 19334 19768 19340 19780
rect 19024 19740 19340 19768
rect 19024 19728 19030 19740
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 19622 19771 19680 19777
rect 19622 19737 19634 19771
rect 19668 19768 19680 19771
rect 20464 19768 20492 19876
rect 25682 19864 25688 19876
rect 25740 19864 25746 19916
rect 26418 19864 26424 19916
rect 26476 19904 26482 19916
rect 26476 19876 28948 19904
rect 26476 19864 26482 19876
rect 20898 19796 20904 19848
rect 20956 19836 20962 19848
rect 20993 19839 21051 19845
rect 20993 19836 21005 19839
rect 20956 19808 21005 19836
rect 20956 19796 20962 19808
rect 20993 19805 21005 19808
rect 21039 19805 21051 19839
rect 20993 19799 21051 19805
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 21634 19836 21640 19848
rect 21232 19808 21404 19836
rect 21595 19808 21640 19836
rect 21232 19796 21238 19808
rect 21266 19768 21272 19780
rect 19668 19740 20492 19768
rect 20640 19740 21272 19768
rect 19668 19737 19680 19740
rect 19622 19731 19680 19737
rect 20640 19700 20668 19740
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 21376 19768 21404 19808
rect 21634 19796 21640 19808
rect 21692 19796 21698 19848
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19836 23627 19839
rect 23750 19836 23756 19848
rect 23615 19808 23756 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 24210 19796 24216 19848
rect 24268 19836 24274 19848
rect 24486 19836 24492 19848
rect 24268 19808 24492 19836
rect 24268 19796 24274 19808
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 24581 19839 24639 19845
rect 24581 19805 24593 19839
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 22462 19768 22468 19780
rect 21376 19740 21864 19768
rect 22423 19740 22468 19768
rect 18892 19672 20668 19700
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 21729 19703 21787 19709
rect 21729 19700 21741 19703
rect 21232 19672 21741 19700
rect 21232 19660 21238 19672
rect 21729 19669 21741 19672
rect 21775 19669 21787 19703
rect 21836 19700 21864 19740
rect 22462 19728 22468 19740
rect 22520 19728 22526 19780
rect 22554 19728 22560 19780
rect 22612 19768 22618 19780
rect 22612 19740 22657 19768
rect 22612 19728 22618 19740
rect 22922 19728 22928 19780
rect 22980 19768 22986 19780
rect 23109 19771 23167 19777
rect 23109 19768 23121 19771
rect 22980 19740 23121 19768
rect 22980 19728 22986 19740
rect 23109 19737 23121 19740
rect 23155 19737 23167 19771
rect 23658 19768 23664 19780
rect 23109 19731 23167 19737
rect 23216 19740 23664 19768
rect 23216 19700 23244 19740
rect 23658 19728 23664 19740
rect 23716 19768 23722 19780
rect 24596 19768 24624 19799
rect 25038 19796 25044 19848
rect 25096 19836 25102 19848
rect 26329 19839 26387 19845
rect 26329 19836 26341 19839
rect 25096 19808 26341 19836
rect 25096 19796 25102 19808
rect 26329 19805 26341 19808
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19836 27031 19839
rect 27246 19836 27252 19848
rect 27019 19808 27252 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27246 19796 27252 19808
rect 27304 19836 27310 19848
rect 27617 19839 27675 19845
rect 27617 19836 27629 19839
rect 27304 19808 27629 19836
rect 27304 19796 27310 19808
rect 27617 19805 27629 19808
rect 27663 19805 27675 19839
rect 28258 19836 28264 19848
rect 28219 19808 28264 19836
rect 27617 19799 27675 19805
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 28920 19845 28948 19876
rect 28905 19839 28963 19845
rect 28905 19805 28917 19839
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19836 31079 19839
rect 37826 19836 37832 19848
rect 31067 19808 37832 19836
rect 31067 19805 31079 19808
rect 31021 19799 31079 19805
rect 37826 19796 37832 19808
rect 37884 19796 37890 19848
rect 38286 19836 38292 19848
rect 38247 19808 38292 19836
rect 38286 19796 38292 19808
rect 38344 19796 38350 19848
rect 23716 19740 24624 19768
rect 23716 19728 23722 19740
rect 24854 19728 24860 19780
rect 24912 19768 24918 19780
rect 25685 19771 25743 19777
rect 25685 19768 25697 19771
rect 24912 19740 25697 19768
rect 24912 19728 24918 19740
rect 25685 19737 25697 19740
rect 25731 19737 25743 19771
rect 29914 19768 29920 19780
rect 29875 19740 29920 19768
rect 25685 19731 25743 19737
rect 29914 19728 29920 19740
rect 29972 19728 29978 19780
rect 30006 19728 30012 19780
rect 30064 19768 30070 19780
rect 30064 19740 30109 19768
rect 30064 19728 30070 19740
rect 30374 19728 30380 19780
rect 30432 19768 30438 19780
rect 30561 19771 30619 19777
rect 30561 19768 30573 19771
rect 30432 19740 30573 19768
rect 30432 19728 30438 19740
rect 30561 19737 30573 19740
rect 30607 19768 30619 19771
rect 31386 19768 31392 19780
rect 30607 19740 31392 19768
rect 30607 19737 30619 19740
rect 30561 19731 30619 19737
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 21836 19672 23244 19700
rect 21729 19663 21787 19669
rect 23382 19660 23388 19712
rect 23440 19700 23446 19712
rect 24673 19703 24731 19709
rect 24673 19700 24685 19703
rect 23440 19672 24685 19700
rect 23440 19660 23446 19672
rect 24673 19669 24685 19672
rect 24719 19669 24731 19703
rect 25774 19700 25780 19712
rect 25735 19672 25780 19700
rect 24673 19663 24731 19669
rect 25774 19660 25780 19672
rect 25832 19660 25838 19712
rect 26418 19700 26424 19712
rect 26379 19672 26424 19700
rect 26418 19660 26424 19672
rect 26476 19660 26482 19712
rect 27062 19700 27068 19712
rect 27023 19672 27068 19700
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 28353 19703 28411 19709
rect 28353 19700 28365 19703
rect 27856 19672 28365 19700
rect 27856 19660 27862 19672
rect 28353 19669 28365 19672
rect 28399 19669 28411 19703
rect 28353 19663 28411 19669
rect 28534 19660 28540 19712
rect 28592 19700 28598 19712
rect 28997 19703 29055 19709
rect 28997 19700 29009 19703
rect 28592 19672 29009 19700
rect 28592 19660 28598 19672
rect 28997 19669 29009 19672
rect 29043 19669 29055 19703
rect 28997 19663 29055 19669
rect 29086 19660 29092 19712
rect 29144 19700 29150 19712
rect 31113 19703 31171 19709
rect 31113 19700 31125 19703
rect 29144 19672 31125 19700
rect 29144 19660 29150 19672
rect 31113 19669 31125 19672
rect 31159 19669 31171 19703
rect 31113 19663 31171 19669
rect 31478 19660 31484 19712
rect 31536 19700 31542 19712
rect 38105 19703 38163 19709
rect 38105 19700 38117 19703
rect 31536 19672 38117 19700
rect 31536 19660 31542 19672
rect 38105 19669 38117 19672
rect 38151 19669 38163 19703
rect 38105 19663 38163 19669
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1946 19456 1952 19508
rect 2004 19496 2010 19508
rect 3513 19499 3571 19505
rect 3513 19496 3525 19499
rect 2004 19468 3525 19496
rect 2004 19456 2010 19468
rect 3513 19465 3525 19468
rect 3559 19465 3571 19499
rect 11238 19496 11244 19508
rect 3513 19459 3571 19465
rect 4632 19468 11244 19496
rect 4632 19428 4660 19468
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 13170 19496 13176 19508
rect 12176 19468 13176 19496
rect 3266 19400 4660 19428
rect 5997 19431 6055 19437
rect 5997 19397 6009 19431
rect 6043 19428 6055 19431
rect 6730 19428 6736 19440
rect 6043 19400 6736 19428
rect 6043 19397 6055 19400
rect 5997 19391 6055 19397
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 7742 19428 7748 19440
rect 6840 19400 7748 19428
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 5350 19320 5356 19372
rect 5408 19320 5414 19372
rect 6840 19369 6868 19400
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 9490 19428 9496 19440
rect 9451 19400 9496 19428
rect 9490 19388 9496 19400
rect 9548 19388 9554 19440
rect 10134 19428 10140 19440
rect 10095 19400 10140 19428
rect 10134 19388 10140 19400
rect 10192 19388 10198 19440
rect 10226 19388 10232 19440
rect 10284 19428 10290 19440
rect 10594 19428 10600 19440
rect 10284 19400 10600 19428
rect 10284 19388 10290 19400
rect 10594 19388 10600 19400
rect 10652 19428 10658 19440
rect 11606 19428 11612 19440
rect 10652 19400 11612 19428
rect 10652 19388 10658 19400
rect 11606 19388 11612 19400
rect 11664 19388 11670 19440
rect 12176 19437 12204 19468
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 13504 19468 13768 19496
rect 13504 19456 13510 19468
rect 12161 19431 12219 19437
rect 12161 19397 12173 19431
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 12250 19388 12256 19440
rect 12308 19428 12314 19440
rect 12308 19400 12353 19428
rect 12308 19388 12314 19400
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 13538 19428 13544 19440
rect 12492 19400 13544 19428
rect 12492 19388 12498 19400
rect 13538 19388 13544 19400
rect 13596 19388 13602 19440
rect 13740 19437 13768 19468
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 14976 19468 15424 19496
rect 14976 19456 14982 19468
rect 13725 19431 13783 19437
rect 13725 19397 13737 19431
rect 13771 19397 13783 19431
rect 13725 19391 13783 19397
rect 13814 19388 13820 19440
rect 13872 19428 13878 19440
rect 13872 19400 13917 19428
rect 13872 19388 13878 19400
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 14737 19431 14795 19437
rect 14737 19428 14749 19431
rect 14608 19400 14749 19428
rect 14608 19388 14614 19400
rect 14737 19397 14749 19400
rect 14783 19397 14795 19431
rect 14737 19391 14795 19397
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 15396 19437 15424 19468
rect 16022 19456 16028 19508
rect 16080 19496 16086 19508
rect 16482 19496 16488 19508
rect 16080 19468 16488 19496
rect 16080 19456 16086 19468
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 18506 19496 18512 19508
rect 17052 19468 18512 19496
rect 15289 19431 15347 19437
rect 15289 19428 15301 19431
rect 14884 19400 15301 19428
rect 14884 19388 14890 19400
rect 15289 19397 15301 19400
rect 15335 19397 15347 19431
rect 15289 19391 15347 19397
rect 15381 19431 15439 19437
rect 15381 19397 15393 19431
rect 15427 19397 15439 19431
rect 15381 19391 15439 19397
rect 15562 19388 15568 19440
rect 15620 19428 15626 19440
rect 16301 19431 16359 19437
rect 16301 19428 16313 19431
rect 15620 19400 16313 19428
rect 15620 19388 15626 19400
rect 16301 19397 16313 19400
rect 16347 19397 16359 19431
rect 16942 19428 16948 19440
rect 16903 19400 16948 19428
rect 16301 19391 16359 19397
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 17052 19437 17080 19468
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 18966 19496 18972 19508
rect 18616 19468 18972 19496
rect 17037 19431 17095 19437
rect 17037 19397 17049 19431
rect 17083 19397 17095 19431
rect 17037 19391 17095 19397
rect 17218 19388 17224 19440
rect 17276 19428 17282 19440
rect 18616 19428 18644 19468
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 19978 19496 19984 19508
rect 19537 19468 19984 19496
rect 17276 19400 18644 19428
rect 18693 19431 18751 19437
rect 17276 19388 17282 19400
rect 18693 19397 18705 19431
rect 18739 19428 18751 19431
rect 18782 19428 18788 19440
rect 18739 19400 18788 19428
rect 18739 19397 18751 19400
rect 18693 19391 18751 19397
rect 18782 19388 18788 19400
rect 18840 19388 18846 19440
rect 19537 19428 19565 19468
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20162 19496 20168 19508
rect 20123 19468 20168 19496
rect 20162 19456 20168 19468
rect 20220 19456 20226 19508
rect 20438 19456 20444 19508
rect 20496 19496 20502 19508
rect 20496 19468 20576 19496
rect 20496 19456 20502 19468
rect 19444 19400 19565 19428
rect 6825 19363 6883 19369
rect 6825 19329 6837 19363
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 6972 19332 7481 19360
rect 6972 19320 6978 19332
rect 7469 19329 7481 19332
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 3970 19292 3976 19304
rect 2087 19264 3832 19292
rect 3931 19264 3976 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 3804 19156 3832 19264
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19292 4307 19295
rect 5994 19292 6000 19304
rect 4295 19264 6000 19292
rect 4295 19261 4307 19264
rect 4249 19255 4307 19261
rect 5994 19252 6000 19264
rect 6052 19252 6058 19304
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 7800 19264 7845 19292
rect 7800 19252 7806 19264
rect 5810 19184 5816 19236
rect 5868 19224 5874 19236
rect 6270 19224 6276 19236
rect 5868 19196 6276 19224
rect 5868 19184 5874 19196
rect 6270 19184 6276 19196
rect 6328 19184 6334 19236
rect 8864 19224 8892 19346
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 11296 19332 12020 19360
rect 11296 19320 11302 19332
rect 9030 19252 9036 19304
rect 9088 19292 9094 19304
rect 9674 19292 9680 19304
rect 9088 19264 9680 19292
rect 9088 19252 9094 19264
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 9916 19264 10057 19292
rect 9916 19252 9922 19264
rect 10045 19261 10057 19264
rect 10091 19292 10103 19295
rect 10410 19292 10416 19304
rect 10091 19264 10416 19292
rect 10091 19261 10103 19264
rect 10045 19255 10103 19261
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 10873 19295 10931 19301
rect 10873 19261 10885 19295
rect 10919 19261 10931 19295
rect 11992 19292 12020 19332
rect 13078 19320 13084 19372
rect 13136 19320 13142 19372
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 18196 19332 18460 19360
rect 18196 19320 18202 19332
rect 12434 19292 12440 19304
rect 11992 19264 12440 19292
rect 10873 19255 10931 19261
rect 9950 19224 9956 19236
rect 8864 19196 9956 19224
rect 9950 19184 9956 19196
rect 10008 19184 10014 19236
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 10888 19224 10916 19255
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 13096 19292 13124 19320
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 13096 19264 13185 19292
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13173 19255 13231 19261
rect 13446 19252 13452 19304
rect 13504 19292 13510 19304
rect 17126 19292 17132 19304
rect 13504 19264 17132 19292
rect 13504 19252 13510 19264
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17586 19292 17592 19304
rect 17547 19264 17592 19292
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18432 19292 18460 19332
rect 18601 19295 18659 19301
rect 18601 19292 18613 19295
rect 17920 19264 18276 19292
rect 18432 19264 18613 19292
rect 17920 19252 17926 19264
rect 12526 19224 12532 19236
rect 10836 19196 10916 19224
rect 11164 19196 12532 19224
rect 10836 19184 10842 19196
rect 5902 19156 5908 19168
rect 3804 19128 5908 19156
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 6917 19159 6975 19165
rect 6917 19125 6929 19159
rect 6963 19156 6975 19159
rect 8294 19156 8300 19168
rect 6963 19128 8300 19156
rect 6963 19125 6975 19128
rect 6917 19119 6975 19125
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8478 19116 8484 19168
rect 8536 19156 8542 19168
rect 11164 19156 11192 19196
rect 12526 19184 12532 19196
rect 12584 19184 12590 19236
rect 18138 19224 18144 19236
rect 12636 19196 18144 19224
rect 8536 19128 11192 19156
rect 8536 19116 8542 19128
rect 11238 19116 11244 19168
rect 11296 19156 11302 19168
rect 12636 19156 12664 19196
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18248 19224 18276 19264
rect 18601 19261 18613 19264
rect 18647 19261 18659 19295
rect 18874 19292 18880 19304
rect 18835 19264 18880 19292
rect 18601 19255 18659 19261
rect 18874 19252 18880 19264
rect 18932 19252 18938 19304
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19444 19292 19472 19400
rect 19610 19388 19616 19440
rect 19668 19428 19674 19440
rect 20548 19428 20576 19468
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 20680 19468 20944 19496
rect 20680 19456 20686 19468
rect 20916 19437 20944 19468
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22244 19468 22600 19496
rect 22244 19456 22250 19468
rect 20809 19431 20867 19437
rect 20809 19428 20821 19431
rect 19668 19400 20392 19428
rect 20548 19400 20821 19428
rect 19668 19388 19674 19400
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19360 20131 19363
rect 20254 19360 20260 19372
rect 20119 19332 20260 19360
rect 20119 19329 20131 19332
rect 20073 19323 20131 19329
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20364 19360 20392 19400
rect 20809 19397 20821 19400
rect 20855 19397 20867 19431
rect 20809 19391 20867 19397
rect 20901 19431 20959 19437
rect 20901 19397 20913 19431
rect 20947 19397 20959 19431
rect 22462 19428 22468 19440
rect 22423 19400 22468 19428
rect 20901 19391 20959 19397
rect 22462 19388 22468 19400
rect 22520 19388 22526 19440
rect 22572 19437 22600 19468
rect 23934 19456 23940 19508
rect 23992 19496 23998 19508
rect 23992 19468 28948 19496
rect 23992 19456 23998 19468
rect 22557 19431 22615 19437
rect 22557 19397 22569 19431
rect 22603 19397 22615 19431
rect 24026 19428 24032 19440
rect 22557 19391 22615 19397
rect 23308 19400 24032 19428
rect 20622 19360 20628 19372
rect 20364 19332 20628 19360
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 19024 19264 19472 19292
rect 19024 19252 19030 19264
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 20438 19292 20444 19304
rect 19668 19264 20444 19292
rect 19668 19252 19674 19264
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 20530 19252 20536 19304
rect 20588 19292 20594 19304
rect 21085 19295 21143 19301
rect 21085 19292 21097 19295
rect 20588 19264 21097 19292
rect 20588 19252 20594 19264
rect 21085 19261 21097 19264
rect 21131 19261 21143 19295
rect 21085 19255 21143 19261
rect 21266 19252 21272 19304
rect 21324 19292 21330 19304
rect 23308 19292 23336 19400
rect 24026 19388 24032 19400
rect 24084 19388 24090 19440
rect 24121 19431 24179 19437
rect 24121 19397 24133 19431
rect 24167 19428 24179 19431
rect 25590 19428 25596 19440
rect 24167 19400 25452 19428
rect 25551 19400 25596 19428
rect 24167 19397 24179 19400
rect 24121 19391 24179 19397
rect 21324 19264 23336 19292
rect 23385 19295 23443 19301
rect 21324 19252 21330 19264
rect 23385 19261 23397 19295
rect 23431 19292 23443 19295
rect 24670 19292 24676 19304
rect 23431 19264 24676 19292
rect 23431 19261 23443 19264
rect 23385 19255 23443 19261
rect 19628 19224 19656 19252
rect 18248 19196 19656 19224
rect 19702 19184 19708 19236
rect 19760 19224 19766 19236
rect 21634 19224 21640 19236
rect 19760 19196 21640 19224
rect 19760 19184 19766 19196
rect 21634 19184 21640 19196
rect 21692 19184 21698 19236
rect 11296 19128 12664 19156
rect 11296 19116 11302 19128
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 20438 19156 20444 19168
rect 12952 19128 20444 19156
rect 12952 19116 12958 19128
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 20714 19116 20720 19168
rect 20772 19156 20778 19168
rect 23400 19156 23428 19255
rect 24670 19252 24676 19264
rect 24728 19252 24734 19304
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 25314 19292 25320 19304
rect 25188 19264 25320 19292
rect 25188 19252 25194 19264
rect 25314 19252 25320 19264
rect 25372 19252 25378 19304
rect 24486 19184 24492 19236
rect 24544 19224 24550 19236
rect 24581 19227 24639 19233
rect 24581 19224 24593 19227
rect 24544 19196 24593 19224
rect 24544 19184 24550 19196
rect 24581 19193 24593 19196
rect 24627 19193 24639 19227
rect 25424 19224 25452 19400
rect 25590 19388 25596 19400
rect 25648 19388 25654 19440
rect 25685 19431 25743 19437
rect 25685 19397 25697 19431
rect 25731 19428 25743 19431
rect 26418 19428 26424 19440
rect 25731 19400 26424 19428
rect 25731 19397 25743 19400
rect 25685 19391 25743 19397
rect 26418 19388 26424 19400
rect 26476 19388 26482 19440
rect 26605 19431 26663 19437
rect 26605 19397 26617 19431
rect 26651 19428 26663 19431
rect 26970 19428 26976 19440
rect 26651 19400 26976 19428
rect 26651 19397 26663 19400
rect 26605 19391 26663 19397
rect 26970 19388 26976 19400
rect 27028 19388 27034 19440
rect 27338 19428 27344 19440
rect 27299 19400 27344 19428
rect 27338 19388 27344 19400
rect 27396 19388 27402 19440
rect 27614 19388 27620 19440
rect 27672 19428 27678 19440
rect 28261 19431 28319 19437
rect 28261 19428 28273 19431
rect 27672 19400 28273 19428
rect 27672 19388 27678 19400
rect 28261 19397 28273 19400
rect 28307 19397 28319 19431
rect 28810 19428 28816 19440
rect 28771 19400 28816 19428
rect 28261 19391 28319 19397
rect 28810 19388 28816 19400
rect 28868 19388 28874 19440
rect 28920 19437 28948 19468
rect 29914 19456 29920 19508
rect 29972 19496 29978 19508
rect 31573 19499 31631 19505
rect 31573 19496 31585 19499
rect 29972 19468 31585 19496
rect 29972 19456 29978 19468
rect 31573 19465 31585 19468
rect 31619 19465 31631 19499
rect 31573 19459 31631 19465
rect 37645 19499 37703 19505
rect 37645 19465 37657 19499
rect 37691 19496 37703 19499
rect 37918 19496 37924 19508
rect 37691 19468 37924 19496
rect 37691 19465 37703 19468
rect 37645 19459 37703 19465
rect 37918 19456 37924 19468
rect 37976 19456 37982 19508
rect 28905 19431 28963 19437
rect 28905 19397 28917 19431
rect 28951 19397 28963 19431
rect 29822 19428 29828 19440
rect 29783 19400 29828 19428
rect 28905 19391 28963 19397
rect 29822 19388 29828 19400
rect 29880 19428 29886 19440
rect 30190 19428 30196 19440
rect 29880 19400 30196 19428
rect 29880 19388 29886 19400
rect 30190 19388 30196 19400
rect 30248 19388 30254 19440
rect 30374 19428 30380 19440
rect 30335 19400 30380 19428
rect 30374 19388 30380 19400
rect 30432 19388 30438 19440
rect 30469 19431 30527 19437
rect 30469 19397 30481 19431
rect 30515 19428 30527 19431
rect 30558 19428 30564 19440
rect 30515 19400 30564 19428
rect 30515 19397 30527 19400
rect 30469 19391 30527 19397
rect 30558 19388 30564 19400
rect 30616 19388 30622 19440
rect 31478 19360 31484 19372
rect 31439 19332 31484 19360
rect 31478 19320 31484 19332
rect 31536 19320 31542 19372
rect 37826 19360 37832 19372
rect 37787 19332 37832 19360
rect 37826 19320 37832 19332
rect 37884 19320 37890 19372
rect 25590 19252 25596 19304
rect 25648 19292 25654 19304
rect 27249 19295 27307 19301
rect 27249 19292 27261 19295
rect 25648 19264 27261 19292
rect 25648 19252 25654 19264
rect 27249 19261 27261 19264
rect 27295 19261 27307 19295
rect 27249 19255 27307 19261
rect 29454 19252 29460 19304
rect 29512 19292 29518 19304
rect 30098 19292 30104 19304
rect 29512 19264 30104 19292
rect 29512 19252 29518 19264
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 30650 19292 30656 19304
rect 30611 19264 30656 19292
rect 30650 19252 30656 19264
rect 30708 19252 30714 19304
rect 26878 19224 26884 19236
rect 25424 19196 26884 19224
rect 24581 19187 24639 19193
rect 26878 19184 26884 19196
rect 26936 19184 26942 19236
rect 27062 19184 27068 19236
rect 27120 19224 27126 19236
rect 28074 19224 28080 19236
rect 27120 19196 28080 19224
rect 27120 19184 27126 19196
rect 28074 19184 28080 19196
rect 28132 19184 28138 19236
rect 20772 19128 23428 19156
rect 20772 19116 20778 19128
rect 26786 19116 26792 19168
rect 26844 19156 26850 19168
rect 28258 19156 28264 19168
rect 26844 19128 28264 19156
rect 26844 19116 26850 19128
rect 28258 19116 28264 19128
rect 28316 19116 28322 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 2096 18924 3341 18952
rect 2096 18912 2102 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 3329 18915 3387 18921
rect 9309 18955 9367 18961
rect 9309 18921 9321 18955
rect 9355 18952 9367 18955
rect 14918 18952 14924 18964
rect 9355 18924 14924 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 14918 18912 14924 18924
rect 14976 18912 14982 18964
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 15838 18952 15844 18964
rect 15528 18924 15844 18952
rect 15528 18912 15534 18924
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 17862 18952 17868 18964
rect 16908 18924 17868 18952
rect 16908 18912 16914 18924
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18966 18952 18972 18964
rect 18064 18924 18972 18952
rect 8110 18844 8116 18896
rect 8168 18884 8174 18896
rect 9858 18884 9864 18896
rect 8168 18856 9864 18884
rect 8168 18844 8174 18856
rect 9858 18844 9864 18856
rect 9916 18844 9922 18896
rect 11609 18887 11667 18893
rect 11609 18853 11621 18887
rect 11655 18884 11667 18887
rect 11974 18884 11980 18896
rect 11655 18856 11980 18884
rect 11655 18853 11667 18856
rect 11609 18847 11667 18853
rect 11974 18844 11980 18856
rect 12032 18884 12038 18896
rect 12250 18884 12256 18896
rect 12032 18856 12256 18884
rect 12032 18844 12038 18856
rect 12250 18844 12256 18856
rect 12308 18844 12314 18896
rect 14090 18884 14096 18896
rect 12360 18856 14096 18884
rect 1581 18819 1639 18825
rect 1581 18785 1593 18819
rect 1627 18816 1639 18819
rect 1854 18816 1860 18828
rect 1627 18788 1860 18816
rect 1627 18785 1639 18788
rect 1581 18779 1639 18785
rect 1854 18776 1860 18788
rect 1912 18816 1918 18828
rect 3970 18816 3976 18828
rect 1912 18788 3976 18816
rect 1912 18776 1918 18788
rect 3970 18776 3976 18788
rect 4028 18776 4034 18828
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18816 4307 18819
rect 4798 18816 4804 18828
rect 4295 18788 4804 18816
rect 4295 18785 4307 18788
rect 4249 18779 4307 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 5994 18816 6000 18828
rect 5907 18788 6000 18816
rect 5994 18776 6000 18788
rect 6052 18816 6058 18828
rect 11146 18816 11152 18828
rect 6052 18788 11152 18816
rect 6052 18776 6058 18788
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 12360 18825 12388 18856
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 17218 18884 17224 18896
rect 14200 18856 17224 18884
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 13446 18816 13452 18828
rect 12584 18788 13452 18816
rect 12584 18776 12590 18788
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14200 18816 14228 18856
rect 17218 18844 17224 18856
rect 17276 18844 17282 18896
rect 17402 18844 17408 18896
rect 17460 18884 17466 18896
rect 18064 18884 18092 18924
rect 18966 18912 18972 18924
rect 19024 18912 19030 18964
rect 19537 18924 19741 18952
rect 17460 18856 18092 18884
rect 17460 18844 17466 18856
rect 18138 18844 18144 18896
rect 18196 18884 18202 18896
rect 19537 18884 19565 18924
rect 18196 18856 19565 18884
rect 19713 18884 19741 18924
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 26418 18952 26424 18964
rect 20036 18924 26424 18952
rect 20036 18912 20042 18924
rect 26418 18912 26424 18924
rect 26476 18912 26482 18964
rect 26878 18952 26884 18964
rect 26839 18924 26884 18952
rect 26878 18912 26884 18924
rect 26936 18912 26942 18964
rect 27062 18912 27068 18964
rect 27120 18952 27126 18964
rect 27120 18924 30144 18952
rect 27120 18912 27126 18924
rect 22002 18884 22008 18896
rect 19713 18856 22008 18884
rect 18196 18844 18202 18856
rect 22002 18844 22008 18856
rect 22060 18844 22066 18896
rect 24946 18844 24952 18896
rect 25004 18884 25010 18896
rect 30006 18884 30012 18896
rect 25004 18856 30012 18884
rect 25004 18844 25010 18856
rect 30006 18844 30012 18856
rect 30064 18844 30070 18896
rect 17954 18816 17960 18828
rect 13872 18788 14228 18816
rect 15304 18788 17960 18816
rect 13872 18776 13878 18788
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 6546 18748 6552 18760
rect 6507 18720 6552 18748
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 7958 18720 9168 18748
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 2866 18640 2872 18692
rect 2924 18640 2930 18692
rect 6825 18683 6883 18689
rect 6825 18649 6837 18683
rect 6871 18649 6883 18683
rect 6825 18643 6883 18649
rect 8573 18683 8631 18689
rect 8573 18649 8585 18683
rect 8619 18680 8631 18683
rect 8754 18680 8760 18692
rect 8619 18652 8760 18680
rect 8619 18649 8631 18652
rect 8573 18643 8631 18649
rect 6840 18612 6868 18643
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 9140 18680 9168 18720
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9272 18720 9317 18748
rect 9272 18708 9278 18720
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9732 18720 9873 18748
rect 9732 18708 9738 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 10042 18680 10048 18692
rect 9140 18652 10048 18680
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10137 18683 10195 18689
rect 10137 18649 10149 18683
rect 10183 18649 10195 18683
rect 11362 18652 11836 18680
rect 10137 18643 10195 18649
rect 8478 18612 8484 18624
rect 6840 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 10152 18612 10180 18643
rect 11422 18612 11428 18624
rect 10152 18584 11428 18612
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 11808 18612 11836 18652
rect 11882 18640 11888 18692
rect 11940 18680 11946 18692
rect 12437 18683 12495 18689
rect 12437 18680 12449 18683
rect 11940 18652 12449 18680
rect 11940 18640 11946 18652
rect 12437 18649 12449 18652
rect 12483 18649 12495 18683
rect 12437 18643 12495 18649
rect 13170 18640 13176 18692
rect 13228 18680 13234 18692
rect 13357 18683 13415 18689
rect 13357 18680 13369 18683
rect 13228 18652 13369 18680
rect 13228 18640 13234 18652
rect 13357 18649 13369 18652
rect 13403 18680 13415 18683
rect 13403 18652 14136 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13814 18612 13820 18624
rect 11808 18584 13820 18612
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 14108 18612 14136 18652
rect 14182 18640 14188 18692
rect 14240 18680 14246 18692
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 14240 18652 14381 18680
rect 14240 18640 14246 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14461 18683 14519 18689
rect 14461 18649 14473 18683
rect 14507 18680 14519 18683
rect 15304 18680 15332 18788
rect 17954 18776 17960 18788
rect 18012 18776 18018 18828
rect 18230 18816 18236 18828
rect 18064 18788 18236 18816
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15528 18720 15853 18748
rect 15528 18708 15534 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18748 17739 18751
rect 18064 18748 18092 18788
rect 18230 18776 18236 18788
rect 18288 18776 18294 18828
rect 18877 18819 18935 18825
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 19334 18816 19340 18828
rect 18923 18788 19340 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 19610 18776 19616 18828
rect 19668 18816 19674 18828
rect 19889 18819 19947 18825
rect 19889 18816 19901 18819
rect 19668 18788 19901 18816
rect 19668 18776 19674 18788
rect 19889 18785 19901 18788
rect 19935 18785 19947 18819
rect 20530 18816 20536 18828
rect 20491 18788 20536 18816
rect 19889 18779 19947 18785
rect 20530 18776 20536 18788
rect 20588 18776 20594 18828
rect 21085 18819 21143 18825
rect 21085 18785 21097 18819
rect 21131 18816 21143 18819
rect 21266 18816 21272 18828
rect 21131 18788 21272 18816
rect 21131 18785 21143 18788
rect 21085 18779 21143 18785
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 22281 18819 22339 18825
rect 22281 18785 22293 18819
rect 22327 18816 22339 18819
rect 22462 18816 22468 18828
rect 22327 18788 22468 18816
rect 22327 18785 22339 18788
rect 22281 18779 22339 18785
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 22922 18816 22928 18828
rect 22883 18788 22928 18816
rect 22922 18776 22928 18788
rect 22980 18776 22986 18828
rect 25498 18816 25504 18828
rect 23768 18788 25504 18816
rect 17727 18720 18092 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 14507 18652 15332 18680
rect 14507 18649 14519 18652
rect 14461 18643 14519 18649
rect 15378 18640 15384 18692
rect 15436 18680 15442 18692
rect 15436 18652 15481 18680
rect 15436 18640 15442 18652
rect 15562 18640 15568 18692
rect 15620 18680 15626 18692
rect 16117 18683 16175 18689
rect 16117 18680 16129 18683
rect 15620 18652 16129 18680
rect 15620 18640 15626 18652
rect 16117 18649 16129 18652
rect 16163 18649 16175 18683
rect 16117 18643 16175 18649
rect 15654 18612 15660 18624
rect 14108 18584 15660 18612
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 16132 18612 16160 18643
rect 16850 18640 16856 18692
rect 16908 18680 16914 18692
rect 17026 18683 17084 18689
rect 17026 18680 17038 18683
rect 16908 18652 17038 18680
rect 16908 18640 16914 18652
rect 17026 18649 17038 18652
rect 17072 18649 17084 18683
rect 17026 18643 17084 18649
rect 17122 18683 17180 18689
rect 17122 18649 17134 18683
rect 17168 18680 17180 18683
rect 17402 18680 17408 18692
rect 17168 18652 17408 18680
rect 17168 18649 17180 18652
rect 17122 18643 17180 18649
rect 17402 18640 17408 18652
rect 17460 18640 17466 18692
rect 18064 18624 18092 18720
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19024 18720 19380 18748
rect 19024 18708 19030 18720
rect 18233 18683 18291 18689
rect 18233 18649 18245 18683
rect 18279 18649 18291 18683
rect 18233 18643 18291 18649
rect 18325 18683 18383 18689
rect 18325 18649 18337 18683
rect 18371 18680 18383 18683
rect 19242 18680 19248 18692
rect 18371 18652 19248 18680
rect 18371 18649 18383 18652
rect 18325 18643 18383 18649
rect 17954 18612 17960 18624
rect 16132 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18046 18572 18052 18624
rect 18104 18572 18110 18624
rect 18248 18612 18276 18643
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 19352 18680 19380 18720
rect 19702 18680 19708 18692
rect 19352 18652 19708 18680
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 19971 18680 19977 18692
rect 19932 18652 19977 18680
rect 19971 18640 19977 18652
rect 20029 18640 20035 18692
rect 20548 18680 20576 18776
rect 23474 18748 23480 18760
rect 23124 18720 23480 18748
rect 21177 18683 21235 18689
rect 20548 18652 21036 18680
rect 21008 18624 21036 18652
rect 21177 18649 21189 18683
rect 21223 18649 21235 18683
rect 21177 18643 21235 18649
rect 18966 18612 18972 18624
rect 18248 18584 18972 18612
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 20714 18612 20720 18624
rect 19392 18584 20720 18612
rect 19392 18572 19398 18584
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 20990 18572 20996 18624
rect 21048 18572 21054 18624
rect 21192 18612 21220 18643
rect 21266 18640 21272 18692
rect 21324 18680 21330 18692
rect 21729 18683 21787 18689
rect 21729 18680 21741 18683
rect 21324 18652 21741 18680
rect 21324 18640 21330 18652
rect 21729 18649 21741 18652
rect 21775 18649 21787 18683
rect 21729 18643 21787 18649
rect 22373 18683 22431 18689
rect 22373 18649 22385 18683
rect 22419 18680 22431 18683
rect 23124 18680 23152 18720
rect 23474 18708 23480 18720
rect 23532 18708 23538 18760
rect 23768 18757 23796 18788
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25958 18816 25964 18828
rect 25740 18788 25964 18816
rect 25740 18776 25746 18788
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 29086 18816 29092 18828
rect 27356 18788 29092 18816
rect 23753 18751 23811 18757
rect 23753 18717 23765 18751
rect 23799 18717 23811 18751
rect 26142 18748 26148 18760
rect 26103 18720 26148 18748
rect 23753 18711 23811 18717
rect 26142 18708 26148 18720
rect 26200 18708 26206 18760
rect 26786 18748 26792 18760
rect 26747 18720 26792 18748
rect 26786 18708 26792 18720
rect 26844 18708 26850 18760
rect 22419 18652 23152 18680
rect 22419 18649 22431 18652
rect 22373 18643 22431 18649
rect 24670 18640 24676 18692
rect 24728 18680 24734 18692
rect 25041 18683 25099 18689
rect 25041 18680 25053 18683
rect 24728 18652 25053 18680
rect 24728 18640 24734 18652
rect 25041 18649 25053 18652
rect 25087 18649 25099 18683
rect 25041 18643 25099 18649
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25188 18652 25233 18680
rect 25188 18640 25194 18652
rect 25958 18640 25964 18692
rect 26016 18680 26022 18692
rect 27356 18680 27384 18788
rect 29086 18776 29092 18788
rect 29144 18776 29150 18828
rect 29825 18819 29883 18825
rect 29825 18785 29837 18819
rect 29871 18816 29883 18819
rect 29914 18816 29920 18828
rect 29871 18788 29920 18816
rect 29871 18785 29883 18788
rect 29825 18779 29883 18785
rect 29914 18776 29920 18788
rect 29972 18776 29978 18828
rect 30116 18825 30144 18924
rect 30190 18844 30196 18896
rect 30248 18884 30254 18896
rect 30248 18856 31524 18884
rect 30248 18844 30254 18856
rect 30101 18819 30159 18825
rect 30101 18785 30113 18819
rect 30147 18785 30159 18819
rect 30101 18779 30159 18785
rect 31205 18819 31263 18825
rect 31205 18785 31217 18819
rect 31251 18816 31263 18819
rect 31386 18816 31392 18828
rect 31251 18788 31392 18816
rect 31251 18785 31263 18788
rect 31205 18779 31263 18785
rect 31386 18776 31392 18788
rect 31444 18776 31450 18828
rect 31496 18825 31524 18856
rect 31481 18819 31539 18825
rect 31481 18785 31493 18819
rect 31527 18785 31539 18819
rect 31481 18779 31539 18785
rect 28626 18748 28632 18760
rect 28587 18720 28632 18748
rect 28626 18708 28632 18720
rect 28684 18708 28690 18760
rect 32674 18748 32680 18760
rect 32635 18720 32680 18748
rect 32674 18708 32680 18720
rect 32732 18708 32738 18760
rect 38286 18748 38292 18760
rect 38247 18720 38292 18748
rect 38286 18708 38292 18720
rect 38344 18708 38350 18760
rect 27525 18683 27583 18689
rect 27525 18680 27537 18683
rect 26016 18652 27537 18680
rect 26016 18640 26022 18652
rect 27525 18649 27537 18652
rect 27571 18649 27583 18683
rect 27525 18643 27583 18649
rect 27617 18683 27675 18689
rect 27617 18649 27629 18683
rect 27663 18680 27675 18683
rect 27798 18680 27804 18692
rect 27663 18652 27804 18680
rect 27663 18649 27675 18652
rect 27617 18643 27675 18649
rect 27798 18640 27804 18652
rect 27856 18640 27862 18692
rect 28169 18683 28227 18689
rect 28169 18649 28181 18683
rect 28215 18680 28227 18683
rect 29362 18680 29368 18692
rect 28215 18652 29368 18680
rect 28215 18649 28227 18652
rect 28169 18643 28227 18649
rect 23845 18615 23903 18621
rect 23845 18612 23857 18615
rect 21192 18584 23857 18612
rect 23845 18581 23857 18584
rect 23891 18581 23903 18615
rect 23845 18575 23903 18581
rect 24026 18572 24032 18624
rect 24084 18612 24090 18624
rect 26237 18615 26295 18621
rect 26237 18612 26249 18615
rect 24084 18584 26249 18612
rect 24084 18572 24090 18584
rect 26237 18581 26249 18584
rect 26283 18581 26295 18615
rect 26237 18575 26295 18581
rect 26326 18572 26332 18624
rect 26384 18612 26390 18624
rect 28184 18612 28212 18643
rect 29362 18640 29368 18652
rect 29420 18640 29426 18692
rect 29914 18640 29920 18692
rect 29972 18680 29978 18692
rect 31294 18680 31300 18692
rect 29972 18652 30017 18680
rect 31255 18652 31300 18680
rect 29972 18640 29978 18652
rect 31294 18640 31300 18652
rect 31352 18640 31358 18692
rect 28718 18612 28724 18624
rect 26384 18584 28212 18612
rect 28679 18584 28724 18612
rect 26384 18572 26390 18584
rect 28718 18572 28724 18584
rect 28776 18572 28782 18624
rect 28810 18572 28816 18624
rect 28868 18612 28874 18624
rect 32769 18615 32827 18621
rect 32769 18612 32781 18615
rect 28868 18584 32781 18612
rect 28868 18572 28874 18584
rect 32769 18581 32781 18584
rect 32815 18581 32827 18615
rect 32769 18575 32827 18581
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 34572 18584 38117 18612
rect 34572 18572 34578 18584
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 12342 18408 12348 18420
rect 1912 18380 8708 18408
rect 1912 18368 1918 18380
rect 2222 18340 2228 18352
rect 2183 18312 2228 18340
rect 2222 18300 2228 18312
rect 2280 18300 2286 18352
rect 3145 18343 3203 18349
rect 3145 18309 3157 18343
rect 3191 18340 3203 18343
rect 4154 18340 4160 18352
rect 3191 18312 4160 18340
rect 3191 18309 3203 18312
rect 3145 18303 3203 18309
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 5644 18349 5672 18380
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18309 5687 18343
rect 8680 18340 8708 18380
rect 9416 18380 12348 18408
rect 9416 18340 9444 18380
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 18874 18408 18880 18420
rect 13372 18380 18880 18408
rect 8680 18312 9444 18340
rect 5629 18303 5687 18309
rect 10134 18300 10140 18352
rect 10192 18300 10198 18352
rect 12437 18343 12495 18349
rect 12437 18340 12449 18343
rect 10888 18312 12449 18340
rect 6454 18272 6460 18284
rect 5014 18244 6460 18272
rect 6454 18232 6460 18244
rect 6512 18232 6518 18284
rect 8202 18232 8208 18284
rect 8260 18232 8266 18284
rect 9316 18275 9374 18281
rect 9316 18272 9328 18275
rect 9232 18244 9328 18272
rect 9232 18216 9260 18244
rect 9316 18241 9328 18244
rect 9362 18241 9374 18275
rect 10888 18272 10916 18312
rect 12437 18309 12449 18312
rect 12483 18309 12495 18343
rect 12437 18303 12495 18309
rect 12526 18300 12532 18352
rect 12584 18340 12590 18352
rect 13262 18340 13268 18352
rect 12584 18312 13268 18340
rect 12584 18300 12590 18312
rect 13262 18300 13268 18312
rect 13320 18300 13326 18352
rect 13372 18349 13400 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 18969 18411 19027 18417
rect 18969 18377 18981 18411
rect 19015 18408 19027 18411
rect 19426 18408 19432 18420
rect 19015 18380 19432 18408
rect 19015 18377 19027 18380
rect 18969 18371 19027 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 20806 18408 20812 18420
rect 19628 18380 20812 18408
rect 19628 18352 19656 18380
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 20925 18380 21404 18408
rect 13357 18343 13415 18349
rect 13357 18309 13369 18343
rect 13403 18309 13415 18343
rect 13357 18303 13415 18309
rect 9316 18235 9374 18241
rect 10796 18244 10916 18272
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 2314 18204 2320 18216
rect 2179 18176 2320 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 3605 18207 3663 18213
rect 3605 18173 3617 18207
rect 3651 18204 3663 18207
rect 3878 18204 3884 18216
rect 3651 18176 3740 18204
rect 3839 18176 3884 18204
rect 3651 18173 3663 18176
rect 3605 18167 3663 18173
rect 3712 18068 3740 18176
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4246 18164 4252 18216
rect 4304 18204 4310 18216
rect 6822 18204 6828 18216
rect 4304 18176 5488 18204
rect 6783 18176 6828 18204
rect 4304 18164 4310 18176
rect 5460 18148 5488 18176
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 7101 18207 7159 18213
rect 7101 18173 7113 18207
rect 7147 18204 7159 18207
rect 7834 18204 7840 18216
rect 7147 18176 7840 18204
rect 7147 18173 7159 18176
rect 7101 18167 7159 18173
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8628 18176 8861 18204
rect 8628 18164 8634 18176
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 8849 18167 8907 18173
rect 9214 18164 9220 18216
rect 9272 18164 9278 18216
rect 10796 18204 10824 18244
rect 11606 18232 11612 18284
rect 11664 18272 11670 18284
rect 11664 18244 12020 18272
rect 11664 18232 11670 18244
rect 9416 18176 10824 18204
rect 5442 18096 5448 18148
rect 5500 18136 5506 18148
rect 9416 18136 9444 18176
rect 10870 18164 10876 18216
rect 10928 18204 10934 18216
rect 11882 18204 11888 18216
rect 10928 18176 11888 18204
rect 10928 18164 10934 18176
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 11992 18204 12020 18244
rect 12345 18207 12403 18213
rect 12345 18204 12357 18207
rect 11992 18176 12357 18204
rect 12345 18173 12357 18176
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 12986 18204 12992 18216
rect 12768 18176 12992 18204
rect 12768 18164 12774 18176
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 5500 18108 6960 18136
rect 5500 18096 5506 18108
rect 6932 18080 6960 18108
rect 8496 18108 9444 18136
rect 4614 18068 4620 18080
rect 3712 18040 4620 18068
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 6086 18068 6092 18080
rect 5408 18040 6092 18068
rect 5408 18028 5414 18040
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6914 18028 6920 18080
rect 6972 18028 6978 18080
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 8496 18068 8524 18108
rect 12066 18096 12072 18148
rect 12124 18136 12130 18148
rect 13372 18136 13400 18303
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 14185 18343 14243 18349
rect 14185 18340 14197 18343
rect 13504 18312 14197 18340
rect 13504 18300 13510 18312
rect 14185 18309 14197 18312
rect 14231 18309 14243 18343
rect 14185 18303 14243 18309
rect 15381 18343 15439 18349
rect 15381 18309 15393 18343
rect 15427 18340 15439 18343
rect 16942 18340 16948 18352
rect 15427 18312 16804 18340
rect 16903 18312 16948 18340
rect 15427 18309 15439 18312
rect 15381 18303 15439 18309
rect 16666 18272 16672 18284
rect 16132 18244 16672 18272
rect 14093 18207 14151 18213
rect 14093 18173 14105 18207
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 12124 18108 13400 18136
rect 14108 18136 14136 18167
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14240 18176 14381 18204
rect 14240 18164 14246 18176
rect 14369 18173 14381 18176
rect 14415 18204 14427 18207
rect 14918 18204 14924 18216
rect 14415 18176 14924 18204
rect 14415 18173 14427 18176
rect 14369 18167 14427 18173
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18204 15347 18207
rect 15470 18204 15476 18216
rect 15335 18176 15476 18204
rect 15335 18173 15347 18176
rect 15289 18167 15347 18173
rect 15304 18136 15332 18167
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 14108 18108 15332 18136
rect 12124 18096 12130 18108
rect 9582 18077 9588 18080
rect 7156 18040 8524 18068
rect 9566 18071 9588 18077
rect 7156 18028 7162 18040
rect 9566 18037 9578 18071
rect 9566 18031 9588 18037
rect 9582 18028 9588 18031
rect 9640 18028 9646 18080
rect 11057 18071 11115 18077
rect 11057 18037 11069 18071
rect 11103 18068 11115 18071
rect 11238 18068 11244 18080
rect 11103 18040 11244 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 16132 18068 16160 18244
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 16301 18207 16359 18213
rect 16301 18173 16313 18207
rect 16347 18204 16359 18207
rect 16482 18204 16488 18216
rect 16347 18176 16488 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 16776 18204 16804 18312
rect 16942 18300 16948 18312
rect 17000 18300 17006 18352
rect 17037 18343 17095 18349
rect 17037 18309 17049 18343
rect 17083 18340 17095 18343
rect 17954 18340 17960 18352
rect 17083 18312 17960 18340
rect 17083 18309 17095 18312
rect 17037 18303 17095 18309
rect 17954 18300 17960 18312
rect 18012 18300 18018 18352
rect 18506 18300 18512 18352
rect 18564 18340 18570 18352
rect 19242 18340 19248 18352
rect 18564 18312 19248 18340
rect 18564 18300 18570 18312
rect 19242 18300 19248 18312
rect 19300 18300 19306 18352
rect 19610 18340 19616 18352
rect 19523 18312 19616 18340
rect 19610 18300 19616 18312
rect 19668 18300 19674 18352
rect 19705 18343 19763 18349
rect 19705 18309 19717 18343
rect 19751 18340 19763 18343
rect 20346 18340 20352 18352
rect 19751 18312 20352 18340
rect 19751 18309 19763 18312
rect 19705 18303 19763 18309
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 20925 18349 20953 18380
rect 20901 18343 20959 18349
rect 20901 18309 20913 18343
rect 20947 18309 20959 18343
rect 21376 18340 21404 18380
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 21508 18380 25268 18408
rect 21508 18368 21514 18380
rect 21376 18312 22416 18340
rect 20901 18303 20959 18309
rect 18414 18272 18420 18284
rect 17880 18244 18420 18272
rect 17880 18204 17908 18244
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 18877 18275 18935 18281
rect 18877 18272 18889 18275
rect 18748 18244 18889 18272
rect 18748 18232 18754 18244
rect 18877 18241 18889 18244
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18272 20315 18275
rect 20622 18272 20628 18284
rect 20303 18244 20628 18272
rect 20303 18241 20315 18244
rect 20257 18235 20315 18241
rect 16776 18176 17908 18204
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18012 18176 18057 18204
rect 18012 18164 18018 18176
rect 18966 18164 18972 18216
rect 19024 18204 19030 18216
rect 20272 18204 20300 18235
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 19024 18192 20017 18204
rect 20180 18192 20300 18204
rect 19024 18176 20300 18192
rect 20809 18207 20867 18213
rect 19024 18164 19030 18176
rect 19989 18164 20208 18176
rect 20809 18173 20821 18207
rect 20855 18204 20867 18207
rect 21450 18204 21456 18216
rect 20855 18192 20953 18204
rect 21008 18192 21456 18204
rect 20855 18176 21456 18192
rect 20855 18173 20867 18176
rect 20809 18167 20867 18173
rect 20925 18164 21036 18176
rect 21450 18164 21456 18176
rect 21508 18164 21514 18216
rect 21634 18164 21640 18216
rect 21692 18204 21698 18216
rect 22094 18204 22100 18216
rect 21692 18176 22100 18204
rect 21692 18164 21698 18176
rect 22094 18164 22100 18176
rect 22152 18164 22158 18216
rect 22388 18204 22416 18312
rect 22462 18300 22468 18352
rect 22520 18340 22526 18352
rect 23201 18343 23259 18349
rect 23201 18340 23213 18343
rect 22520 18312 23213 18340
rect 22520 18300 22526 18312
rect 23201 18309 23213 18312
rect 23247 18309 23259 18343
rect 23201 18303 23259 18309
rect 23293 18343 23351 18349
rect 23293 18309 23305 18343
rect 23339 18340 23351 18343
rect 24026 18340 24032 18352
rect 23339 18312 24032 18340
rect 23339 18309 23351 18312
rect 23293 18303 23351 18309
rect 24026 18300 24032 18312
rect 24084 18300 24090 18352
rect 24854 18340 24860 18352
rect 24815 18312 24860 18340
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 25240 18340 25268 18380
rect 25314 18368 25320 18420
rect 25372 18408 25378 18420
rect 25372 18380 27844 18408
rect 25372 18368 25378 18380
rect 25958 18340 25964 18352
rect 25240 18312 25964 18340
rect 25958 18300 25964 18312
rect 26016 18300 26022 18352
rect 26053 18343 26111 18349
rect 26053 18309 26065 18343
rect 26099 18340 26111 18343
rect 27522 18340 27528 18352
rect 26099 18312 27528 18340
rect 26099 18309 26111 18312
rect 26053 18303 26111 18309
rect 27522 18300 27528 18312
rect 27580 18300 27586 18352
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18272 25467 18275
rect 25682 18272 25688 18284
rect 25455 18244 25688 18272
rect 25455 18241 25467 18244
rect 25409 18235 25467 18241
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 26694 18232 26700 18284
rect 26752 18272 26758 18284
rect 27816 18281 27844 18380
rect 29914 18368 29920 18420
rect 29972 18408 29978 18420
rect 30837 18411 30895 18417
rect 30837 18408 30849 18411
rect 29972 18380 30849 18408
rect 29972 18368 29978 18380
rect 30837 18377 30849 18380
rect 30883 18377 30895 18411
rect 30837 18371 30895 18377
rect 28721 18343 28779 18349
rect 28721 18309 28733 18343
rect 28767 18340 28779 18343
rect 29730 18340 29736 18352
rect 28767 18312 29736 18340
rect 28767 18309 28779 18312
rect 28721 18303 28779 18309
rect 29730 18300 29736 18312
rect 29788 18300 29794 18352
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26752 18244 27169 18272
rect 26752 18232 26758 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27801 18275 27859 18281
rect 27801 18241 27813 18275
rect 27847 18241 27859 18275
rect 30098 18272 30104 18284
rect 30059 18244 30104 18272
rect 27801 18235 27859 18241
rect 30098 18232 30104 18244
rect 30156 18232 30162 18284
rect 30558 18232 30564 18284
rect 30616 18272 30622 18284
rect 30745 18275 30803 18281
rect 30745 18272 30757 18275
rect 30616 18244 30757 18272
rect 30616 18232 30622 18244
rect 30745 18241 30757 18244
rect 30791 18241 30803 18275
rect 30745 18235 30803 18241
rect 30834 18232 30840 18284
rect 30892 18272 30898 18284
rect 31389 18275 31447 18281
rect 31389 18272 31401 18275
rect 30892 18244 31401 18272
rect 30892 18232 30898 18244
rect 31389 18241 31401 18244
rect 31435 18241 31447 18275
rect 31389 18235 31447 18241
rect 24026 18204 24032 18216
rect 22388 18176 24032 18204
rect 24026 18164 24032 18176
rect 24084 18164 24090 18216
rect 24213 18207 24271 18213
rect 24213 18173 24225 18207
rect 24259 18173 24271 18207
rect 24213 18167 24271 18173
rect 16942 18096 16948 18148
rect 17000 18136 17006 18148
rect 19150 18136 19156 18148
rect 17000 18108 19156 18136
rect 17000 18096 17006 18108
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 20438 18136 20444 18148
rect 19893 18108 20444 18136
rect 12492 18040 16160 18068
rect 12492 18028 12498 18040
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 18230 18068 18236 18080
rect 16448 18040 18236 18068
rect 16448 18028 16454 18040
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 18414 18028 18420 18080
rect 18472 18068 18478 18080
rect 18874 18068 18880 18080
rect 18472 18040 18880 18068
rect 18472 18028 18478 18040
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 19893 18068 19921 18108
rect 20438 18096 20444 18108
rect 20496 18096 20502 18148
rect 21082 18136 21088 18148
rect 20732 18108 21088 18136
rect 19576 18040 19921 18068
rect 19576 18028 19582 18040
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20732 18068 20760 18108
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 21358 18136 21364 18148
rect 21319 18108 21364 18136
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 23474 18136 23480 18148
rect 22020 18108 23480 18136
rect 20220 18040 20760 18068
rect 20220 18028 20226 18040
rect 20806 18028 20812 18080
rect 20864 18068 20870 18080
rect 22020 18068 22048 18108
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 24228 18136 24256 18167
rect 24486 18164 24492 18216
rect 24544 18204 24550 18216
rect 24765 18207 24823 18213
rect 24765 18204 24777 18207
rect 24544 18176 24777 18204
rect 24544 18164 24550 18176
rect 24765 18173 24777 18176
rect 24811 18204 24823 18207
rect 26326 18204 26332 18216
rect 24811 18176 25912 18204
rect 26287 18176 26332 18204
rect 24811 18173 24823 18176
rect 24765 18167 24823 18173
rect 25038 18136 25044 18148
rect 24228 18108 25044 18136
rect 25038 18096 25044 18108
rect 25096 18096 25102 18148
rect 25884 18136 25912 18176
rect 26326 18164 26332 18176
rect 26384 18164 26390 18216
rect 28629 18207 28687 18213
rect 28629 18173 28641 18207
rect 28675 18204 28687 18207
rect 28994 18204 29000 18216
rect 28675 18176 29000 18204
rect 28675 18173 28687 18176
rect 28629 18167 28687 18173
rect 28994 18164 29000 18176
rect 29052 18164 29058 18216
rect 29641 18207 29699 18213
rect 29104 18176 29500 18204
rect 26510 18136 26516 18148
rect 25884 18108 26516 18136
rect 26510 18096 26516 18108
rect 26568 18096 26574 18148
rect 27246 18136 27252 18148
rect 27207 18108 27252 18136
rect 27246 18096 27252 18108
rect 27304 18096 27310 18148
rect 29104 18136 29132 18176
rect 29472 18148 29500 18176
rect 29641 18173 29653 18207
rect 29687 18204 29699 18207
rect 30006 18204 30012 18216
rect 29687 18176 30012 18204
rect 29687 18173 29699 18176
rect 29641 18167 29699 18173
rect 30006 18164 30012 18176
rect 30064 18164 30070 18216
rect 27356 18108 29132 18136
rect 20864 18040 22048 18068
rect 22097 18071 22155 18077
rect 20864 18028 20870 18040
rect 22097 18037 22109 18071
rect 22143 18068 22155 18071
rect 27356 18068 27384 18108
rect 29454 18096 29460 18148
rect 29512 18096 29518 18148
rect 22143 18040 27384 18068
rect 22143 18037 22155 18040
rect 22097 18031 22155 18037
rect 27614 18028 27620 18080
rect 27672 18068 27678 18080
rect 27893 18071 27951 18077
rect 27893 18068 27905 18071
rect 27672 18040 27905 18068
rect 27672 18028 27678 18040
rect 27893 18037 27905 18040
rect 27939 18037 27951 18071
rect 27893 18031 27951 18037
rect 28074 18028 28080 18080
rect 28132 18068 28138 18080
rect 29178 18068 29184 18080
rect 28132 18040 29184 18068
rect 28132 18028 28138 18040
rect 29178 18028 29184 18040
rect 29236 18028 29242 18080
rect 30190 18068 30196 18080
rect 30151 18040 30196 18068
rect 30190 18028 30196 18040
rect 30248 18028 30254 18080
rect 30374 18028 30380 18080
rect 30432 18068 30438 18080
rect 31481 18071 31539 18077
rect 31481 18068 31493 18071
rect 30432 18040 31493 18068
rect 30432 18028 30438 18040
rect 31481 18037 31493 18040
rect 31527 18037 31539 18071
rect 31481 18031 31539 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1936 17867 1994 17873
rect 1936 17833 1948 17867
rect 1982 17864 1994 17867
rect 1982 17836 8156 17864
rect 1982 17833 1994 17836
rect 1936 17827 1994 17833
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 6362 17796 6368 17808
rect 3467 17768 4108 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 2314 17728 2320 17740
rect 1719 17700 2320 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 2314 17688 2320 17700
rect 2372 17728 2378 17740
rect 3973 17731 4031 17737
rect 3973 17728 3985 17731
rect 2372 17700 3985 17728
rect 2372 17688 2378 17700
rect 3973 17697 3985 17700
rect 4019 17697 4031 17731
rect 4080 17728 4108 17768
rect 5276 17768 6368 17796
rect 4982 17728 4988 17740
rect 4080 17700 4988 17728
rect 3973 17691 4031 17697
rect 4982 17688 4988 17700
rect 5040 17728 5046 17740
rect 5276 17728 5304 17768
rect 6362 17756 6368 17768
rect 6420 17756 6426 17808
rect 8128 17796 8156 17836
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 14826 17864 14832 17876
rect 8352 17836 14832 17864
rect 8352 17824 8358 17836
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 16574 17864 16580 17876
rect 15304 17836 16580 17864
rect 8754 17796 8760 17808
rect 8128 17768 8760 17796
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 9398 17796 9404 17808
rect 8864 17768 9404 17796
rect 5040 17700 5304 17728
rect 5040 17688 5046 17700
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5592 17700 6009 17728
rect 5592 17688 5598 17700
rect 5997 17697 6009 17700
rect 6043 17697 6055 17731
rect 6454 17728 6460 17740
rect 6367 17700 6460 17728
rect 5997 17691 6055 17697
rect 6454 17688 6460 17700
rect 6512 17728 6518 17740
rect 6822 17728 6828 17740
rect 6512 17700 6828 17728
rect 6512 17688 6518 17700
rect 6822 17688 6828 17700
rect 6880 17728 6886 17740
rect 6880 17700 8340 17728
rect 6880 17688 6886 17700
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 3694 17592 3700 17604
rect 3174 17564 3700 17592
rect 3694 17552 3700 17564
rect 3752 17552 3758 17604
rect 4246 17592 4252 17604
rect 4207 17564 4252 17592
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 6730 17592 6736 17604
rect 6691 17564 6736 17592
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 8202 17592 8208 17604
rect 7958 17564 8208 17592
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 8312 17592 8340 17700
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 8864 17728 8892 17768
rect 9398 17756 9404 17768
rect 9456 17756 9462 17808
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 12894 17796 12900 17808
rect 11940 17768 12900 17796
rect 11940 17756 11946 17768
rect 12894 17756 12900 17768
rect 12952 17756 12958 17808
rect 15304 17796 15332 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 17954 17864 17960 17876
rect 16908 17836 17960 17864
rect 16908 17824 16914 17836
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 19610 17864 19616 17876
rect 18892 17836 19616 17864
rect 18414 17796 18420 17808
rect 13280 17768 15332 17796
rect 16132 17768 18420 17796
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 8628 17700 8892 17728
rect 9048 17700 9873 17728
rect 8628 17688 8634 17700
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 9048 17660 9076 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 13280 17728 13308 17768
rect 10008 17700 13308 17728
rect 13357 17731 13415 17737
rect 10008 17688 10014 17700
rect 13357 17697 13369 17731
rect 13403 17728 13415 17731
rect 14366 17728 14372 17740
rect 13403 17700 14372 17728
rect 13403 17697 13415 17700
rect 13357 17691 13415 17697
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 15381 17731 15439 17737
rect 15381 17697 15393 17731
rect 15427 17728 15439 17731
rect 15746 17728 15752 17740
rect 15427 17700 15752 17728
rect 15427 17697 15439 17700
rect 15381 17691 15439 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 16132 17737 16160 17768
rect 18414 17756 18420 17768
rect 18472 17756 18478 17808
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17697 16175 17731
rect 17034 17728 17040 17740
rect 16995 17700 17040 17728
rect 16117 17691 16175 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17728 17739 17731
rect 18782 17728 18788 17740
rect 17727 17700 18788 17728
rect 17727 17697 17739 17700
rect 17681 17691 17739 17697
rect 18782 17688 18788 17700
rect 18840 17728 18846 17740
rect 18892 17728 18920 17836
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 19886 17824 19892 17876
rect 19944 17864 19950 17876
rect 22005 17867 22063 17873
rect 22005 17864 22017 17867
rect 19944 17836 22017 17864
rect 19944 17824 19950 17836
rect 22005 17833 22017 17836
rect 22051 17833 22063 17867
rect 22005 17827 22063 17833
rect 24118 17824 24124 17876
rect 24176 17864 24182 17876
rect 24670 17864 24676 17876
rect 24176 17836 24676 17864
rect 24176 17824 24182 17836
rect 24670 17824 24676 17836
rect 24728 17824 24734 17876
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25869 17867 25927 17873
rect 25869 17864 25881 17867
rect 24912 17836 25881 17864
rect 24912 17824 24918 17836
rect 25869 17833 25881 17836
rect 25915 17833 25927 17867
rect 25869 17827 25927 17833
rect 25958 17824 25964 17876
rect 26016 17864 26022 17876
rect 30742 17864 30748 17876
rect 26016 17836 30748 17864
rect 26016 17824 26022 17836
rect 30742 17824 30748 17836
rect 30800 17824 30806 17876
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 20438 17796 20444 17808
rect 19024 17768 20444 17796
rect 19024 17756 19030 17768
rect 20438 17756 20444 17768
rect 20496 17756 20502 17808
rect 21358 17796 21364 17808
rect 20548 17768 20953 17796
rect 21319 17768 21364 17796
rect 20548 17728 20576 17768
rect 20925 17740 20953 17768
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 21910 17756 21916 17808
rect 21968 17796 21974 17808
rect 29822 17796 29828 17808
rect 21968 17768 29828 17796
rect 21968 17756 21974 17768
rect 29822 17756 29828 17768
rect 29880 17796 29886 17808
rect 31665 17799 31723 17805
rect 31665 17796 31677 17799
rect 29880 17768 31677 17796
rect 29880 17756 29886 17768
rect 31665 17765 31677 17768
rect 31711 17765 31723 17799
rect 31665 17759 31723 17765
rect 20806 17728 20812 17740
rect 18840 17700 18920 17728
rect 18984 17700 20576 17728
rect 20767 17700 20812 17728
rect 18840 17688 18846 17700
rect 8588 17632 9076 17660
rect 8588 17592 8616 17632
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 10594 17660 10600 17672
rect 9456 17632 10600 17660
rect 9456 17620 9462 17632
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12584 17632 12633 17660
rect 12584 17620 12590 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 13078 17660 13084 17672
rect 13039 17632 13084 17660
rect 12621 17623 12679 17629
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17660 18383 17663
rect 18414 17660 18420 17672
rect 18371 17632 18420 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 8312 17564 8616 17592
rect 9142 17595 9200 17601
rect 9142 17561 9154 17595
rect 9188 17592 9200 17595
rect 9766 17592 9772 17604
rect 9188 17564 9772 17592
rect 9188 17561 9200 17564
rect 9142 17555 9200 17561
rect 9766 17552 9772 17564
rect 9824 17552 9830 17604
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 10873 17595 10931 17601
rect 10873 17592 10885 17595
rect 10560 17564 10885 17592
rect 10560 17552 10566 17564
rect 10873 17561 10885 17564
rect 10919 17561 10931 17595
rect 12158 17592 12164 17604
rect 12098 17564 12164 17592
rect 10873 17555 10931 17561
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 14182 17592 14188 17604
rect 12452 17564 14188 17592
rect 1026 17484 1032 17536
rect 1084 17524 1090 17536
rect 2682 17524 2688 17536
rect 1084 17496 2688 17524
rect 1084 17484 1090 17496
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 4338 17524 4344 17536
rect 3936 17496 4344 17524
rect 3936 17484 3942 17496
rect 4338 17484 4344 17496
rect 4396 17524 4402 17536
rect 11790 17524 11796 17536
rect 4396 17496 11796 17524
rect 4396 17484 4402 17496
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 12452 17524 12480 17564
rect 14182 17552 14188 17564
rect 14240 17552 14246 17604
rect 14366 17592 14372 17604
rect 14327 17564 14372 17592
rect 14366 17552 14372 17564
rect 14424 17552 14430 17604
rect 14461 17595 14519 17601
rect 14461 17561 14473 17595
rect 14507 17561 14519 17595
rect 14461 17555 14519 17561
rect 12308 17496 12480 17524
rect 12308 17484 12314 17496
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 14476 17524 14504 17555
rect 14642 17552 14648 17604
rect 14700 17592 14706 17604
rect 15562 17592 15568 17604
rect 14700 17564 15568 17592
rect 14700 17552 14706 17564
rect 15562 17552 15568 17564
rect 15620 17552 15626 17604
rect 17770 17601 17776 17604
rect 16209 17595 16267 17601
rect 16209 17592 16221 17595
rect 16040 17564 16221 17592
rect 12584 17496 14504 17524
rect 12584 17484 12590 17496
rect 14826 17484 14832 17536
rect 14884 17524 14890 17536
rect 16040 17524 16068 17564
rect 16209 17561 16221 17564
rect 16255 17561 16267 17595
rect 17766 17592 17776 17601
rect 17731 17564 17776 17592
rect 16209 17555 16267 17561
rect 17766 17555 17776 17564
rect 17770 17552 17776 17555
rect 17828 17552 17834 17604
rect 17862 17552 17868 17604
rect 17920 17592 17926 17604
rect 18984 17592 19012 17700
rect 20806 17688 20812 17700
rect 20864 17688 20870 17740
rect 20925 17728 21036 17740
rect 26513 17731 26571 17737
rect 26513 17728 26525 17731
rect 20925 17712 26525 17728
rect 21008 17700 26525 17712
rect 26513 17697 26525 17700
rect 26559 17697 26571 17731
rect 26513 17691 26571 17697
rect 27246 17688 27252 17740
rect 27304 17728 27310 17740
rect 27525 17731 27583 17737
rect 27525 17728 27537 17731
rect 27304 17700 27537 17728
rect 27304 17688 27310 17700
rect 27525 17697 27537 17700
rect 27571 17728 27583 17731
rect 27890 17728 27896 17740
rect 27571 17700 27896 17728
rect 27571 17697 27583 17700
rect 27525 17691 27583 17697
rect 27890 17688 27896 17700
rect 27948 17688 27954 17740
rect 30190 17728 30196 17740
rect 28184 17700 30196 17728
rect 21913 17663 21971 17669
rect 21913 17629 21925 17663
rect 21959 17660 21971 17663
rect 22278 17660 22284 17672
rect 21959 17632 22284 17660
rect 21959 17629 21971 17632
rect 21913 17623 21971 17629
rect 22278 17620 22284 17632
rect 22336 17620 22342 17672
rect 22554 17660 22560 17672
rect 22515 17632 22560 17660
rect 22554 17620 22560 17632
rect 22612 17660 22618 17672
rect 23106 17660 23112 17672
rect 22612 17632 23112 17660
rect 22612 17620 22618 17632
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 23201 17663 23259 17669
rect 23201 17629 23213 17663
rect 23247 17660 23259 17663
rect 23290 17660 23296 17672
rect 23247 17632 23296 17660
rect 23247 17629 23259 17632
rect 23201 17623 23259 17629
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 23842 17660 23848 17672
rect 23803 17632 23848 17660
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 25777 17663 25835 17669
rect 25777 17629 25789 17663
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 26421 17663 26479 17669
rect 26421 17629 26433 17663
rect 26467 17660 26479 17663
rect 26786 17660 26792 17672
rect 26467 17632 26792 17660
rect 26467 17629 26479 17632
rect 26421 17623 26479 17629
rect 19518 17592 19524 17604
rect 17920 17564 19012 17592
rect 19479 17564 19524 17592
rect 17920 17552 17926 17564
rect 19518 17552 19524 17564
rect 19576 17552 19582 17604
rect 19613 17595 19671 17601
rect 19613 17561 19625 17595
rect 19659 17592 19671 17595
rect 20165 17595 20223 17601
rect 19659 17564 20116 17592
rect 19659 17561 19671 17564
rect 19613 17555 19671 17561
rect 14884 17496 16068 17524
rect 14884 17484 14890 17496
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17310 17524 17316 17536
rect 16632 17496 17316 17524
rect 16632 17484 16638 17496
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 19978 17524 19984 17536
rect 18012 17496 19984 17524
rect 18012 17484 18018 17496
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20088 17524 20116 17564
rect 20165 17561 20177 17595
rect 20211 17592 20223 17595
rect 20806 17592 20812 17604
rect 20211 17564 20812 17592
rect 20211 17561 20223 17564
rect 20165 17555 20223 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 20910 17595 20968 17601
rect 20910 17561 20922 17595
rect 20956 17592 20968 17595
rect 21174 17592 21180 17604
rect 20956 17564 21180 17592
rect 20956 17561 20968 17564
rect 20910 17555 20968 17561
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 24486 17592 24492 17604
rect 22020 17564 24492 17592
rect 22020 17524 22048 17564
rect 24486 17552 24492 17564
rect 24544 17552 24550 17604
rect 24670 17592 24676 17604
rect 24631 17564 24676 17592
rect 24670 17552 24676 17564
rect 24728 17552 24734 17604
rect 24762 17552 24768 17604
rect 24820 17592 24826 17604
rect 25317 17595 25375 17601
rect 24820 17564 24865 17592
rect 24820 17552 24826 17564
rect 25317 17561 25329 17595
rect 25363 17592 25375 17595
rect 25406 17592 25412 17604
rect 25363 17564 25412 17592
rect 25363 17561 25375 17564
rect 25317 17555 25375 17561
rect 25406 17552 25412 17564
rect 25464 17552 25470 17604
rect 20088 17496 22048 17524
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22649 17527 22707 17533
rect 22649 17524 22661 17527
rect 22152 17496 22661 17524
rect 22152 17484 22158 17496
rect 22649 17493 22661 17496
rect 22695 17493 22707 17527
rect 23290 17524 23296 17536
rect 23251 17496 23296 17524
rect 22649 17487 22707 17493
rect 23290 17484 23296 17496
rect 23348 17484 23354 17536
rect 23934 17524 23940 17536
rect 23895 17496 23940 17524
rect 23934 17484 23940 17496
rect 23992 17484 23998 17536
rect 24118 17484 24124 17536
rect 24176 17524 24182 17536
rect 25792 17524 25820 17623
rect 26786 17620 26792 17632
rect 26844 17660 26850 17672
rect 27062 17660 27068 17672
rect 26844 17632 27068 17660
rect 26844 17620 26850 17632
rect 27062 17620 27068 17632
rect 27120 17620 27126 17672
rect 27246 17592 27252 17604
rect 27207 17564 27252 17592
rect 27246 17552 27252 17564
rect 27304 17552 27310 17604
rect 27341 17595 27399 17601
rect 27341 17561 27353 17595
rect 27387 17592 27399 17595
rect 28184 17592 28212 17700
rect 30190 17688 30196 17700
rect 30248 17688 30254 17740
rect 37366 17728 37372 17740
rect 31128 17700 37372 17728
rect 31128 17672 31156 17700
rect 37366 17688 37372 17700
rect 37424 17688 37430 17740
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17629 28779 17663
rect 31110 17660 31116 17672
rect 31071 17632 31116 17660
rect 28721 17623 28779 17629
rect 27387 17564 28212 17592
rect 27387 17561 27399 17564
rect 27341 17555 27399 17561
rect 24176 17496 25820 17524
rect 24176 17484 24182 17496
rect 27430 17484 27436 17536
rect 27488 17524 27494 17536
rect 28736 17524 28764 17623
rect 31110 17620 31116 17632
rect 31168 17620 31174 17672
rect 31573 17663 31631 17669
rect 31573 17629 31585 17663
rect 31619 17660 31631 17663
rect 34514 17660 34520 17672
rect 31619 17632 34520 17660
rect 31619 17629 31631 17632
rect 31573 17623 31631 17629
rect 34514 17620 34520 17632
rect 34572 17620 34578 17672
rect 29822 17592 29828 17604
rect 29783 17564 29828 17592
rect 29822 17552 29828 17564
rect 29880 17552 29886 17604
rect 29917 17595 29975 17601
rect 29917 17561 29929 17595
rect 29963 17561 29975 17595
rect 29917 17555 29975 17561
rect 27488 17496 28764 17524
rect 27488 17484 27494 17496
rect 28810 17484 28816 17536
rect 28868 17524 28874 17536
rect 29932 17524 29960 17555
rect 30006 17552 30012 17604
rect 30064 17592 30070 17604
rect 30466 17592 30472 17604
rect 30064 17564 30472 17592
rect 30064 17552 30070 17564
rect 30466 17552 30472 17564
rect 30524 17552 30530 17604
rect 30374 17524 30380 17536
rect 28868 17496 28913 17524
rect 29932 17496 30380 17524
rect 28868 17484 28874 17496
rect 30374 17484 30380 17496
rect 30432 17484 30438 17536
rect 30650 17484 30656 17536
rect 30708 17524 30714 17536
rect 30929 17527 30987 17533
rect 30929 17524 30941 17527
rect 30708 17496 30941 17524
rect 30708 17484 30714 17496
rect 30929 17493 30941 17496
rect 30975 17493 30987 17527
rect 30929 17487 30987 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2682 17280 2688 17332
rect 2740 17320 2746 17332
rect 11422 17320 11428 17332
rect 2740 17292 5028 17320
rect 2740 17280 2746 17292
rect 566 17212 572 17264
rect 624 17252 630 17264
rect 4338 17252 4344 17264
rect 624 17224 3082 17252
rect 4299 17224 4344 17252
rect 624 17212 630 17224
rect 4338 17212 4344 17224
rect 4396 17212 4402 17264
rect 4890 17252 4896 17264
rect 4851 17224 4896 17252
rect 4890 17212 4896 17224
rect 4948 17212 4954 17264
rect 5000 17261 5028 17292
rect 6932 17292 11428 17320
rect 6932 17261 6960 17292
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 16574 17320 16580 17332
rect 11756 17292 14044 17320
rect 11756 17280 11762 17292
rect 4985 17255 5043 17261
rect 4985 17221 4997 17255
rect 5031 17221 5043 17255
rect 4985 17215 5043 17221
rect 6917 17255 6975 17261
rect 6917 17221 6929 17255
rect 6963 17221 6975 17255
rect 8754 17252 8760 17264
rect 8142 17224 8760 17252
rect 6917 17215 6975 17221
rect 8754 17212 8760 17224
rect 8812 17212 8818 17264
rect 9030 17252 9036 17264
rect 8864 17224 9036 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17153 1639 17187
rect 2314 17184 2320 17196
rect 2275 17156 2320 17184
rect 1581 17147 1639 17153
rect 1596 17116 1624 17147
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 8864 17193 8892 17224
rect 9030 17212 9036 17224
rect 9088 17212 9094 17264
rect 9122 17212 9128 17264
rect 9180 17252 9186 17264
rect 9180 17224 9225 17252
rect 9180 17212 9186 17224
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 11974 17252 11980 17264
rect 9456 17224 9614 17252
rect 11935 17224 11980 17252
rect 9456 17212 9462 17224
rect 11974 17212 11980 17224
rect 12032 17212 12038 17264
rect 14016 17252 14044 17292
rect 15120 17292 16580 17320
rect 14093 17255 14151 17261
rect 14093 17252 14105 17255
rect 14016 17224 14105 17252
rect 14093 17221 14105 17224
rect 14139 17221 14151 17255
rect 14093 17215 14151 17221
rect 6641 17187 6699 17193
rect 6641 17184 6653 17187
rect 6512 17156 6653 17184
rect 6512 17144 6518 17156
rect 6641 17153 6653 17156
rect 6687 17153 6699 17187
rect 6641 17147 6699 17153
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 10962 17184 10968 17196
rect 10652 17156 10968 17184
rect 10652 17144 10658 17156
rect 10962 17144 10968 17156
rect 11020 17184 11026 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11020 17156 11713 17184
rect 11020 17144 11026 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 13110 17156 13860 17184
rect 11701 17147 11759 17153
rect 2593 17119 2651 17125
rect 2593 17116 2605 17119
rect 1596 17088 2268 17116
rect 2240 16992 2268 17088
rect 2424 17088 2605 17116
rect 2424 16992 2452 17088
rect 2593 17085 2605 17088
rect 2639 17085 2651 17119
rect 5166 17116 5172 17128
rect 5127 17088 5172 17116
rect 2593 17079 2651 17085
rect 5166 17076 5172 17088
rect 5224 17116 5230 17128
rect 5224 17088 10456 17116
rect 5224 17076 5230 17088
rect 8389 17051 8447 17057
rect 8389 17017 8401 17051
rect 8435 17048 8447 17051
rect 8570 17048 8576 17060
rect 8435 17020 8576 17048
rect 8435 17017 8447 17020
rect 8389 17011 8447 17017
rect 8570 17008 8576 17020
rect 8628 17008 8634 17060
rect 2222 16980 2228 16992
rect 2183 16952 2228 16980
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 2406 16940 2412 16992
rect 2464 16940 2470 16992
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 5074 16980 5080 16992
rect 4948 16952 5080 16980
rect 4948 16940 4954 16952
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 10134 16980 10140 16992
rect 8812 16952 10140 16980
rect 8812 16940 8818 16952
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10428 16980 10456 17088
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10836 17088 10885 17116
rect 10836 17076 10842 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 13354 17116 13360 17128
rect 11480 17088 13360 17116
rect 11480 17076 11486 17088
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17116 13507 17119
rect 13722 17116 13728 17128
rect 13495 17088 13728 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 13832 17048 13860 17156
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 15120 17116 15148 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 16868 17292 17540 17320
rect 15378 17252 15384 17264
rect 15339 17224 15384 17252
rect 15378 17212 15384 17224
rect 15436 17212 15442 17264
rect 16301 17255 16359 17261
rect 16301 17221 16313 17255
rect 16347 17252 16359 17255
rect 16868 17252 16896 17292
rect 17034 17252 17040 17264
rect 16347 17224 16896 17252
rect 16995 17224 17040 17252
rect 16347 17221 16359 17224
rect 16301 17215 16359 17221
rect 17034 17212 17040 17224
rect 17092 17212 17098 17264
rect 17512 17252 17540 17292
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18506 17320 18512 17332
rect 17644 17292 18512 17320
rect 17644 17280 17650 17292
rect 18506 17280 18512 17292
rect 18564 17280 18570 17332
rect 18598 17280 18604 17332
rect 18656 17280 18662 17332
rect 23934 17320 23940 17332
rect 18800 17292 23940 17320
rect 18616 17252 18644 17280
rect 18800 17261 18828 17292
rect 23934 17280 23940 17292
rect 23992 17280 23998 17332
rect 24026 17280 24032 17332
rect 24084 17320 24090 17332
rect 24084 17292 24129 17320
rect 24084 17280 24090 17292
rect 25130 17280 25136 17332
rect 25188 17320 25194 17332
rect 27430 17320 27436 17332
rect 25188 17292 27436 17320
rect 25188 17280 25194 17292
rect 27430 17280 27436 17292
rect 27488 17280 27494 17332
rect 27522 17280 27528 17332
rect 27580 17320 27586 17332
rect 28445 17323 28503 17329
rect 28445 17320 28457 17323
rect 27580 17292 28457 17320
rect 27580 17280 27586 17292
rect 28445 17289 28457 17292
rect 28491 17289 28503 17323
rect 30558 17320 30564 17332
rect 28445 17283 28503 17289
rect 28966 17292 30564 17320
rect 17512 17224 18644 17252
rect 18785 17255 18843 17261
rect 18785 17221 18797 17255
rect 18831 17221 18843 17255
rect 18785 17215 18843 17221
rect 19058 17212 19064 17264
rect 19116 17252 19122 17264
rect 19705 17255 19763 17261
rect 19705 17252 19717 17255
rect 19116 17224 19717 17252
rect 19116 17212 19122 17224
rect 19705 17221 19717 17224
rect 19751 17252 19763 17255
rect 20070 17252 20076 17264
rect 19751 17224 20076 17252
rect 19751 17221 19763 17224
rect 19705 17215 19763 17221
rect 20070 17212 20076 17224
rect 20128 17212 20134 17264
rect 20533 17255 20591 17261
rect 20533 17221 20545 17255
rect 20579 17252 20591 17255
rect 20898 17252 20904 17264
rect 20579 17224 20904 17252
rect 20579 17221 20591 17224
rect 20533 17215 20591 17221
rect 20898 17212 20904 17224
rect 20956 17212 20962 17264
rect 22186 17252 22192 17264
rect 22147 17224 22192 17252
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22281 17255 22339 17261
rect 22281 17221 22293 17255
rect 22327 17252 22339 17255
rect 23106 17252 23112 17264
rect 22327 17224 23112 17252
rect 22327 17221 22339 17224
rect 22281 17215 22339 17221
rect 23106 17212 23112 17224
rect 23164 17212 23170 17264
rect 23385 17255 23443 17261
rect 23385 17221 23397 17255
rect 23431 17252 23443 17255
rect 24857 17255 24915 17261
rect 24857 17252 24869 17255
rect 23431 17224 24869 17252
rect 23431 17221 23443 17224
rect 23385 17215 23443 17221
rect 24857 17221 24869 17224
rect 24903 17221 24915 17255
rect 24857 17215 24915 17221
rect 24946 17212 24952 17264
rect 25004 17252 25010 17264
rect 25409 17255 25467 17261
rect 25409 17252 25421 17255
rect 25004 17224 25421 17252
rect 25004 17212 25010 17224
rect 25409 17221 25421 17224
rect 25455 17221 25467 17255
rect 25409 17215 25467 17221
rect 27341 17255 27399 17261
rect 27341 17221 27353 17255
rect 27387 17252 27399 17255
rect 28534 17252 28540 17264
rect 27387 17224 28540 17252
rect 27387 17221 27399 17224
rect 27341 17215 27399 17221
rect 28534 17212 28540 17224
rect 28592 17212 28598 17264
rect 20162 17184 20168 17196
rect 19536 17156 20168 17184
rect 14047 17088 15148 17116
rect 15289 17119 15347 17125
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 16574 17116 16580 17128
rect 15335 17088 16580 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 17862 17116 17868 17128
rect 16991 17088 17868 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 14553 17051 14611 17057
rect 13832 17020 14504 17048
rect 11974 16980 11980 16992
rect 10428 16952 11980 16980
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 14366 16980 14372 16992
rect 12124 16952 14372 16980
rect 12124 16940 12130 16952
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 14476 16980 14504 17020
rect 14553 17017 14565 17051
rect 14599 17048 14611 17051
rect 15194 17048 15200 17060
rect 14599 17020 15200 17048
rect 14599 17017 14611 17020
rect 14553 17011 14611 17017
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 15470 17008 15476 17060
rect 15528 17048 15534 17060
rect 16960 17048 16988 17079
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18012 17088 18057 17116
rect 18012 17076 18018 17088
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 18693 17119 18751 17125
rect 18693 17116 18705 17119
rect 18564 17088 18705 17116
rect 18564 17076 18570 17088
rect 18693 17085 18705 17088
rect 18739 17085 18751 17119
rect 18693 17079 18751 17085
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 19536 17116 19564 17156
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 21910 17184 21916 17196
rect 21376 17156 21916 17184
rect 20441 17119 20499 17125
rect 18932 17088 19564 17116
rect 19621 17088 19741 17116
rect 18932 17076 18938 17088
rect 15528 17020 16988 17048
rect 15528 17008 15534 17020
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 17586 17048 17592 17060
rect 17184 17020 17592 17048
rect 17184 17008 17190 17020
rect 17586 17008 17592 17020
rect 17644 17008 17650 17060
rect 17770 17008 17776 17060
rect 17828 17048 17834 17060
rect 19621 17048 19649 17088
rect 17828 17020 19649 17048
rect 19713 17048 19741 17088
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 21376 17116 21404 17156
rect 21910 17144 21916 17156
rect 21968 17144 21974 17196
rect 22830 17144 22836 17196
rect 22888 17184 22894 17196
rect 22888 17156 22933 17184
rect 22888 17144 22894 17156
rect 23198 17144 23204 17196
rect 23256 17184 23262 17196
rect 23293 17187 23351 17193
rect 23293 17184 23305 17187
rect 23256 17156 23305 17184
rect 23256 17144 23262 17156
rect 23293 17153 23305 17156
rect 23339 17153 23351 17187
rect 23934 17184 23940 17196
rect 23895 17156 23940 17184
rect 23293 17147 23351 17153
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 25869 17187 25927 17193
rect 25869 17153 25881 17187
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17184 28411 17187
rect 28966 17184 28994 17292
rect 30558 17280 30564 17292
rect 30616 17280 30622 17332
rect 29457 17255 29515 17261
rect 29457 17221 29469 17255
rect 29503 17252 29515 17255
rect 31570 17252 31576 17264
rect 29503 17224 31576 17252
rect 29503 17221 29515 17224
rect 29457 17215 29515 17221
rect 31570 17212 31576 17224
rect 31628 17212 31634 17264
rect 28399 17156 28994 17184
rect 30469 17187 30527 17193
rect 28399 17153 28411 17156
rect 28353 17147 28411 17153
rect 30469 17153 30481 17187
rect 30515 17184 30527 17187
rect 31110 17184 31116 17196
rect 30515 17156 31116 17184
rect 30515 17153 30527 17156
rect 30469 17147 30527 17153
rect 20487 17088 21404 17116
rect 21453 17119 21511 17125
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 21453 17085 21465 17119
rect 21499 17116 21511 17119
rect 22646 17116 22652 17128
rect 21499 17088 22652 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 23952 17116 23980 17144
rect 24765 17119 24823 17125
rect 23952 17088 24716 17116
rect 24688 17048 24716 17088
rect 24765 17085 24777 17119
rect 24811 17116 24823 17119
rect 25130 17116 25136 17128
rect 24811 17088 25136 17116
rect 24811 17085 24823 17088
rect 24765 17079 24823 17085
rect 25130 17076 25136 17088
rect 25188 17076 25194 17128
rect 25884 17048 25912 17147
rect 26234 17076 26240 17128
rect 26292 17116 26298 17128
rect 27246 17116 27252 17128
rect 26292 17088 27252 17116
rect 26292 17076 26298 17088
rect 27246 17076 27252 17088
rect 27304 17076 27310 17128
rect 27522 17116 27528 17128
rect 27483 17088 27528 17116
rect 27522 17076 27528 17088
rect 27580 17076 27586 17128
rect 27706 17076 27712 17128
rect 27764 17116 27770 17128
rect 28368 17116 28396 17147
rect 31110 17144 31116 17156
rect 31168 17144 31174 17196
rect 37737 17187 37795 17193
rect 37737 17184 37749 17187
rect 35866 17156 37749 17184
rect 27764 17088 28396 17116
rect 27764 17076 27770 17088
rect 28994 17076 29000 17128
rect 29052 17116 29058 17128
rect 29365 17119 29423 17125
rect 29365 17116 29377 17119
rect 29052 17088 29377 17116
rect 29052 17076 29058 17088
rect 29365 17085 29377 17088
rect 29411 17116 29423 17119
rect 30098 17116 30104 17128
rect 29411 17088 30104 17116
rect 29411 17085 29423 17088
rect 29365 17079 29423 17085
rect 30098 17076 30104 17088
rect 30156 17076 30162 17128
rect 19713 17020 24164 17048
rect 24688 17020 25912 17048
rect 17828 17008 17834 17020
rect 24026 16980 24032 16992
rect 14476 16952 24032 16980
rect 24026 16940 24032 16952
rect 24084 16940 24090 16992
rect 24136 16980 24164 17020
rect 25961 16983 26019 16989
rect 25961 16980 25973 16983
rect 24136 16952 25973 16980
rect 25961 16949 25973 16952
rect 26007 16949 26019 16983
rect 27264 16980 27292 17076
rect 28902 17008 28908 17060
rect 28960 17048 28966 17060
rect 29917 17051 29975 17057
rect 29917 17048 29929 17051
rect 28960 17020 29929 17048
rect 28960 17008 28966 17020
rect 29917 17017 29929 17020
rect 29963 17017 29975 17051
rect 29917 17011 29975 17017
rect 30742 17008 30748 17060
rect 30800 17048 30806 17060
rect 35866 17048 35894 17156
rect 37737 17153 37749 17156
rect 37783 17153 37795 17187
rect 37737 17147 37795 17153
rect 37458 17116 37464 17128
rect 37419 17088 37464 17116
rect 37458 17076 37464 17088
rect 37516 17076 37522 17128
rect 30800 17020 35894 17048
rect 30800 17008 30806 17020
rect 30561 16983 30619 16989
rect 30561 16980 30573 16983
rect 27264 16952 30573 16980
rect 25961 16943 26019 16949
rect 30561 16949 30573 16952
rect 30607 16949 30619 16983
rect 30561 16943 30619 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 4065 16779 4123 16785
rect 4065 16745 4077 16779
rect 4111 16776 4123 16779
rect 5810 16776 5816 16788
rect 4111 16748 5816 16776
rect 4111 16745 4123 16748
rect 4065 16739 4123 16745
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6086 16736 6092 16788
rect 6144 16776 6150 16788
rect 6144 16748 8248 16776
rect 6144 16736 6150 16748
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 1673 16643 1731 16649
rect 1673 16640 1685 16643
rect 1636 16612 1685 16640
rect 1636 16600 1642 16612
rect 1673 16609 1685 16612
rect 1719 16640 1731 16643
rect 2314 16640 2320 16652
rect 1719 16612 2320 16640
rect 1719 16609 1731 16612
rect 1673 16603 1731 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 2682 16600 2688 16652
rect 2740 16640 2746 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 2740 16612 4353 16640
rect 2740 16600 2746 16612
rect 4341 16609 4353 16612
rect 4387 16640 4399 16643
rect 4614 16640 4620 16652
rect 4387 16612 4620 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 4614 16600 4620 16612
rect 4672 16640 4678 16652
rect 5350 16640 5356 16652
rect 4672 16612 5356 16640
rect 4672 16600 4678 16612
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 6546 16640 6552 16652
rect 6507 16612 6552 16640
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6825 16643 6883 16649
rect 6825 16609 6837 16643
rect 6871 16640 6883 16643
rect 7558 16640 7564 16652
rect 6871 16612 7564 16640
rect 6871 16609 6883 16612
rect 6825 16603 6883 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8220 16640 8248 16748
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 16942 16776 16948 16788
rect 9916 16748 12434 16776
rect 9916 16736 9922 16748
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8352 16680 10732 16708
rect 8352 16668 8358 16680
rect 8754 16640 8760 16652
rect 8220 16612 8760 16640
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 9674 16600 9680 16652
rect 9732 16640 9738 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9732 16612 9873 16640
rect 9732 16600 9738 16612
rect 9861 16609 9873 16612
rect 9907 16640 9919 16643
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 9907 16612 10609 16640
rect 9907 16609 9919 16612
rect 9861 16603 9919 16609
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10704 16640 10732 16680
rect 11974 16668 11980 16720
rect 12032 16708 12038 16720
rect 12406 16708 12434 16748
rect 14936 16748 16948 16776
rect 14936 16708 14964 16748
rect 16942 16736 16948 16748
rect 17000 16736 17006 16788
rect 17034 16736 17040 16788
rect 17092 16776 17098 16788
rect 22922 16776 22928 16788
rect 17092 16748 22928 16776
rect 17092 16736 17098 16748
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 23017 16779 23075 16785
rect 23017 16745 23029 16779
rect 23063 16776 23075 16779
rect 23106 16776 23112 16788
rect 23063 16748 23112 16776
rect 23063 16745 23075 16748
rect 23017 16739 23075 16745
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 23198 16736 23204 16788
rect 23256 16776 23262 16788
rect 23661 16779 23719 16785
rect 23661 16776 23673 16779
rect 23256 16748 23673 16776
rect 23256 16736 23262 16748
rect 23661 16745 23673 16748
rect 23707 16745 23719 16779
rect 23661 16739 23719 16745
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 27246 16776 27252 16788
rect 24084 16748 27252 16776
rect 24084 16736 24090 16748
rect 27246 16736 27252 16748
rect 27304 16736 27310 16788
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 28350 16776 28356 16788
rect 27488 16748 28356 16776
rect 27488 16736 27494 16748
rect 28350 16736 28356 16748
rect 28408 16736 28414 16788
rect 33502 16736 33508 16788
rect 33560 16776 33566 16788
rect 38197 16779 38255 16785
rect 38197 16776 38209 16779
rect 33560 16748 38209 16776
rect 33560 16736 33566 16748
rect 38197 16745 38209 16748
rect 38243 16745 38255 16779
rect 38197 16739 38255 16745
rect 12032 16680 12304 16708
rect 12406 16680 14964 16708
rect 12032 16668 12038 16680
rect 12276 16640 12304 16680
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 28810 16708 28816 16720
rect 15436 16680 28816 16708
rect 15436 16668 15442 16680
rect 28810 16668 28816 16680
rect 28868 16668 28874 16720
rect 29638 16668 29644 16720
rect 29696 16708 29702 16720
rect 30834 16708 30840 16720
rect 29696 16680 30840 16708
rect 29696 16668 29702 16680
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 10704 16612 12112 16640
rect 12276 16612 15485 16640
rect 10597 16603 10655 16609
rect 3418 16532 3424 16584
rect 3476 16572 3482 16584
rect 8570 16572 8576 16584
rect 3476 16544 4384 16572
rect 8531 16544 8576 16572
rect 3476 16532 3482 16544
rect 4356 16516 4384 16544
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 12084 16572 12112 16612
rect 15473 16609 15485 16612
rect 15519 16640 15531 16643
rect 15562 16640 15568 16652
rect 15519 16612 15568 16640
rect 15519 16609 15531 16612
rect 15473 16603 15531 16609
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 16632 16612 17325 16640
rect 16632 16600 16638 16612
rect 17313 16609 17325 16612
rect 17359 16640 17371 16643
rect 17494 16640 17500 16652
rect 17359 16612 17500 16640
rect 17359 16609 17371 16612
rect 17313 16603 17371 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 17770 16640 17776 16652
rect 17644 16612 17776 16640
rect 17644 16600 17650 16612
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 19702 16640 19708 16652
rect 18248 16612 19708 16640
rect 12084 16544 12296 16572
rect 1949 16507 2007 16513
rect 1949 16473 1961 16507
rect 1995 16473 2007 16507
rect 4062 16504 4068 16516
rect 3174 16476 4068 16504
rect 1949 16467 2007 16473
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 1964 16436 1992 16467
rect 4062 16464 4068 16476
rect 4120 16464 4126 16516
rect 4338 16464 4344 16516
rect 4396 16464 4402 16516
rect 4617 16507 4675 16513
rect 4617 16473 4629 16507
rect 4663 16473 4675 16507
rect 6730 16504 6736 16516
rect 5842 16476 6736 16504
rect 4617 16467 4675 16473
rect 1820 16408 1992 16436
rect 1820 16396 1826 16408
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3292 16408 3433 16436
rect 3292 16396 3298 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 4632 16436 4660 16467
rect 6730 16464 6736 16476
rect 6788 16464 6794 16516
rect 8202 16504 8208 16516
rect 8050 16476 8208 16504
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 8662 16464 8668 16516
rect 8720 16504 8726 16516
rect 9030 16504 9036 16516
rect 8720 16476 9036 16504
rect 8720 16464 8726 16476
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 9125 16507 9183 16513
rect 9125 16473 9137 16507
rect 9171 16504 9183 16507
rect 9766 16504 9772 16516
rect 9171 16476 9772 16504
rect 9171 16473 9183 16476
rect 9125 16467 9183 16473
rect 9766 16464 9772 16476
rect 9824 16504 9830 16516
rect 10134 16504 10140 16516
rect 9824 16476 10140 16504
rect 9824 16464 9830 16476
rect 10134 16464 10140 16476
rect 10192 16464 10198 16516
rect 10502 16464 10508 16516
rect 10560 16504 10566 16516
rect 10778 16504 10784 16516
rect 10560 16476 10784 16504
rect 10560 16464 10566 16476
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 10870 16464 10876 16516
rect 10928 16504 10934 16516
rect 12158 16504 12164 16516
rect 10928 16476 10973 16504
rect 12098 16476 12164 16504
rect 10928 16464 10934 16476
rect 12158 16464 12164 16476
rect 12216 16464 12222 16516
rect 12268 16504 12296 16544
rect 12342 16532 12348 16584
rect 12400 16572 12406 16584
rect 12400 16544 12940 16572
rect 12400 16532 12406 16544
rect 12434 16504 12440 16516
rect 12268 16476 12440 16504
rect 12434 16464 12440 16476
rect 12492 16464 12498 16516
rect 12621 16507 12679 16513
rect 12621 16473 12633 16507
rect 12667 16504 12679 16507
rect 12802 16504 12808 16516
rect 12667 16476 12808 16504
rect 12667 16473 12679 16476
rect 12621 16467 12679 16473
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 12912 16504 12940 16544
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13906 16572 13912 16584
rect 13136 16544 13912 16572
rect 13136 16532 13142 16544
rect 13906 16532 13912 16544
rect 13964 16532 13970 16584
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14461 16575 14519 16581
rect 14461 16572 14473 16575
rect 14148 16544 14473 16572
rect 14148 16532 14154 16544
rect 14461 16541 14473 16544
rect 14507 16572 14519 16575
rect 14642 16572 14648 16584
rect 14507 16544 14648 16572
rect 14507 16541 14519 16544
rect 14461 16535 14519 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12912 16476 13369 16504
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 13357 16467 13415 16473
rect 13630 16464 13636 16516
rect 13688 16504 13694 16516
rect 14553 16507 14611 16513
rect 14553 16504 14565 16507
rect 13688 16476 14565 16504
rect 13688 16464 13694 16476
rect 14553 16473 14565 16476
rect 14599 16473 14611 16507
rect 15194 16504 15200 16516
rect 15155 16476 15200 16504
rect 14553 16467 14611 16473
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15289 16507 15347 16513
rect 15289 16473 15301 16507
rect 15335 16504 15347 16507
rect 17310 16504 17316 16516
rect 15335 16476 17316 16504
rect 15335 16473 15347 16476
rect 15289 16467 15347 16473
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 17405 16507 17463 16513
rect 17405 16473 17417 16507
rect 17451 16504 17463 16507
rect 18248 16504 18276 16612
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 20530 16640 20536 16652
rect 19852 16612 20536 16640
rect 19852 16600 19858 16612
rect 20530 16600 20536 16612
rect 20588 16640 20594 16652
rect 20588 16612 20668 16640
rect 20588 16600 20594 16612
rect 18598 16532 18604 16584
rect 18656 16572 18662 16584
rect 20640 16581 20668 16612
rect 20714 16600 20720 16652
rect 20772 16640 20778 16652
rect 21453 16643 21511 16649
rect 20772 16612 20817 16640
rect 20772 16600 20778 16612
rect 21453 16609 21465 16643
rect 21499 16640 21511 16643
rect 22278 16640 22284 16652
rect 21499 16612 22284 16640
rect 21499 16609 21511 16612
rect 21453 16603 21511 16609
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 20625 16575 20683 16581
rect 18656 16544 19380 16572
rect 18656 16532 18662 16544
rect 17451 16476 18276 16504
rect 18325 16507 18383 16513
rect 17451 16473 17463 16476
rect 17405 16467 17463 16473
rect 18325 16473 18337 16507
rect 18371 16504 18383 16507
rect 19058 16504 19064 16516
rect 18371 16476 19064 16504
rect 18371 16473 18383 16476
rect 18325 16467 18383 16473
rect 19058 16464 19064 16476
rect 19116 16464 19122 16516
rect 4706 16436 4712 16448
rect 4619 16408 4712 16436
rect 3421 16399 3479 16405
rect 4706 16396 4712 16408
rect 4764 16436 4770 16448
rect 4982 16436 4988 16448
rect 4764 16408 4988 16436
rect 4764 16396 4770 16408
rect 4982 16396 4988 16408
rect 5040 16396 5046 16448
rect 6089 16439 6147 16445
rect 6089 16405 6101 16439
rect 6135 16436 6147 16439
rect 6178 16436 6184 16448
rect 6135 16408 6184 16436
rect 6135 16405 6147 16408
rect 6089 16399 6147 16405
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 14458 16436 14464 16448
rect 8904 16408 14464 16436
rect 8904 16396 8910 16408
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 15010 16396 15016 16448
rect 15068 16436 15074 16448
rect 16298 16436 16304 16448
rect 15068 16408 16304 16436
rect 15068 16396 15074 16408
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16482 16396 16488 16448
rect 16540 16436 16546 16448
rect 18874 16436 18880 16448
rect 16540 16408 18880 16436
rect 16540 16396 16546 16408
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 19352 16436 19380 16544
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 22480 16572 22508 16603
rect 22738 16600 22744 16652
rect 22796 16640 22802 16652
rect 22796 16612 22968 16640
rect 22796 16600 22802 16612
rect 22830 16572 22836 16584
rect 22480 16544 22836 16572
rect 20625 16535 20683 16541
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 22940 16581 22968 16612
rect 26068 16612 27108 16640
rect 22925 16575 22983 16581
rect 22925 16541 22937 16575
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 23382 16532 23388 16584
rect 23440 16572 23446 16584
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 23440 16544 23581 16572
rect 23440 16532 23446 16544
rect 23569 16541 23581 16544
rect 23615 16572 23627 16575
rect 23658 16572 23664 16584
rect 23615 16544 23664 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 23658 16532 23664 16544
rect 23716 16532 23722 16584
rect 26068 16574 26096 16612
rect 25884 16572 26096 16574
rect 25608 16546 26096 16572
rect 27080 16572 27108 16612
rect 27890 16600 27896 16652
rect 27948 16640 27954 16652
rect 27948 16612 29040 16640
rect 27948 16600 27954 16612
rect 27614 16572 27620 16584
rect 25608 16544 25912 16546
rect 27080 16544 27620 16572
rect 19518 16504 19524 16516
rect 19479 16476 19524 16504
rect 19518 16464 19524 16476
rect 19576 16464 19582 16516
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16504 19671 16507
rect 19978 16504 19984 16516
rect 19659 16476 19984 16504
rect 19659 16473 19671 16476
rect 19613 16467 19671 16473
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 20165 16507 20223 16513
rect 20165 16473 20177 16507
rect 20211 16504 20223 16507
rect 20346 16504 20352 16516
rect 20211 16476 20352 16504
rect 20211 16473 20223 16476
rect 20165 16467 20223 16473
rect 20346 16464 20352 16476
rect 20404 16464 20410 16516
rect 21082 16464 21088 16516
rect 21140 16504 21146 16516
rect 21545 16507 21603 16513
rect 21545 16504 21557 16507
rect 21140 16476 21557 16504
rect 21140 16464 21146 16476
rect 21545 16473 21557 16476
rect 21591 16473 21603 16507
rect 24670 16504 24676 16516
rect 21545 16467 21603 16473
rect 22756 16476 24676 16504
rect 22094 16436 22100 16448
rect 19352 16408 22100 16436
rect 22094 16396 22100 16408
rect 22152 16436 22158 16448
rect 22756 16436 22784 16476
rect 24670 16464 24676 16476
rect 24728 16464 24734 16516
rect 24765 16507 24823 16513
rect 24765 16473 24777 16507
rect 24811 16504 24823 16507
rect 25608 16504 25636 16544
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 27706 16532 27712 16584
rect 27764 16572 27770 16584
rect 28368 16581 28396 16612
rect 28353 16575 28411 16581
rect 27764 16544 27809 16572
rect 27764 16532 27770 16544
rect 28353 16541 28365 16575
rect 28399 16541 28411 16575
rect 28353 16535 28411 16541
rect 28442 16532 28448 16584
rect 28500 16572 28506 16584
rect 29012 16581 29040 16612
rect 28997 16575 29055 16581
rect 28500 16544 28545 16572
rect 28500 16532 28506 16544
rect 28997 16541 29009 16575
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 29086 16532 29092 16584
rect 29144 16572 29150 16584
rect 29748 16581 29776 16680
rect 30834 16668 30840 16680
rect 30892 16668 30898 16720
rect 30282 16600 30288 16652
rect 30340 16640 30346 16652
rect 37182 16640 37188 16652
rect 30340 16612 30420 16640
rect 30340 16600 30346 16612
rect 30392 16581 30420 16612
rect 31036 16612 37188 16640
rect 31036 16581 31064 16612
rect 37182 16600 37188 16612
rect 37240 16600 37246 16652
rect 29733 16575 29791 16581
rect 29144 16544 29189 16572
rect 29144 16532 29150 16544
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 30377 16575 30435 16581
rect 30377 16541 30389 16575
rect 30423 16541 30435 16575
rect 30377 16535 30435 16541
rect 31021 16575 31079 16581
rect 31021 16541 31033 16575
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 24811 16476 25636 16504
rect 25685 16507 25743 16513
rect 24811 16473 24823 16476
rect 24765 16467 24823 16473
rect 25685 16473 25697 16507
rect 25731 16504 25743 16507
rect 26050 16504 26056 16516
rect 25731 16476 26056 16504
rect 25731 16473 25743 16476
rect 25685 16467 25743 16473
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 26234 16504 26240 16516
rect 26195 16476 26240 16504
rect 26234 16464 26240 16476
rect 26292 16464 26298 16516
rect 26329 16507 26387 16513
rect 26329 16473 26341 16507
rect 26375 16473 26387 16507
rect 26329 16467 26387 16473
rect 22152 16408 22784 16436
rect 22152 16396 22158 16408
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 25866 16436 25872 16448
rect 22888 16408 25872 16436
rect 22888 16396 22894 16408
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 26344 16436 26372 16467
rect 27062 16464 27068 16516
rect 27120 16504 27126 16516
rect 27249 16507 27307 16513
rect 27249 16504 27261 16507
rect 27120 16476 27261 16504
rect 27120 16464 27126 16476
rect 27249 16473 27261 16476
rect 27295 16473 27307 16507
rect 29825 16507 29883 16513
rect 29825 16504 29837 16507
rect 27249 16467 27307 16473
rect 27586 16476 29837 16504
rect 27586 16436 27614 16476
rect 29825 16473 29837 16476
rect 29871 16473 29883 16507
rect 38102 16504 38108 16516
rect 38063 16476 38108 16504
rect 29825 16467 29883 16473
rect 38102 16464 38108 16476
rect 38160 16464 38166 16516
rect 27798 16436 27804 16448
rect 26344 16408 27614 16436
rect 27759 16408 27804 16436
rect 27798 16396 27804 16408
rect 27856 16396 27862 16448
rect 28074 16396 28080 16448
rect 28132 16436 28138 16448
rect 29730 16436 29736 16448
rect 28132 16408 29736 16436
rect 28132 16396 28138 16408
rect 29730 16396 29736 16408
rect 29788 16396 29794 16448
rect 30466 16436 30472 16448
rect 30427 16408 30472 16436
rect 30466 16396 30472 16408
rect 30524 16396 30530 16448
rect 31110 16436 31116 16448
rect 31071 16408 31116 16436
rect 31110 16396 31116 16408
rect 31168 16396 31174 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 5399 16235 5457 16241
rect 5399 16232 5411 16235
rect 5224 16204 5411 16232
rect 5224 16192 5230 16204
rect 5399 16201 5411 16204
rect 5445 16201 5457 16235
rect 7098 16232 7104 16244
rect 7059 16204 7104 16232
rect 5399 16195 5457 16201
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 10502 16232 10508 16244
rect 7944 16204 10508 16232
rect 4338 16124 4344 16176
rect 4396 16164 4402 16176
rect 7650 16164 7656 16176
rect 4396 16136 7656 16164
rect 4396 16124 4402 16136
rect 7650 16124 7656 16136
rect 7708 16124 7714 16176
rect 7944 16173 7972 16204
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10796 16204 13308 16232
rect 7929 16167 7987 16173
rect 7929 16133 7941 16167
rect 7975 16133 7987 16167
rect 7929 16127 7987 16133
rect 9582 16124 9588 16176
rect 9640 16164 9646 16176
rect 10796 16164 10824 16204
rect 10962 16164 10968 16176
rect 9640 16136 10824 16164
rect 10923 16136 10968 16164
rect 9640 16124 9646 16136
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11330 16164 11336 16176
rect 11112 16136 11336 16164
rect 11112 16124 11118 16136
rect 11330 16124 11336 16136
rect 11388 16164 11394 16176
rect 11974 16164 11980 16176
rect 11388 16136 11980 16164
rect 11388 16124 11394 16136
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 12434 16124 12440 16176
rect 12492 16124 12498 16176
rect 13280 16164 13308 16204
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 16390 16232 16396 16244
rect 13596 16204 16396 16232
rect 13596 16192 13602 16204
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 26237 16235 26295 16241
rect 26237 16232 26249 16235
rect 17045 16204 26249 16232
rect 15010 16164 15016 16176
rect 13280 16136 15016 16164
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 15378 16124 15384 16176
rect 15436 16164 15442 16176
rect 16301 16167 16359 16173
rect 15436 16136 15481 16164
rect 15436 16124 15442 16136
rect 16301 16133 16313 16167
rect 16347 16164 16359 16167
rect 16758 16164 16764 16176
rect 16347 16136 16764 16164
rect 16347 16133 16359 16136
rect 16301 16127 16359 16133
rect 16758 16124 16764 16136
rect 16816 16124 16822 16176
rect 17045 16173 17073 16204
rect 26237 16201 26249 16204
rect 26283 16201 26295 16235
rect 27246 16232 27252 16244
rect 27207 16204 27252 16232
rect 26237 16195 26295 16201
rect 27246 16192 27252 16204
rect 27304 16192 27310 16244
rect 31110 16232 31116 16244
rect 27908 16204 31116 16232
rect 17030 16167 17088 16173
rect 17030 16133 17042 16167
rect 17076 16133 17088 16167
rect 17030 16127 17088 16133
rect 17402 16124 17408 16176
rect 17460 16164 17466 16176
rect 18598 16164 18604 16176
rect 17460 16136 18604 16164
rect 17460 16124 17466 16136
rect 18598 16124 18604 16136
rect 18656 16124 18662 16176
rect 18782 16164 18788 16176
rect 18743 16136 18788 16164
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16164 18935 16167
rect 19242 16164 19248 16176
rect 18923 16136 19248 16164
rect 18923 16133 18935 16136
rect 18877 16127 18935 16133
rect 19242 16124 19248 16136
rect 19300 16124 19306 16176
rect 19794 16164 19800 16176
rect 19444 16136 19800 16164
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2682 16096 2688 16108
rect 2643 16068 2688 16096
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 3007 16000 4016 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 1765 15895 1823 15901
rect 1765 15861 1777 15895
rect 1811 15892 1823 15895
rect 3694 15892 3700 15904
rect 1811 15864 3700 15892
rect 1811 15861 1823 15864
rect 1765 15855 1823 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 3988 15892 4016 16000
rect 4080 15960 4108 16082
rect 4246 16056 4252 16108
rect 4304 16096 4310 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4304 16068 5181 16096
rect 4304 16056 4310 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 7006 16096 7012 16108
rect 6967 16068 7012 16096
rect 5169 16059 5227 16065
rect 7006 16056 7012 16068
rect 7064 16056 7070 16108
rect 4706 16028 4712 16040
rect 4667 16000 4712 16028
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 7653 16031 7711 16037
rect 7653 16028 7665 16031
rect 6604 16000 7665 16028
rect 6604 15988 6610 16000
rect 7653 15997 7665 16000
rect 7699 16028 7711 16031
rect 8662 16028 8668 16040
rect 7699 16000 8668 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 9048 15960 9076 16082
rect 9490 16056 9496 16108
rect 9548 16096 9554 16108
rect 10042 16096 10048 16108
rect 9548 16068 10048 16096
rect 9548 16056 9554 16068
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10229 16099 10287 16105
rect 10229 16096 10241 16099
rect 10192 16068 10241 16096
rect 10192 16056 10198 16068
rect 10229 16065 10241 16068
rect 10275 16065 10287 16099
rect 10980 16096 11008 16124
rect 19444 16108 19472 16136
rect 19794 16124 19800 16136
rect 19852 16124 19858 16176
rect 19978 16124 19984 16176
rect 20036 16164 20042 16176
rect 20625 16167 20683 16173
rect 20625 16164 20637 16167
rect 20036 16136 20637 16164
rect 20036 16124 20042 16136
rect 20625 16133 20637 16136
rect 20671 16133 20683 16167
rect 20625 16127 20683 16133
rect 20898 16124 20904 16176
rect 20956 16164 20962 16176
rect 21269 16167 21327 16173
rect 21269 16164 21281 16167
rect 20956 16136 21281 16164
rect 20956 16124 20962 16136
rect 21269 16133 21281 16136
rect 21315 16133 21327 16167
rect 22094 16164 22100 16176
rect 22055 16136 22100 16164
rect 21269 16127 21327 16133
rect 22094 16124 22100 16136
rect 22152 16124 22158 16176
rect 22189 16167 22247 16173
rect 22189 16133 22201 16167
rect 22235 16164 22247 16167
rect 23198 16164 23204 16176
rect 22235 16136 23204 16164
rect 22235 16133 22247 16136
rect 22189 16127 22247 16133
rect 23198 16124 23204 16136
rect 23256 16124 23262 16176
rect 24302 16164 24308 16176
rect 24263 16136 24308 16164
rect 24302 16124 24308 16136
rect 24360 16124 24366 16176
rect 24762 16124 24768 16176
rect 24820 16164 24826 16176
rect 27798 16164 27804 16176
rect 24820 16136 27804 16164
rect 24820 16124 24826 16136
rect 27798 16124 27804 16136
rect 27856 16124 27862 16176
rect 11514 16096 11520 16108
rect 10980 16068 11520 16096
rect 10229 16059 10287 16065
rect 11514 16056 11520 16068
rect 11572 16096 11578 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11572 16068 11713 16096
rect 11572 16056 11578 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13964 16068 14197 16096
rect 13964 16056 13970 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 19426 16056 19432 16108
rect 19484 16056 19490 16108
rect 19610 16056 19616 16108
rect 19668 16096 19674 16108
rect 19889 16099 19947 16105
rect 19889 16096 19901 16099
rect 19668 16068 19901 16096
rect 19668 16056 19674 16068
rect 19889 16065 19901 16068
rect 19935 16096 19947 16099
rect 20438 16096 20444 16108
rect 19935 16068 20444 16096
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16096 20591 16099
rect 20714 16096 20720 16108
rect 20579 16068 20720 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 23382 16096 23388 16108
rect 21185 16089 21243 16095
rect 21185 16055 21197 16089
rect 21231 16086 21243 16089
rect 21231 16058 21312 16086
rect 21231 16055 21243 16058
rect 21185 16049 21243 16055
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 11054 16028 11060 16040
rect 9723 16000 11060 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 11054 15988 11060 16000
rect 11112 15988 11118 16040
rect 11330 15988 11336 16040
rect 11388 16028 11394 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11388 16000 11989 16028
rect 11388 15988 11394 16000
rect 11977 15997 11989 16000
rect 12023 16028 12035 16031
rect 13630 16028 13636 16040
rect 12023 16000 13636 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 14366 16028 14372 16040
rect 13780 16000 13825 16028
rect 14327 16000 14372 16028
rect 13780 15988 13786 16000
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 15997 15347 16031
rect 16942 16028 16948 16040
rect 16903 16000 16948 16028
rect 15289 15991 15347 15997
rect 10962 15960 10968 15972
rect 4080 15932 7788 15960
rect 9048 15932 10968 15960
rect 5258 15892 5264 15904
rect 3988 15864 5264 15892
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 6638 15892 6644 15904
rect 6236 15864 6644 15892
rect 6236 15852 6242 15864
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 7760 15892 7788 15932
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 13998 15920 14004 15972
rect 14056 15960 14062 15972
rect 14826 15960 14832 15972
rect 14056 15932 14832 15960
rect 14056 15920 14062 15932
rect 14826 15920 14832 15932
rect 14884 15920 14890 15972
rect 15304 15960 15332 15991
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 17402 16028 17408 16040
rect 17144 16000 17408 16028
rect 17144 15960 17172 16000
rect 17402 15988 17408 16000
rect 17460 16028 17466 16040
rect 17862 16028 17868 16040
rect 17460 16000 17868 16028
rect 17460 15988 17466 16000
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18012 16000 18057 16028
rect 18012 15988 18018 16000
rect 18874 15988 18880 16040
rect 18932 16028 18938 16040
rect 18932 16000 20714 16028
rect 18932 15988 18938 16000
rect 15304 15932 17172 15960
rect 17218 15920 17224 15972
rect 17276 15960 17282 15972
rect 19337 15963 19395 15969
rect 19337 15960 19349 15963
rect 17276 15932 19349 15960
rect 17276 15920 17282 15932
rect 19337 15929 19349 15932
rect 19383 15929 19395 15963
rect 20686 15960 20714 16000
rect 20898 15988 20904 16040
rect 20956 16028 20962 16040
rect 20956 16016 21128 16028
rect 21284 16016 21312 16058
rect 22940 16068 23388 16096
rect 21634 16028 21640 16040
rect 20956 16000 21312 16016
rect 20956 15988 20962 16000
rect 21100 15988 21312 16000
rect 21376 16000 21640 16028
rect 21376 15960 21404 16000
rect 21634 15988 21640 16000
rect 21692 16028 21698 16040
rect 21910 16028 21916 16040
rect 21692 16000 21916 16028
rect 21692 15988 21698 16000
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 22940 16028 22968 16068
rect 23382 16056 23388 16068
rect 23440 16056 23446 16108
rect 23569 16099 23627 16105
rect 23569 16065 23581 16099
rect 23615 16065 23627 16099
rect 23569 16059 23627 16065
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16065 24271 16099
rect 24854 16096 24860 16108
rect 24815 16068 24860 16096
rect 24213 16059 24271 16065
rect 23106 16028 23112 16040
rect 22152 16000 22968 16028
rect 23067 16000 23112 16028
rect 22152 15988 22158 16000
rect 23106 15988 23112 16000
rect 23164 15988 23170 16040
rect 23584 16028 23612 16059
rect 23216 16000 23612 16028
rect 19337 15923 19395 15929
rect 19444 15932 20116 15960
rect 20686 15932 21404 15960
rect 13170 15892 13176 15904
rect 7760 15864 13176 15892
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 19444 15892 19472 15932
rect 19978 15892 19984 15904
rect 13320 15864 19472 15892
rect 19939 15864 19984 15892
rect 13320 15852 13326 15864
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20088 15892 20116 15932
rect 21818 15920 21824 15972
rect 21876 15960 21882 15972
rect 23216 15960 23244 16000
rect 24228 15960 24256 16059
rect 24854 16056 24860 16068
rect 24912 16056 24918 16108
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25501 16099 25559 16105
rect 25501 16096 25513 16099
rect 25096 16068 25513 16096
rect 25096 16056 25102 16068
rect 25501 16065 25513 16068
rect 25547 16065 25559 16099
rect 26142 16096 26148 16108
rect 26103 16068 26148 16096
rect 25501 16059 25559 16065
rect 26142 16056 26148 16068
rect 26200 16056 26206 16108
rect 27157 16099 27215 16105
rect 27157 16065 27169 16099
rect 27203 16096 27215 16099
rect 27246 16096 27252 16108
rect 27203 16068 27252 16096
rect 27203 16065 27215 16068
rect 27157 16059 27215 16065
rect 27246 16056 27252 16068
rect 27304 16056 27310 16108
rect 24670 15988 24676 16040
rect 24728 16028 24734 16040
rect 27908 16028 27936 16204
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 31570 16232 31576 16244
rect 31531 16204 31576 16232
rect 31570 16192 31576 16204
rect 31628 16192 31634 16244
rect 35897 16235 35955 16241
rect 35897 16201 35909 16235
rect 35943 16232 35955 16235
rect 38010 16232 38016 16244
rect 35943 16204 38016 16232
rect 35943 16201 35955 16204
rect 35897 16195 35955 16201
rect 38010 16192 38016 16204
rect 38068 16192 38074 16244
rect 28258 16164 28264 16176
rect 28219 16136 28264 16164
rect 28258 16124 28264 16136
rect 28316 16124 28322 16176
rect 29178 16164 29184 16176
rect 29139 16136 29184 16164
rect 29178 16124 29184 16136
rect 29236 16124 29242 16176
rect 29546 16124 29552 16176
rect 29604 16164 29610 16176
rect 29733 16167 29791 16173
rect 29733 16164 29745 16167
rect 29604 16136 29745 16164
rect 29604 16124 29610 16136
rect 29733 16133 29745 16136
rect 29779 16133 29791 16167
rect 29733 16127 29791 16133
rect 29825 16167 29883 16173
rect 29825 16133 29837 16167
rect 29871 16164 29883 16167
rect 30466 16164 30472 16176
rect 29871 16136 30472 16164
rect 29871 16133 29883 16136
rect 29825 16127 29883 16133
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 30834 16096 30840 16108
rect 30795 16068 30840 16096
rect 30834 16056 30840 16068
rect 30892 16056 30898 16108
rect 31110 16056 31116 16108
rect 31168 16096 31174 16108
rect 31481 16099 31539 16105
rect 31481 16096 31493 16099
rect 31168 16068 31493 16096
rect 31168 16056 31174 16068
rect 31481 16065 31493 16068
rect 31527 16065 31539 16099
rect 31481 16059 31539 16065
rect 35894 16056 35900 16108
rect 35952 16096 35958 16108
rect 36081 16099 36139 16105
rect 36081 16096 36093 16099
rect 35952 16068 36093 16096
rect 35952 16056 35958 16068
rect 36081 16065 36093 16068
rect 36127 16065 36139 16099
rect 36081 16059 36139 16065
rect 24728 16000 27936 16028
rect 28169 16031 28227 16037
rect 24728 15988 24734 16000
rect 28169 15997 28181 16031
rect 28215 16028 28227 16031
rect 28994 16028 29000 16040
rect 28215 16000 29000 16028
rect 28215 15997 28227 16000
rect 28169 15991 28227 15997
rect 28994 15988 29000 16000
rect 29052 15988 29058 16040
rect 30006 16028 30012 16040
rect 29919 16000 30012 16028
rect 30006 15988 30012 16000
rect 30064 15988 30070 16040
rect 21876 15932 23244 15960
rect 23584 15932 24256 15960
rect 21876 15920 21882 15932
rect 23584 15892 23612 15932
rect 24486 15920 24492 15972
rect 24544 15960 24550 15972
rect 25593 15963 25651 15969
rect 25593 15960 25605 15963
rect 24544 15932 25605 15960
rect 24544 15920 24550 15932
rect 25593 15929 25605 15932
rect 25639 15929 25651 15963
rect 25593 15923 25651 15929
rect 25866 15920 25872 15972
rect 25924 15960 25930 15972
rect 28074 15960 28080 15972
rect 25924 15932 28080 15960
rect 25924 15920 25930 15932
rect 28074 15920 28080 15932
rect 28132 15920 28138 15972
rect 29086 15960 29092 15972
rect 28368 15932 29092 15960
rect 20088 15864 23612 15892
rect 23658 15852 23664 15904
rect 23716 15892 23722 15904
rect 24946 15892 24952 15904
rect 23716 15864 23761 15892
rect 24907 15864 24952 15892
rect 23716 15852 23722 15864
rect 24946 15852 24952 15864
rect 25004 15852 25010 15904
rect 25130 15852 25136 15904
rect 25188 15892 25194 15904
rect 28368 15892 28396 15932
rect 29086 15920 29092 15932
rect 29144 15920 29150 15972
rect 29178 15920 29184 15972
rect 29236 15960 29242 15972
rect 30024 15960 30052 15988
rect 29236 15932 30052 15960
rect 29236 15920 29242 15932
rect 25188 15864 28396 15892
rect 25188 15852 25194 15864
rect 28442 15852 28448 15904
rect 28500 15892 28506 15904
rect 30929 15895 30987 15901
rect 30929 15892 30941 15895
rect 28500 15864 30941 15892
rect 28500 15852 28506 15864
rect 30929 15861 30941 15864
rect 30975 15861 30987 15895
rect 30929 15855 30987 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 934 15648 940 15700
rect 992 15688 998 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 992 15660 3341 15688
rect 992 15648 998 15660
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 4062 15688 4068 15700
rect 3975 15660 4068 15688
rect 3329 15651 3387 15657
rect 4062 15648 4068 15660
rect 4120 15688 4126 15700
rect 11057 15691 11115 15697
rect 4120 15660 11008 15688
rect 4120 15648 4126 15660
rect 4246 15620 4252 15632
rect 3988 15592 4252 15620
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15552 1642 15564
rect 3988 15552 4016 15592
rect 4246 15580 4252 15592
rect 4304 15620 4310 15632
rect 9214 15620 9220 15632
rect 4304 15592 4936 15620
rect 4304 15580 4310 15592
rect 4908 15561 4936 15592
rect 6656 15592 9220 15620
rect 1636 15524 4016 15552
rect 4893 15555 4951 15561
rect 1636 15512 1642 15524
rect 4893 15521 4905 15555
rect 4939 15521 4951 15555
rect 4893 15515 4951 15521
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15552 5687 15555
rect 5718 15552 5724 15564
rect 5675 15524 5724 15552
rect 5675 15521 5687 15524
rect 5629 15515 5687 15521
rect 5718 15512 5724 15524
rect 5776 15512 5782 15564
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6656 15552 6684 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 10980 15620 11008 15660
rect 11057 15657 11069 15691
rect 11103 15688 11115 15691
rect 11422 15688 11428 15700
rect 11103 15660 11428 15688
rect 11103 15657 11115 15660
rect 11057 15651 11115 15657
rect 11422 15648 11428 15660
rect 11480 15648 11486 15700
rect 12342 15688 12348 15700
rect 11532 15660 12348 15688
rect 11532 15620 11560 15660
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 22094 15688 22100 15700
rect 13688 15660 22100 15688
rect 13688 15648 13694 15660
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 26142 15688 26148 15700
rect 22244 15660 26148 15688
rect 22244 15648 22250 15660
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 26418 15648 26424 15700
rect 26476 15688 26482 15700
rect 26513 15691 26571 15697
rect 26513 15688 26525 15691
rect 26476 15660 26525 15688
rect 26476 15648 26482 15660
rect 26513 15657 26525 15660
rect 26559 15657 26571 15691
rect 27154 15688 27160 15700
rect 27115 15660 27160 15688
rect 26513 15651 26571 15657
rect 27154 15648 27160 15660
rect 27212 15648 27218 15700
rect 27614 15648 27620 15700
rect 27672 15688 27678 15700
rect 33502 15688 33508 15700
rect 27672 15660 33508 15688
rect 27672 15648 27678 15660
rect 33502 15648 33508 15660
rect 33560 15648 33566 15700
rect 10980 15592 11560 15620
rect 13078 15580 13084 15632
rect 13136 15620 13142 15632
rect 16025 15623 16083 15629
rect 13136 15592 14412 15620
rect 13136 15580 13142 15592
rect 6420 15524 6684 15552
rect 6420 15512 6426 15524
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 7340 15524 7389 15552
rect 7340 15512 7346 15524
rect 7377 15521 7389 15524
rect 7423 15552 7435 15555
rect 7926 15552 7932 15564
rect 7423 15524 7932 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 8662 15512 8668 15564
rect 8720 15552 8726 15564
rect 9309 15555 9367 15561
rect 9309 15552 9321 15555
rect 8720 15524 9321 15552
rect 8720 15512 8726 15524
rect 9309 15521 9321 15524
rect 9355 15552 9367 15555
rect 9674 15552 9680 15564
rect 9355 15524 9680 15552
rect 9355 15521 9367 15524
rect 9309 15515 9367 15521
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 10042 15512 10048 15564
rect 10100 15552 10106 15564
rect 10100 15524 10916 15552
rect 10100 15512 10106 15524
rect 5350 15484 5356 15496
rect 5311 15456 5356 15484
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 8754 15484 8760 15496
rect 8619 15456 8760 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 1857 15419 1915 15425
rect 1857 15385 1869 15419
rect 1903 15385 1915 15419
rect 4062 15416 4068 15428
rect 3082 15388 4068 15416
rect 1857 15379 1915 15385
rect 1872 15348 1900 15379
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 4157 15419 4215 15425
rect 4157 15385 4169 15419
rect 4203 15416 4215 15419
rect 4614 15416 4620 15428
rect 4203 15388 4620 15416
rect 4203 15385 4215 15388
rect 4157 15379 4215 15385
rect 4614 15376 4620 15388
rect 4672 15376 4678 15428
rect 5902 15376 5908 15428
rect 5960 15416 5966 15428
rect 5960 15388 6118 15416
rect 5960 15376 5966 15388
rect 7650 15376 7656 15428
rect 7708 15416 7714 15428
rect 7929 15419 7987 15425
rect 7929 15416 7941 15419
rect 7708 15388 7941 15416
rect 7708 15376 7714 15388
rect 7929 15385 7941 15388
rect 7975 15385 7987 15419
rect 7929 15379 7987 15385
rect 8021 15419 8079 15425
rect 8021 15385 8033 15419
rect 8067 15416 8079 15419
rect 8110 15416 8116 15428
rect 8067 15388 8116 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 8110 15376 8116 15388
rect 8168 15376 8174 15428
rect 8386 15376 8392 15428
rect 8444 15416 8450 15428
rect 8588 15416 8616 15447
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 8444 15388 8616 15416
rect 8444 15376 8450 15388
rect 8662 15376 8668 15428
rect 8720 15416 8726 15428
rect 9490 15416 9496 15428
rect 8720 15388 9496 15416
rect 8720 15376 8726 15388
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 9585 15419 9643 15425
rect 9585 15385 9597 15419
rect 9631 15416 9643 15419
rect 9631 15388 9996 15416
rect 9631 15385 9643 15388
rect 9585 15379 9643 15385
rect 3234 15348 3240 15360
rect 1872 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 3694 15308 3700 15360
rect 3752 15348 3758 15360
rect 6362 15348 6368 15360
rect 3752 15320 6368 15348
rect 3752 15308 3758 15320
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 9674 15348 9680 15360
rect 6696 15320 9680 15348
rect 6696 15308 6702 15320
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 9968 15348 9996 15388
rect 10042 15376 10048 15428
rect 10100 15376 10106 15428
rect 10888 15416 10916 15524
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11330 15552 11336 15564
rect 11112 15524 11336 15552
rect 11112 15512 11118 15524
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11514 15552 11520 15564
rect 11475 15524 11520 15552
rect 11514 15512 11520 15524
rect 11572 15552 11578 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 11572 15524 14289 15552
rect 11572 15512 11578 15524
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 14384 15552 14412 15592
rect 16025 15589 16037 15623
rect 16071 15620 16083 15623
rect 16298 15620 16304 15632
rect 16071 15592 16304 15620
rect 16071 15589 16083 15592
rect 16025 15583 16083 15589
rect 16298 15580 16304 15592
rect 16356 15580 16362 15632
rect 16390 15580 16396 15632
rect 16448 15620 16454 15632
rect 22738 15620 22744 15632
rect 16448 15592 22744 15620
rect 16448 15580 16454 15592
rect 22738 15580 22744 15592
rect 22796 15580 22802 15632
rect 24578 15580 24584 15632
rect 24636 15580 24642 15632
rect 26970 15580 26976 15632
rect 27028 15620 27034 15632
rect 27798 15620 27804 15632
rect 27028 15592 27804 15620
rect 27028 15580 27034 15592
rect 27798 15580 27804 15592
rect 27856 15580 27862 15632
rect 28905 15623 28963 15629
rect 28905 15589 28917 15623
rect 28951 15620 28963 15623
rect 31386 15620 31392 15632
rect 28951 15592 31392 15620
rect 28951 15589 28963 15592
rect 28905 15583 28963 15589
rect 31386 15580 31392 15592
rect 31444 15580 31450 15632
rect 14384 15524 17440 15552
rect 14277 15515 14335 15521
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17412 15484 17440 15524
rect 17494 15512 17500 15564
rect 17552 15552 17558 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17552 15524 17877 15552
rect 17552 15512 17558 15524
rect 17865 15521 17877 15524
rect 17911 15552 17923 15555
rect 18877 15555 18935 15561
rect 17911 15524 18744 15552
rect 17911 15521 17923 15524
rect 17865 15515 17923 15521
rect 17586 15484 17592 15496
rect 17276 15456 17321 15484
rect 17412 15456 17592 15484
rect 17276 15444 17282 15456
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 18716 15484 18744 15524
rect 18877 15521 18889 15555
rect 18923 15552 18935 15555
rect 18966 15552 18972 15564
rect 18923 15524 18972 15552
rect 18923 15521 18935 15524
rect 18877 15515 18935 15521
rect 18966 15512 18972 15524
rect 19024 15512 19030 15564
rect 19076 15552 19334 15564
rect 19076 15536 22221 15552
rect 19076 15484 19104 15536
rect 19306 15524 22221 15536
rect 18716 15456 19104 15484
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 20254 15484 20260 15496
rect 19475 15456 20260 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20530 15444 20536 15496
rect 20588 15484 20594 15496
rect 20806 15484 20812 15496
rect 20588 15456 20812 15484
rect 20588 15444 20594 15456
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 22193 15484 22221 15524
rect 22278 15512 22284 15564
rect 22336 15552 22342 15564
rect 23937 15555 23995 15561
rect 22336 15524 23796 15552
rect 22336 15512 22342 15524
rect 22646 15484 22652 15496
rect 22193 15456 22652 15484
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23768 15484 23796 15524
rect 23937 15521 23949 15555
rect 23983 15552 23995 15555
rect 24596 15552 24624 15580
rect 23983 15524 24624 15552
rect 25317 15555 25375 15561
rect 23983 15521 23995 15524
rect 23937 15515 23995 15521
rect 25317 15521 25329 15555
rect 25363 15552 25375 15555
rect 27522 15552 27528 15564
rect 25363 15524 27528 15552
rect 25363 15521 25375 15524
rect 25317 15515 25375 15521
rect 27522 15512 27528 15524
rect 27580 15512 27586 15564
rect 28350 15552 28356 15564
rect 28311 15524 28356 15552
rect 28350 15512 28356 15524
rect 28408 15512 28414 15564
rect 37734 15552 37740 15564
rect 35866 15524 37740 15552
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23768 15456 24593 15484
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 25961 15487 26019 15493
rect 25961 15453 25973 15487
rect 26007 15484 26019 15487
rect 26326 15484 26332 15496
rect 26007 15456 26332 15484
rect 26007 15453 26019 15456
rect 25961 15447 26019 15453
rect 26326 15444 26332 15456
rect 26384 15444 26390 15496
rect 26421 15487 26479 15493
rect 26421 15453 26433 15487
rect 26467 15484 26479 15487
rect 26970 15484 26976 15496
rect 26467 15456 26976 15484
rect 26467 15453 26479 15456
rect 26421 15447 26479 15453
rect 26970 15444 26976 15456
rect 27028 15444 27034 15496
rect 27065 15487 27123 15493
rect 27065 15453 27077 15487
rect 27111 15453 27123 15487
rect 27065 15447 27123 15453
rect 11790 15416 11796 15428
rect 10888 15388 11796 15416
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 11882 15376 11888 15428
rect 11940 15376 11946 15428
rect 13018 15388 13952 15416
rect 11146 15348 11152 15360
rect 9968 15320 11152 15348
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11900 15348 11928 15376
rect 13265 15351 13323 15357
rect 13265 15348 13277 15351
rect 11900 15320 13277 15348
rect 13265 15317 13277 15320
rect 13311 15317 13323 15351
rect 13924 15348 13952 15388
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 14553 15419 14611 15425
rect 14553 15416 14565 15419
rect 14056 15388 14565 15416
rect 14056 15376 14062 15388
rect 14553 15385 14565 15388
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 14642 15376 14648 15428
rect 14700 15416 14706 15428
rect 16574 15416 16580 15428
rect 14700 15388 15042 15416
rect 16535 15388 16580 15416
rect 14700 15376 14706 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 16669 15419 16727 15425
rect 16669 15385 16681 15419
rect 16715 15385 16727 15419
rect 16669 15379 16727 15385
rect 17957 15419 18015 15425
rect 17957 15385 17969 15419
rect 18003 15416 18015 15419
rect 20070 15416 20076 15428
rect 18003 15388 20076 15416
rect 18003 15385 18015 15388
rect 17957 15379 18015 15385
rect 16390 15348 16396 15360
rect 13924 15320 16396 15348
rect 13265 15311 13323 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 16684 15348 16712 15379
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 20625 15419 20683 15425
rect 20625 15385 20637 15419
rect 20671 15385 20683 15419
rect 20625 15379 20683 15385
rect 21361 15419 21419 15425
rect 21361 15385 21373 15419
rect 21407 15385 21419 15419
rect 21361 15379 21419 15385
rect 18874 15348 18880 15360
rect 16684 15320 18880 15348
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19150 15308 19156 15360
rect 19208 15348 19214 15360
rect 19521 15351 19579 15357
rect 19521 15348 19533 15351
rect 19208 15320 19533 15348
rect 19208 15308 19214 15320
rect 19521 15317 19533 15320
rect 19567 15317 19579 15351
rect 19521 15311 19579 15317
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 20640 15348 20668 15379
rect 19944 15320 20668 15348
rect 20717 15351 20775 15357
rect 19944 15308 19950 15320
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 21266 15348 21272 15360
rect 20763 15320 21272 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21376 15348 21404 15379
rect 21450 15376 21456 15428
rect 21508 15416 21514 15428
rect 22373 15419 22431 15425
rect 21508 15388 21553 15416
rect 21508 15376 21514 15388
rect 22373 15385 22385 15419
rect 22419 15416 22431 15419
rect 22554 15416 22560 15428
rect 22419 15388 22560 15416
rect 22419 15385 22431 15388
rect 22373 15379 22431 15385
rect 22554 15376 22560 15388
rect 22612 15376 22618 15428
rect 22922 15416 22928 15428
rect 22883 15388 22928 15416
rect 22922 15376 22928 15388
rect 22980 15376 22986 15428
rect 23014 15376 23020 15428
rect 23072 15416 23078 15428
rect 23072 15388 23117 15416
rect 23072 15376 23078 15388
rect 23198 15376 23204 15428
rect 23256 15416 23262 15428
rect 25130 15416 25136 15428
rect 23256 15388 25136 15416
rect 23256 15376 23262 15388
rect 25130 15376 25136 15388
rect 25188 15376 25194 15428
rect 25409 15419 25467 15425
rect 25409 15385 25421 15419
rect 25455 15385 25467 15419
rect 25409 15379 25467 15385
rect 22002 15348 22008 15360
rect 21376 15320 22008 15348
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22186 15308 22192 15360
rect 22244 15348 22250 15360
rect 24673 15351 24731 15357
rect 24673 15348 24685 15351
rect 22244 15320 24685 15348
rect 22244 15308 22250 15320
rect 24673 15317 24685 15320
rect 24719 15317 24731 15351
rect 25424 15348 25452 15379
rect 26234 15376 26240 15428
rect 26292 15416 26298 15428
rect 26292 15388 26556 15416
rect 26292 15376 26298 15388
rect 26418 15348 26424 15360
rect 25424 15320 26424 15348
rect 24673 15311 24731 15317
rect 26418 15308 26424 15320
rect 26476 15308 26482 15360
rect 26528 15348 26556 15388
rect 26602 15376 26608 15428
rect 26660 15416 26666 15428
rect 27080 15416 27108 15447
rect 29270 15444 29276 15496
rect 29328 15484 29334 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29328 15456 29745 15484
rect 29328 15444 29334 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 29822 15444 29828 15496
rect 29880 15484 29886 15496
rect 30377 15487 30435 15493
rect 30377 15484 30389 15487
rect 29880 15456 30389 15484
rect 29880 15444 29886 15456
rect 30377 15453 30389 15456
rect 30423 15453 30435 15487
rect 30377 15447 30435 15453
rect 31021 15487 31079 15493
rect 31021 15453 31033 15487
rect 31067 15484 31079 15487
rect 35866 15484 35894 15524
rect 37734 15512 37740 15524
rect 37792 15512 37798 15564
rect 31067 15456 35894 15484
rect 31067 15453 31079 15456
rect 31021 15447 31079 15453
rect 37366 15444 37372 15496
rect 37424 15484 37430 15496
rect 38013 15487 38071 15493
rect 38013 15484 38025 15487
rect 37424 15456 38025 15484
rect 37424 15444 37430 15456
rect 38013 15453 38025 15456
rect 38059 15453 38071 15487
rect 38013 15447 38071 15453
rect 28166 15416 28172 15428
rect 26660 15388 27108 15416
rect 27586 15388 28172 15416
rect 26660 15376 26666 15388
rect 27586 15348 27614 15388
rect 28166 15376 28172 15388
rect 28224 15376 28230 15428
rect 28442 15376 28448 15428
rect 28500 15416 28506 15428
rect 28500 15388 28545 15416
rect 28500 15376 28506 15388
rect 28810 15376 28816 15428
rect 28868 15416 28874 15428
rect 31113 15419 31171 15425
rect 31113 15416 31125 15419
rect 28868 15388 31125 15416
rect 28868 15376 28874 15388
rect 31113 15385 31125 15388
rect 31159 15385 31171 15419
rect 31113 15379 31171 15385
rect 26528 15320 27614 15348
rect 27982 15308 27988 15360
rect 28040 15348 28046 15360
rect 29825 15351 29883 15357
rect 29825 15348 29837 15351
rect 28040 15320 29837 15348
rect 28040 15308 28046 15320
rect 29825 15317 29837 15320
rect 29871 15317 29883 15351
rect 29825 15311 29883 15317
rect 30469 15351 30527 15357
rect 30469 15317 30481 15351
rect 30515 15348 30527 15351
rect 30558 15348 30564 15360
rect 30515 15320 30564 15348
rect 30515 15317 30527 15320
rect 30469 15311 30527 15317
rect 30558 15308 30564 15320
rect 30616 15308 30622 15360
rect 38194 15348 38200 15360
rect 38155 15320 38200 15348
rect 38194 15308 38200 15320
rect 38252 15308 38258 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 7834 15144 7840 15156
rect 5408 15116 6500 15144
rect 5408 15104 5414 15116
rect 6472 15088 6500 15116
rect 7668 15116 7840 15144
rect 658 15036 664 15088
rect 716 15076 722 15088
rect 1857 15079 1915 15085
rect 1857 15076 1869 15079
rect 716 15048 1869 15076
rect 716 15036 722 15048
rect 1857 15045 1869 15048
rect 1903 15076 1915 15079
rect 2130 15076 2136 15088
rect 1903 15048 2136 15076
rect 1903 15045 1915 15048
rect 1857 15039 1915 15045
rect 2130 15036 2136 15048
rect 2188 15036 2194 15088
rect 3694 15076 3700 15088
rect 3082 15048 3700 15076
rect 3694 15036 3700 15048
rect 3752 15036 3758 15088
rect 5810 15076 5816 15088
rect 5723 15048 5816 15076
rect 5810 15036 5816 15048
rect 5868 15076 5874 15088
rect 6362 15076 6368 15088
rect 5868 15048 6368 15076
rect 5868 15036 5874 15048
rect 6362 15036 6368 15048
rect 6420 15036 6426 15088
rect 6454 15036 6460 15088
rect 6512 15076 6518 15088
rect 7668 15085 7696 15116
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 11054 15144 11060 15156
rect 9876 15116 11060 15144
rect 7653 15079 7711 15085
rect 6512 15048 7420 15076
rect 6512 15036 6518 15048
rect 1578 15008 1584 15020
rect 1539 14980 1584 15008
rect 1578 14968 1584 14980
rect 1636 14968 1642 15020
rect 4246 15008 4252 15020
rect 4207 14980 4252 15008
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 7392 15017 7420 15048
rect 7653 15045 7665 15079
rect 7699 15045 7711 15079
rect 9490 15076 9496 15088
rect 8878 15048 9496 15076
rect 7653 15039 7711 15045
rect 9490 15036 9496 15048
rect 9548 15036 9554 15088
rect 7377 15011 7435 15017
rect 6549 15001 6607 15007
rect 6549 14967 6561 15001
rect 6595 14998 6607 15001
rect 6656 14998 7328 15008
rect 6595 14980 7328 14998
rect 6595 14970 6684 14980
rect 6595 14967 6607 14970
rect 6549 14961 6607 14967
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 4525 14943 4583 14949
rect 3651 14912 4384 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 3694 14764 3700 14816
rect 3752 14804 3758 14816
rect 3881 14807 3939 14813
rect 3881 14804 3893 14807
rect 3752 14776 3893 14804
rect 3752 14764 3758 14776
rect 3881 14773 3893 14776
rect 3927 14773 3939 14807
rect 4356 14804 4384 14912
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 5074 14940 5080 14952
rect 4571 14912 5080 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 7300 14940 7328 14980
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 15008 9459 15011
rect 9876 15008 9904 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 15746 15144 15752 15156
rect 11164 15116 15752 15144
rect 11164 15085 11192 15116
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 17034 15144 17040 15156
rect 16448 15116 17040 15144
rect 16448 15104 16454 15116
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 17129 15147 17187 15153
rect 17129 15113 17141 15147
rect 17175 15144 17187 15147
rect 17678 15144 17684 15156
rect 17175 15116 17684 15144
rect 17175 15113 17187 15116
rect 17129 15107 17187 15113
rect 17678 15104 17684 15116
rect 17736 15104 17742 15156
rect 18138 15144 18144 15156
rect 17777 15116 18144 15144
rect 10229 15079 10287 15085
rect 10229 15045 10241 15079
rect 10275 15076 10287 15079
rect 11149 15079 11207 15085
rect 10275 15048 11100 15076
rect 10275 15045 10287 15048
rect 10229 15039 10287 15045
rect 9447 14980 9904 15008
rect 11072 15008 11100 15048
rect 11149 15045 11161 15079
rect 11195 15045 11207 15079
rect 11882 15076 11888 15088
rect 11149 15039 11207 15045
rect 11440 15048 11888 15076
rect 11440 15008 11468 15048
rect 11882 15036 11888 15048
rect 11940 15036 11946 15088
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 12066 15076 12072 15088
rect 12023 15048 12072 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 12434 15036 12440 15088
rect 12492 15036 12498 15088
rect 13725 15079 13783 15085
rect 13725 15045 13737 15079
rect 13771 15076 13783 15079
rect 15102 15076 15108 15088
rect 13771 15048 15108 15076
rect 13771 15045 13783 15048
rect 13725 15039 13783 15045
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 15381 15079 15439 15085
rect 15381 15045 15393 15079
rect 15427 15076 15439 15079
rect 17494 15076 17500 15088
rect 15427 15048 17500 15076
rect 15427 15045 15439 15048
rect 15381 15039 15439 15045
rect 17494 15036 17500 15048
rect 17552 15036 17558 15088
rect 17777 15076 17805 15116
rect 18138 15104 18144 15116
rect 18196 15144 18202 15156
rect 19150 15144 19156 15156
rect 18196 15116 19156 15144
rect 18196 15104 18202 15116
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 25225 15147 25283 15153
rect 25225 15144 25237 15147
rect 19536 15116 25237 15144
rect 17604 15048 17805 15076
rect 17865 15079 17923 15085
rect 11072 14980 11468 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11572 14980 11713 15008
rect 11572 14968 11578 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13964 14980 14197 15008
rect 13964 14968 13970 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 16666 14968 16672 15020
rect 16724 15008 16730 15020
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 16724 14980 17049 15008
rect 16724 14968 16730 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 17604 15008 17632 15048
rect 17865 15045 17877 15079
rect 17911 15076 17923 15079
rect 18966 15076 18972 15088
rect 17911 15048 18972 15076
rect 17911 15045 17923 15048
rect 17865 15039 17923 15045
rect 18966 15036 18972 15048
rect 19024 15036 19030 15088
rect 19426 15076 19432 15088
rect 19168 15048 19432 15076
rect 19168 15020 19196 15048
rect 19426 15036 19432 15048
rect 19484 15036 19490 15088
rect 19536 15085 19564 15116
rect 25225 15113 25237 15116
rect 25271 15113 25283 15147
rect 26602 15144 26608 15156
rect 25225 15107 25283 15113
rect 25332 15116 26608 15144
rect 19521 15079 19579 15085
rect 19521 15045 19533 15079
rect 19567 15045 19579 15079
rect 19521 15039 19579 15045
rect 19610 15036 19616 15088
rect 19668 15076 19674 15088
rect 20530 15076 20536 15088
rect 19668 15048 20536 15076
rect 19668 15036 19674 15048
rect 20530 15036 20536 15048
rect 20588 15036 20594 15088
rect 20806 15076 20812 15088
rect 20767 15048 20812 15076
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 20898 15036 20904 15088
rect 20956 15076 20962 15088
rect 21910 15076 21916 15088
rect 20956 15048 21916 15076
rect 20956 15036 20962 15048
rect 21910 15036 21916 15048
rect 21968 15036 21974 15088
rect 22186 15076 22192 15088
rect 22147 15048 22192 15076
rect 22186 15036 22192 15048
rect 22244 15036 22250 15088
rect 23106 15076 23112 15088
rect 23067 15048 23112 15076
rect 23106 15036 23112 15048
rect 23164 15036 23170 15088
rect 23290 15036 23296 15088
rect 23348 15076 23354 15088
rect 23661 15079 23719 15085
rect 23661 15076 23673 15079
rect 23348 15048 23673 15076
rect 23348 15036 23354 15048
rect 23661 15045 23673 15048
rect 23707 15045 23719 15079
rect 23661 15039 23719 15045
rect 23753 15079 23811 15085
rect 23753 15045 23765 15079
rect 23799 15076 23811 15079
rect 24946 15076 24952 15088
rect 23799 15048 24952 15076
rect 23799 15045 23811 15048
rect 23753 15039 23811 15045
rect 24946 15036 24952 15048
rect 25004 15036 25010 15088
rect 25332 15076 25360 15116
rect 26602 15104 26608 15116
rect 26660 15104 26666 15156
rect 27522 15104 27528 15156
rect 27580 15144 27586 15156
rect 27801 15147 27859 15153
rect 27801 15144 27813 15147
rect 27580 15116 27813 15144
rect 27580 15104 27586 15116
rect 27801 15113 27813 15116
rect 27847 15113 27859 15147
rect 29917 15147 29975 15153
rect 29917 15144 29929 15147
rect 27801 15107 27859 15113
rect 27908 15116 29929 15144
rect 25148 15048 25360 15076
rect 19058 15008 19064 15020
rect 17184 14980 17632 15008
rect 18616 14980 19064 15008
rect 17184 14968 17190 14980
rect 9858 14940 9864 14952
rect 7300 14912 9864 14940
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 10137 14943 10195 14949
rect 10137 14909 10149 14943
rect 10183 14909 10195 14943
rect 10137 14903 10195 14909
rect 6914 14872 6920 14884
rect 5552 14844 6920 14872
rect 5552 14804 5580 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 4356 14776 5580 14804
rect 3881 14767 3939 14773
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 5997 14807 6055 14813
rect 5997 14804 6009 14807
rect 5776 14776 6009 14804
rect 5776 14764 5782 14776
rect 5997 14773 6009 14776
rect 6043 14804 6055 14807
rect 6178 14804 6184 14816
rect 6043 14776 6184 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 6641 14807 6699 14813
rect 6641 14773 6653 14807
rect 6687 14804 6699 14807
rect 9950 14804 9956 14816
rect 6687 14776 9956 14804
rect 6687 14773 6699 14776
rect 6641 14767 6699 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10152 14804 10180 14903
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 13446 14940 13452 14952
rect 10652 14912 13452 14940
rect 10652 14900 10658 14912
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 13538 14900 13544 14952
rect 13596 14940 13602 14952
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 13596 14912 14381 14940
rect 13596 14900 13602 14912
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 15378 14940 15384 14952
rect 15335 14912 15384 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 15378 14900 15384 14912
rect 15436 14900 15442 14952
rect 15562 14940 15568 14952
rect 15523 14912 15568 14940
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 17310 14940 17316 14952
rect 16356 14912 17316 14940
rect 16356 14900 16362 14912
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 17773 14943 17831 14949
rect 17773 14909 17785 14943
rect 17819 14940 17831 14943
rect 17862 14940 17868 14952
rect 17819 14912 17868 14940
rect 17819 14909 17831 14912
rect 17773 14903 17831 14909
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 18046 14940 18052 14952
rect 17959 14912 18052 14940
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 18616 14940 18644 14980
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 21361 15011 21419 15017
rect 20128 14980 20577 15008
rect 20128 14968 20134 14980
rect 18156 14912 18644 14940
rect 10502 14832 10508 14884
rect 10560 14872 10566 14884
rect 11146 14872 11152 14884
rect 10560 14844 11152 14872
rect 10560 14832 10566 14844
rect 11146 14832 11152 14844
rect 11204 14872 11210 14884
rect 11606 14872 11612 14884
rect 11204 14844 11612 14872
rect 11204 14832 11210 14844
rect 11606 14832 11612 14844
rect 11664 14832 11670 14884
rect 15102 14832 15108 14884
rect 15160 14872 15166 14884
rect 18064 14872 18092 14900
rect 15160 14844 18092 14872
rect 15160 14832 15166 14844
rect 18156 14804 18184 14912
rect 18782 14900 18788 14952
rect 18840 14940 18846 14952
rect 19242 14940 19248 14952
rect 18840 14912 19248 14940
rect 18840 14900 18846 14912
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19429 14943 19487 14949
rect 19429 14909 19441 14943
rect 19475 14940 19487 14943
rect 19475 14912 19840 14940
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 18690 14872 18696 14884
rect 18380 14844 18696 14872
rect 18380 14832 18386 14844
rect 18690 14832 18696 14844
rect 18748 14872 18754 14884
rect 19702 14872 19708 14884
rect 18748 14844 19708 14872
rect 18748 14832 18754 14844
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 19812 14872 19840 14912
rect 19886 14900 19892 14952
rect 19944 14940 19950 14952
rect 20346 14940 20352 14952
rect 19944 14912 20352 14940
rect 19944 14900 19950 14912
rect 20346 14900 20352 14912
rect 20404 14900 20410 14952
rect 20549 14940 20577 14980
rect 21361 14977 21373 15011
rect 21407 15008 21419 15011
rect 21634 15008 21640 15020
rect 21407 14980 21640 15008
rect 21407 14977 21419 14980
rect 21361 14971 21419 14977
rect 21634 14968 21640 14980
rect 21692 14968 21698 15020
rect 25148 15017 25176 15048
rect 25498 15036 25504 15088
rect 25556 15076 25562 15088
rect 27908 15076 27936 15116
rect 29917 15113 29929 15116
rect 29963 15113 29975 15147
rect 29917 15107 29975 15113
rect 25556 15048 27936 15076
rect 25556 15036 25562 15048
rect 28350 15036 28356 15088
rect 28408 15076 28414 15088
rect 28718 15076 28724 15088
rect 28408 15048 28724 15076
rect 28408 15036 28414 15048
rect 28718 15036 28724 15048
rect 28776 15036 28782 15088
rect 28813 15079 28871 15085
rect 28813 15045 28825 15079
rect 28859 15076 28871 15079
rect 30561 15079 30619 15085
rect 30561 15076 30573 15079
rect 28859 15048 30573 15076
rect 28859 15045 28871 15048
rect 28813 15039 28871 15045
rect 30561 15045 30573 15048
rect 30607 15045 30619 15079
rect 30561 15039 30619 15045
rect 25133 15011 25191 15017
rect 25133 14977 25145 15011
rect 25179 14977 25191 15011
rect 25133 14971 25191 14977
rect 25314 14968 25320 15020
rect 25372 15008 25378 15020
rect 25777 15011 25835 15017
rect 25777 15008 25789 15011
rect 25372 14980 25789 15008
rect 25372 14968 25378 14980
rect 25777 14977 25789 14980
rect 25823 14977 25835 15011
rect 25777 14971 25835 14977
rect 26234 14968 26240 15020
rect 26292 15008 26298 15020
rect 26421 15011 26479 15017
rect 26421 15008 26433 15011
rect 26292 14980 26433 15008
rect 26292 14968 26298 14980
rect 26421 14977 26433 14980
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 15008 27215 15011
rect 27338 15008 27344 15020
rect 27203 14980 27344 15008
rect 27203 14977 27215 14980
rect 27157 14971 27215 14977
rect 27338 14968 27344 14980
rect 27396 14968 27402 15020
rect 29825 15011 29883 15017
rect 29825 14977 29837 15011
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 20717 14943 20775 14949
rect 20549 14912 20677 14940
rect 20530 14872 20536 14884
rect 19812 14844 20536 14872
rect 20530 14832 20536 14844
rect 20588 14832 20594 14884
rect 20649 14872 20677 14912
rect 20717 14909 20729 14943
rect 20763 14940 20775 14943
rect 21818 14940 21824 14952
rect 20763 14912 21824 14940
rect 20763 14909 20775 14912
rect 20717 14903 20775 14909
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 22097 14943 22155 14949
rect 22097 14909 22109 14943
rect 22143 14940 22155 14943
rect 22370 14940 22376 14952
rect 22143 14912 22376 14940
rect 22143 14909 22155 14912
rect 22097 14903 22155 14909
rect 22370 14900 22376 14912
rect 22428 14940 22434 14952
rect 24302 14940 24308 14952
rect 22428 14912 24308 14940
rect 22428 14900 22434 14912
rect 24302 14900 24308 14912
rect 24360 14900 24366 14952
rect 24578 14940 24584 14952
rect 24539 14912 24584 14940
rect 24578 14900 24584 14912
rect 24636 14940 24642 14952
rect 26142 14940 26148 14952
rect 24636 14912 26148 14940
rect 24636 14900 24642 14912
rect 26142 14900 26148 14912
rect 26200 14900 26206 14952
rect 26602 14900 26608 14952
rect 26660 14940 26666 14952
rect 27706 14940 27712 14952
rect 26660 14912 27712 14940
rect 26660 14900 26666 14912
rect 27706 14900 27712 14912
rect 27764 14900 27770 14952
rect 29178 14940 29184 14952
rect 29139 14912 29184 14940
rect 29178 14900 29184 14912
rect 29236 14900 29242 14952
rect 27249 14875 27307 14881
rect 27249 14872 27261 14875
rect 20649 14844 27261 14872
rect 27249 14841 27261 14844
rect 27295 14841 27307 14875
rect 27249 14835 27307 14841
rect 27338 14832 27344 14884
rect 27396 14872 27402 14884
rect 29840 14872 29868 14971
rect 30374 14968 30380 15020
rect 30432 15008 30438 15020
rect 30469 15011 30527 15017
rect 30469 15008 30481 15011
rect 30432 14980 30481 15008
rect 30432 14968 30438 14980
rect 30469 14977 30481 14980
rect 30515 14977 30527 15011
rect 31110 15008 31116 15020
rect 31071 14980 31116 15008
rect 30469 14971 30527 14977
rect 31110 14968 31116 14980
rect 31168 14968 31174 15020
rect 37734 14968 37740 15020
rect 37792 15008 37798 15020
rect 38013 15011 38071 15017
rect 38013 15008 38025 15011
rect 37792 14980 38025 15008
rect 37792 14968 37798 14980
rect 38013 14977 38025 14980
rect 38059 14977 38071 15011
rect 38013 14971 38071 14977
rect 27396 14844 29868 14872
rect 27396 14832 27402 14844
rect 10152 14776 18184 14804
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 23382 14804 23388 14816
rect 19024 14776 23388 14804
rect 19024 14764 19030 14776
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 23566 14764 23572 14816
rect 23624 14804 23630 14816
rect 24486 14804 24492 14816
rect 23624 14776 24492 14804
rect 23624 14764 23630 14776
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 25682 14764 25688 14816
rect 25740 14804 25746 14816
rect 25869 14807 25927 14813
rect 25869 14804 25881 14807
rect 25740 14776 25881 14804
rect 25740 14764 25746 14776
rect 25869 14773 25881 14776
rect 25915 14773 25927 14807
rect 25869 14767 25927 14773
rect 26513 14807 26571 14813
rect 26513 14773 26525 14807
rect 26559 14804 26571 14807
rect 26878 14804 26884 14816
rect 26559 14776 26884 14804
rect 26559 14773 26571 14776
rect 26513 14767 26571 14773
rect 26878 14764 26884 14776
rect 26936 14764 26942 14816
rect 27062 14764 27068 14816
rect 27120 14804 27126 14816
rect 29822 14804 29828 14816
rect 27120 14776 29828 14804
rect 27120 14764 27126 14776
rect 29822 14764 29828 14776
rect 29880 14764 29886 14816
rect 31202 14804 31208 14816
rect 31163 14776 31208 14804
rect 31202 14764 31208 14776
rect 31260 14764 31266 14816
rect 37829 14807 37887 14813
rect 37829 14773 37841 14807
rect 37875 14804 37887 14807
rect 38010 14804 38016 14816
rect 37875 14776 38016 14804
rect 37875 14773 37887 14776
rect 37829 14767 37887 14773
rect 38010 14764 38016 14776
rect 38068 14764 38074 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 10778 14600 10784 14612
rect 7616 14572 10784 14600
rect 7616 14560 7622 14572
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 10952 14603 11010 14609
rect 10952 14569 10964 14603
rect 10998 14600 11010 14603
rect 11422 14600 11428 14612
rect 10998 14572 11428 14600
rect 10998 14569 11010 14572
rect 10952 14563 11010 14569
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 15102 14600 15108 14612
rect 11664 14572 15108 14600
rect 11664 14560 11670 14572
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 18690 14600 18696 14612
rect 15252 14572 18696 14600
rect 15252 14560 15258 14572
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 21542 14600 21548 14612
rect 18840 14572 21548 14600
rect 18840 14560 18846 14572
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 22152 14572 22197 14600
rect 22152 14560 22158 14572
rect 23290 14560 23296 14612
rect 23348 14600 23354 14612
rect 23753 14603 23811 14609
rect 23753 14600 23765 14603
rect 23348 14572 23765 14600
rect 23348 14560 23354 14572
rect 23753 14569 23765 14572
rect 23799 14569 23811 14603
rect 23753 14563 23811 14569
rect 26418 14560 26424 14612
rect 26476 14600 26482 14612
rect 27065 14603 27123 14609
rect 27065 14600 27077 14603
rect 26476 14572 27077 14600
rect 26476 14560 26482 14572
rect 27065 14569 27077 14572
rect 27111 14569 27123 14603
rect 27706 14600 27712 14612
rect 27667 14572 27712 14600
rect 27065 14563 27123 14569
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 37366 14600 37372 14612
rect 37327 14572 37372 14600
rect 37366 14560 37372 14572
rect 37424 14560 37430 14612
rect 5350 14492 5356 14544
rect 5408 14492 5414 14544
rect 7926 14492 7932 14544
rect 7984 14532 7990 14544
rect 10502 14532 10508 14544
rect 7984 14504 10508 14532
rect 7984 14492 7990 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 13998 14532 14004 14544
rect 12728 14504 14004 14532
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 1673 14467 1731 14473
rect 1673 14464 1685 14467
rect 1636 14436 1685 14464
rect 1636 14424 1642 14436
rect 1673 14433 1685 14436
rect 1719 14433 1731 14467
rect 1673 14427 1731 14433
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 3142 14464 3148 14476
rect 1995 14436 3148 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14464 4031 14467
rect 5368 14464 5396 14492
rect 5994 14464 6000 14476
rect 4019 14436 5396 14464
rect 5955 14436 6000 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6546 14464 6552 14476
rect 6507 14436 6552 14464
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 7432 14436 9505 14464
rect 7432 14424 7438 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10594 14464 10600 14476
rect 10008 14436 10600 14464
rect 10008 14424 10014 14436
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 11514 14464 11520 14476
rect 10735 14436 11520 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 12728 14473 12756 14504
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 14274 14492 14280 14544
rect 14332 14532 14338 14544
rect 17402 14532 17408 14544
rect 14332 14504 17408 14532
rect 14332 14492 14338 14504
rect 17402 14492 17408 14504
rect 17460 14492 17466 14544
rect 17494 14492 17500 14544
rect 17552 14532 17558 14544
rect 17552 14504 17908 14532
rect 17552 14492 17558 14504
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14433 12771 14467
rect 12713 14427 12771 14433
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 13044 14436 13369 14464
rect 13044 14424 13050 14436
rect 13357 14433 13369 14436
rect 13403 14464 13415 14467
rect 15102 14464 15108 14476
rect 13403 14436 15108 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 16390 14464 16396 14476
rect 15436 14436 16396 14464
rect 15436 14424 15442 14436
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14464 16543 14467
rect 16574 14464 16580 14476
rect 16531 14436 16580 14464
rect 16531 14433 16543 14436
rect 16485 14427 16543 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 17586 14464 17592 14476
rect 16816 14436 17592 14464
rect 16816 14424 16822 14436
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 17880 14473 17908 14504
rect 17954 14492 17960 14544
rect 18012 14492 18018 14544
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 19886 14532 19892 14544
rect 18104 14504 19892 14532
rect 18104 14492 18110 14504
rect 19886 14492 19892 14504
rect 19944 14492 19950 14544
rect 19978 14492 19984 14544
rect 20036 14532 20042 14544
rect 20438 14532 20444 14544
rect 20036 14504 20444 14532
rect 20036 14492 20042 14504
rect 20438 14492 20444 14504
rect 20496 14492 20502 14544
rect 27614 14532 27620 14544
rect 22572 14504 27620 14532
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 17972 14464 18000 14492
rect 17972 14436 20392 14464
rect 17865 14427 17923 14433
rect 5350 14356 5356 14408
rect 5408 14356 5414 14408
rect 8754 14396 8760 14408
rect 8220 14368 8760 14396
rect 3878 14328 3884 14340
rect 3174 14300 3884 14328
rect 3878 14288 3884 14300
rect 3936 14288 3942 14340
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14297 4307 14331
rect 6822 14328 6828 14340
rect 6783 14300 6828 14328
rect 4249 14291 4307 14297
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3421 14263 3479 14269
rect 3421 14260 3433 14263
rect 2832 14232 3433 14260
rect 2832 14220 2838 14232
rect 3421 14229 3433 14232
rect 3467 14229 3479 14263
rect 4264 14260 4292 14291
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 8110 14328 8116 14340
rect 8050 14300 8116 14328
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 5534 14260 5540 14272
rect 4264 14232 5540 14260
rect 3421 14223 3479 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 8220 14260 8248 14368
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 12860 14368 13185 14396
rect 12860 14356 12866 14368
rect 13173 14365 13185 14368
rect 13219 14396 13231 14399
rect 13906 14396 13912 14408
rect 13219 14368 13912 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 17218 14396 17224 14408
rect 14108 14368 17224 14396
rect 8573 14331 8631 14337
rect 8573 14297 8585 14331
rect 8619 14297 8631 14331
rect 8573 14291 8631 14297
rect 6144 14232 8248 14260
rect 8588 14260 8616 14291
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 10137 14331 10195 14337
rect 9640 14300 9685 14328
rect 9640 14288 9646 14300
rect 10137 14297 10149 14331
rect 10183 14328 10195 14331
rect 11238 14328 11244 14340
rect 10183 14300 11244 14328
rect 10183 14297 10195 14300
rect 10137 14291 10195 14297
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 13630 14328 13636 14340
rect 12190 14300 13636 14328
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 10318 14260 10324 14272
rect 8588 14232 10324 14260
rect 6144 14220 6150 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 14108 14260 14136 14368
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 18892 14396 19104 14406
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 18892 14378 19441 14396
rect 14274 14328 14280 14340
rect 14235 14300 14280 14328
rect 14274 14288 14280 14300
rect 14332 14288 14338 14340
rect 14458 14288 14464 14340
rect 14516 14328 14522 14340
rect 14516 14300 16988 14328
rect 14516 14288 14522 14300
rect 10560 14232 14136 14260
rect 10560 14220 10566 14232
rect 14366 14220 14372 14272
rect 14424 14260 14430 14272
rect 15565 14263 15623 14269
rect 15565 14260 15577 14263
rect 14424 14232 15577 14260
rect 14424 14220 14430 14232
rect 15565 14229 15577 14232
rect 15611 14229 15623 14263
rect 15565 14223 15623 14229
rect 15654 14220 15660 14272
rect 15712 14260 15718 14272
rect 16850 14260 16856 14272
rect 15712 14232 16856 14260
rect 15712 14220 15718 14232
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 16960 14260 16988 14300
rect 17034 14288 17040 14340
rect 17092 14328 17098 14340
rect 17589 14331 17647 14337
rect 17589 14328 17601 14331
rect 17092 14300 17601 14328
rect 17092 14288 17098 14300
rect 17589 14297 17601 14300
rect 17635 14297 17647 14331
rect 17589 14291 17647 14297
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 17736 14300 17781 14328
rect 17736 14288 17742 14300
rect 17494 14260 17500 14272
rect 16960 14232 17500 14260
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 17770 14220 17776 14272
rect 17828 14260 17834 14272
rect 18892 14260 18920 14378
rect 19076 14368 19441 14378
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19444 14328 19472 14359
rect 19444 14300 20300 14328
rect 20272 14272 20300 14300
rect 17828 14232 18920 14260
rect 17828 14220 17834 14232
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19521 14263 19579 14269
rect 19521 14260 19533 14263
rect 19392 14232 19533 14260
rect 19392 14220 19398 14232
rect 19521 14229 19533 14232
rect 19567 14229 19579 14263
rect 19521 14223 19579 14229
rect 20254 14220 20260 14272
rect 20312 14220 20318 14272
rect 20364 14260 20392 14436
rect 20530 14424 20536 14476
rect 20588 14464 20594 14476
rect 20588 14436 21680 14464
rect 20588 14424 20594 14436
rect 21652 14408 21680 14436
rect 21634 14356 21640 14408
rect 21692 14356 21698 14408
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14396 22063 14399
rect 22094 14396 22100 14408
rect 22051 14368 22100 14396
rect 22051 14365 22063 14368
rect 22005 14359 22063 14365
rect 22094 14356 22100 14368
rect 22152 14396 22158 14408
rect 22572 14396 22600 14504
rect 27614 14492 27620 14504
rect 27672 14492 27678 14544
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 24026 14464 24032 14476
rect 22704 14436 24032 14464
rect 22704 14424 22710 14436
rect 24026 14424 24032 14436
rect 24084 14424 24090 14476
rect 24673 14467 24731 14473
rect 24673 14464 24685 14467
rect 24136 14436 24685 14464
rect 22152 14368 22600 14396
rect 22152 14356 22158 14368
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 23658 14396 23664 14408
rect 22796 14368 23152 14396
rect 23619 14368 23664 14396
rect 22796 14356 22802 14368
rect 20634 14331 20692 14337
rect 20634 14297 20646 14331
rect 20680 14328 20692 14331
rect 21542 14328 21548 14340
rect 20680 14300 21220 14328
rect 21455 14300 21548 14328
rect 20680 14297 20692 14300
rect 20634 14291 20692 14297
rect 21192 14272 21220 14300
rect 21542 14288 21548 14300
rect 21600 14328 21606 14340
rect 22278 14328 22284 14340
rect 21600 14300 22284 14328
rect 21600 14288 21606 14300
rect 22278 14288 22284 14300
rect 22336 14288 22342 14340
rect 22370 14288 22376 14340
rect 22428 14328 22434 14340
rect 23017 14331 23075 14337
rect 23017 14328 23029 14331
rect 22428 14300 23029 14328
rect 22428 14288 22434 14300
rect 23017 14297 23029 14300
rect 23063 14297 23075 14331
rect 23124 14328 23152 14368
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 24136 14328 24164 14436
rect 24673 14433 24685 14436
rect 24719 14464 24731 14467
rect 24719 14436 25544 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 25317 14399 25375 14405
rect 25317 14365 25329 14399
rect 25363 14396 25375 14399
rect 25406 14396 25412 14408
rect 25363 14368 25412 14396
rect 25363 14365 25375 14368
rect 25317 14359 25375 14365
rect 23124 14300 24164 14328
rect 24765 14331 24823 14337
rect 23017 14291 23075 14297
rect 24765 14297 24777 14331
rect 24811 14297 24823 14331
rect 24765 14291 24823 14297
rect 21082 14260 21088 14272
rect 20364 14232 21088 14260
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 21174 14220 21180 14272
rect 21232 14220 21238 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22738 14260 22744 14272
rect 21876 14232 22744 14260
rect 21876 14220 21882 14232
rect 22738 14220 22744 14232
rect 22796 14220 22802 14272
rect 22830 14220 22836 14272
rect 22888 14260 22894 14272
rect 23109 14263 23167 14269
rect 23109 14260 23121 14263
rect 22888 14232 23121 14260
rect 22888 14220 22894 14232
rect 23109 14229 23121 14232
rect 23155 14229 23167 14263
rect 23109 14223 23167 14229
rect 23290 14220 23296 14272
rect 23348 14260 23354 14272
rect 24578 14260 24584 14272
rect 23348 14232 24584 14260
rect 23348 14220 23354 14232
rect 24578 14220 24584 14232
rect 24636 14220 24642 14272
rect 24780 14260 24808 14291
rect 24854 14288 24860 14340
rect 24912 14328 24918 14340
rect 25332 14328 25360 14359
rect 25406 14356 25412 14368
rect 25464 14356 25470 14408
rect 24912 14300 25360 14328
rect 25516 14328 25544 14436
rect 25682 14424 25688 14476
rect 25740 14464 25746 14476
rect 28353 14467 28411 14473
rect 28353 14464 28365 14467
rect 25740 14436 28365 14464
rect 25740 14424 25746 14436
rect 28353 14433 28365 14436
rect 28399 14433 28411 14467
rect 28353 14427 28411 14433
rect 29546 14424 29552 14476
rect 29604 14464 29610 14476
rect 30282 14464 30288 14476
rect 29604 14436 30288 14464
rect 29604 14424 29610 14436
rect 30282 14424 30288 14436
rect 30340 14464 30346 14476
rect 31113 14467 31171 14473
rect 31113 14464 31125 14467
rect 30340 14436 31125 14464
rect 30340 14424 30346 14436
rect 31113 14433 31125 14436
rect 31159 14433 31171 14467
rect 31386 14464 31392 14476
rect 31347 14436 31392 14464
rect 31113 14427 31171 14433
rect 31386 14424 31392 14436
rect 31444 14424 31450 14476
rect 26981 14401 27039 14407
rect 26981 14367 26993 14401
rect 27027 14367 27039 14401
rect 26981 14361 27039 14367
rect 25866 14328 25872 14340
rect 25516 14300 25872 14328
rect 24912 14288 24918 14300
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 25961 14331 26019 14337
rect 25961 14297 25973 14331
rect 26007 14297 26019 14331
rect 26510 14328 26516 14340
rect 26471 14300 26516 14328
rect 25961 14291 26019 14297
rect 25682 14260 25688 14272
rect 24780 14232 25688 14260
rect 25682 14220 25688 14232
rect 25740 14220 25746 14272
rect 25976 14260 26004 14291
rect 26510 14288 26516 14300
rect 26568 14288 26574 14340
rect 26602 14288 26608 14340
rect 26660 14328 26666 14340
rect 26988 14328 27016 14361
rect 27154 14356 27160 14408
rect 27212 14356 27218 14408
rect 27614 14356 27620 14408
rect 27672 14396 27678 14408
rect 28261 14399 28319 14405
rect 28261 14396 28273 14399
rect 27672 14368 27715 14396
rect 28092 14368 28273 14396
rect 27672 14356 27678 14368
rect 26660 14300 27016 14328
rect 26660 14288 26666 14300
rect 27172 14260 27200 14356
rect 25976 14232 27200 14260
rect 27706 14220 27712 14272
rect 27764 14260 27770 14272
rect 27890 14260 27896 14272
rect 27764 14232 27896 14260
rect 27764 14220 27770 14232
rect 27890 14220 27896 14232
rect 27948 14220 27954 14272
rect 28092 14260 28120 14368
rect 28261 14365 28273 14368
rect 28307 14365 28319 14399
rect 28261 14359 28319 14365
rect 28442 14356 28448 14408
rect 28500 14396 28506 14408
rect 28905 14399 28963 14405
rect 28905 14396 28917 14399
rect 28500 14368 28917 14396
rect 28500 14356 28506 14368
rect 28905 14365 28917 14368
rect 28951 14365 28963 14399
rect 28905 14359 28963 14365
rect 29914 14356 29920 14408
rect 29972 14396 29978 14408
rect 30377 14399 30435 14405
rect 30377 14396 30389 14399
rect 29972 14368 30389 14396
rect 29972 14356 29978 14368
rect 30377 14365 30389 14368
rect 30423 14365 30435 14399
rect 30377 14359 30435 14365
rect 37182 14356 37188 14408
rect 37240 14396 37246 14408
rect 37553 14399 37611 14405
rect 37553 14396 37565 14399
rect 37240 14368 37565 14396
rect 37240 14356 37246 14368
rect 37553 14365 37565 14368
rect 37599 14365 37611 14399
rect 37553 14359 37611 14365
rect 37918 14356 37924 14408
rect 37976 14396 37982 14408
rect 38013 14399 38071 14405
rect 38013 14396 38025 14399
rect 37976 14368 38025 14396
rect 37976 14356 37982 14368
rect 38013 14365 38025 14368
rect 38059 14365 38071 14399
rect 38013 14359 38071 14365
rect 28166 14288 28172 14340
rect 28224 14328 28230 14340
rect 28997 14331 29055 14337
rect 28997 14328 29009 14331
rect 28224 14300 29009 14328
rect 28224 14288 28230 14300
rect 28997 14297 29009 14300
rect 29043 14297 29055 14331
rect 31110 14328 31116 14340
rect 28997 14291 29055 14297
rect 29564 14300 31116 14328
rect 28350 14260 28356 14272
rect 28092 14232 28356 14260
rect 28350 14220 28356 14232
rect 28408 14220 28414 14272
rect 28902 14220 28908 14272
rect 28960 14260 28966 14272
rect 29564 14260 29592 14300
rect 31110 14288 31116 14300
rect 31168 14288 31174 14340
rect 31202 14288 31208 14340
rect 31260 14328 31266 14340
rect 31260 14300 31305 14328
rect 31260 14288 31266 14300
rect 29730 14260 29736 14272
rect 28960 14232 29592 14260
rect 29691 14232 29736 14260
rect 28960 14220 28966 14232
rect 29730 14220 29736 14232
rect 29788 14220 29794 14272
rect 30466 14260 30472 14272
rect 30427 14232 30472 14260
rect 30466 14220 30472 14232
rect 30524 14220 30530 14272
rect 38194 14260 38200 14272
rect 38155 14232 38200 14260
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9858 14056 9864 14068
rect 5644 14028 9864 14056
rect 4522 13988 4528 14000
rect 4483 13960 4528 13988
rect 4522 13948 4528 13960
rect 4580 13948 4586 14000
rect 5445 13991 5503 13997
rect 5445 13957 5457 13991
rect 5491 13988 5503 13991
rect 5644 13988 5672 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 20070 14056 20076 14068
rect 11164 14028 16620 14056
rect 7926 13988 7932 14000
rect 5491 13960 5672 13988
rect 6196 13960 7932 13988
rect 5491 13957 5503 13960
rect 5445 13951 5503 13957
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 1854 13920 1860 13932
rect 1627 13892 1860 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 3878 13880 3884 13932
rect 3936 13880 3942 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6086 13920 6092 13932
rect 6043 13892 6092 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 2498 13852 2504 13864
rect 2459 13824 2504 13852
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13852 2835 13855
rect 4062 13852 4068 13864
rect 2823 13824 4068 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 4062 13812 4068 13824
rect 4120 13852 4126 13864
rect 4706 13852 4712 13864
rect 4120 13824 4712 13852
rect 4120 13812 4126 13824
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 6196 13852 6224 13960
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 10502 13988 10508 14000
rect 8878 13960 10508 13988
rect 10502 13948 10508 13960
rect 10560 13948 10566 14000
rect 10594 13948 10600 14000
rect 10652 13988 10658 14000
rect 11164 13997 11192 14028
rect 11149 13991 11207 13997
rect 10652 13960 10697 13988
rect 10652 13948 10658 13960
rect 11149 13957 11161 13991
rect 11195 13957 11207 13991
rect 11974 13988 11980 14000
rect 11935 13960 11980 13988
rect 11149 13951 11207 13957
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 14461 13991 14519 13997
rect 14461 13988 14473 13991
rect 13280 13960 14473 13988
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6328 13892 6561 13920
rect 6328 13880 6334 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 5399 13824 6224 13852
rect 6564 13824 7389 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 6564 13796 6592 13824
rect 7377 13821 7389 13824
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13852 7711 13855
rect 8386 13852 8392 13864
rect 7699 13824 8392 13852
rect 7699 13821 7711 13824
rect 7653 13815 7711 13821
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 9306 13812 9312 13864
rect 9364 13852 9370 13864
rect 9401 13855 9459 13861
rect 9401 13852 9413 13855
rect 9364 13824 9413 13852
rect 9364 13812 9370 13824
rect 9401 13821 9413 13824
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10505 13855 10563 13861
rect 10505 13852 10517 13855
rect 10100 13824 10517 13852
rect 10100 13812 10106 13824
rect 10505 13821 10517 13824
rect 10551 13821 10563 13855
rect 11698 13852 11704 13864
rect 10505 13815 10563 13821
rect 10612 13824 11560 13852
rect 11659 13824 11704 13852
rect 6546 13744 6552 13796
rect 6604 13744 6610 13796
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10612 13784 10640 13824
rect 10376 13756 10640 13784
rect 11532 13784 11560 13824
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 13096 13852 13124 13906
rect 13280 13852 13308 13960
rect 14461 13957 14473 13960
rect 14507 13957 14519 13991
rect 14461 13951 14519 13957
rect 15010 13948 15016 14000
rect 15068 13988 15074 14000
rect 16298 13988 16304 14000
rect 15068 13960 16304 13988
rect 15068 13948 15074 13960
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 15838 13920 15844 13932
rect 15799 13892 15844 13920
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 11808 13824 13124 13852
rect 13188 13824 13308 13852
rect 11808 13784 11836 13824
rect 11532 13756 11836 13784
rect 10376 13744 10382 13756
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 6733 13719 6791 13725
rect 6733 13716 6745 13719
rect 3844 13688 6745 13716
rect 3844 13676 3850 13688
rect 6733 13685 6745 13688
rect 6779 13685 6791 13719
rect 6733 13679 6791 13685
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 11606 13716 11612 13728
rect 6972 13688 11612 13716
rect 6972 13676 6978 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 13188 13716 13216 13824
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13725 13855 13783 13861
rect 13725 13852 13737 13855
rect 13412 13824 13737 13852
rect 13412 13812 13418 13824
rect 13725 13821 13737 13824
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14642 13852 14648 13864
rect 14415 13824 14648 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15194 13852 15200 13864
rect 15155 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13821 16175 13855
rect 16592 13852 16620 14028
rect 17505 14028 20076 14056
rect 16942 13988 16948 14000
rect 16903 13960 16948 13988
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 17505 13988 17533 14028
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 21174 14056 21180 14068
rect 21135 14028 21180 14056
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 22278 14056 22284 14068
rect 21928 14028 22284 14056
rect 21928 14000 21956 14028
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 22554 14016 22560 14068
rect 22612 14056 22618 14068
rect 23290 14056 23296 14068
rect 22612 14028 23296 14056
rect 22612 14016 22618 14028
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 26513 14059 26571 14065
rect 26513 14056 26525 14059
rect 23400 14028 26525 14056
rect 17083 13960 17533 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 18322 13988 18328 14000
rect 17920 13960 18328 13988
rect 17920 13948 17926 13960
rect 18322 13948 18328 13960
rect 18380 13948 18386 14000
rect 18506 13948 18512 14000
rect 18564 13988 18570 14000
rect 19058 13988 19064 14000
rect 18564 13960 19064 13988
rect 18564 13948 18570 13960
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 19150 13948 19156 14000
rect 19208 13988 19214 14000
rect 19521 13991 19579 13997
rect 19521 13988 19533 13991
rect 19208 13960 19533 13988
rect 19208 13948 19214 13960
rect 19521 13957 19533 13960
rect 19567 13957 19579 13991
rect 19521 13951 19579 13957
rect 19613 13991 19671 13997
rect 19613 13957 19625 13991
rect 19659 13988 19671 13991
rect 19886 13988 19892 14000
rect 19659 13960 19892 13988
rect 19659 13957 19671 13960
rect 19613 13951 19671 13957
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20533 13991 20591 13997
rect 20533 13957 20545 13991
rect 20579 13988 20591 13991
rect 20622 13988 20628 14000
rect 20579 13960 20628 13988
rect 20579 13957 20591 13960
rect 20533 13951 20591 13957
rect 20622 13948 20628 13960
rect 20680 13988 20686 14000
rect 21542 13988 21548 14000
rect 20680 13960 21548 13988
rect 20680 13948 20686 13960
rect 21542 13948 21548 13960
rect 21600 13948 21606 14000
rect 21910 13948 21916 14000
rect 21968 13948 21974 14000
rect 22186 13988 22192 14000
rect 22147 13960 22192 13988
rect 22186 13948 22192 13960
rect 22244 13948 22250 14000
rect 23400 13997 23428 14028
rect 26513 14025 26525 14028
rect 26559 14025 26571 14059
rect 26513 14019 26571 14025
rect 26602 14016 26608 14068
rect 26660 14056 26666 14068
rect 28902 14056 28908 14068
rect 26660 14028 28908 14056
rect 26660 14016 26666 14028
rect 23385 13991 23443 13997
rect 23385 13957 23397 13991
rect 23431 13957 23443 13991
rect 23385 13951 23443 13957
rect 25041 13991 25099 13997
rect 25041 13957 25053 13991
rect 25087 13988 25099 13991
rect 27893 13991 27951 13997
rect 27893 13988 27905 13991
rect 25087 13960 27905 13988
rect 25087 13957 25099 13960
rect 25041 13951 25099 13957
rect 27893 13957 27905 13960
rect 27939 13957 27951 13991
rect 27893 13951 27951 13957
rect 18046 13920 18052 13932
rect 18007 13892 18052 13920
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 18196 13892 18241 13920
rect 18196 13880 18202 13892
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 18472 13892 18705 13920
rect 18472 13880 18478 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20990 13920 20996 13932
rect 20496 13892 20996 13920
rect 20496 13880 20502 13892
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13920 21143 13923
rect 21818 13920 21824 13932
rect 21131 13892 21824 13920
rect 21131 13889 21143 13892
rect 21085 13883 21143 13889
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 22738 13880 22744 13932
rect 22796 13920 22802 13932
rect 23106 13920 23112 13932
rect 22796 13892 23112 13920
rect 22796 13880 22802 13892
rect 23106 13880 23112 13892
rect 23164 13880 23170 13932
rect 24578 13920 24584 13932
rect 23952 13892 24584 13920
rect 17310 13852 17316 13864
rect 16592 13824 17316 13852
rect 16117 13815 16175 13821
rect 11848 13688 13216 13716
rect 16132 13716 16160 13815
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 17644 13840 18184 13852
rect 18237 13840 18797 13852
rect 17644 13824 18797 13840
rect 17644 13812 17650 13824
rect 18156 13812 18265 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 20898 13852 20904 13864
rect 19208 13824 20904 13852
rect 19208 13812 19214 13824
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 22094 13852 22100 13864
rect 22055 13824 22100 13852
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 22462 13852 22468 13864
rect 22423 13824 22468 13852
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 23293 13855 23351 13861
rect 23293 13852 23305 13855
rect 22756 13824 23305 13852
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 17497 13787 17555 13793
rect 17497 13784 17509 13787
rect 16264 13756 17509 13784
rect 16264 13744 16270 13756
rect 17497 13753 17509 13756
rect 17543 13784 17555 13787
rect 18046 13784 18052 13796
rect 17543 13756 18052 13784
rect 17543 13753 17555 13756
rect 17497 13747 17555 13753
rect 18046 13744 18052 13756
rect 18104 13744 18110 13796
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 19426 13784 19432 13796
rect 18472 13756 19432 13784
rect 18472 13744 18478 13756
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 19518 13744 19524 13796
rect 19576 13784 19582 13796
rect 19576 13756 22048 13784
rect 19576 13744 19582 13756
rect 17770 13716 17776 13728
rect 16132 13688 17776 13716
rect 11848 13676 11854 13688
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 17862 13676 17868 13728
rect 17920 13716 17926 13728
rect 18322 13716 18328 13728
rect 17920 13688 18328 13716
rect 17920 13676 17926 13688
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 18506 13676 18512 13728
rect 18564 13716 18570 13728
rect 21910 13716 21916 13728
rect 18564 13688 21916 13716
rect 18564 13676 18570 13688
rect 21910 13676 21916 13688
rect 21968 13676 21974 13728
rect 22020 13716 22048 13756
rect 22756 13716 22784 13824
rect 23293 13821 23305 13824
rect 23339 13852 23351 13855
rect 23952 13852 23980 13892
rect 24578 13880 24584 13892
rect 24636 13880 24642 13932
rect 26418 13920 26424 13932
rect 26379 13892 26424 13920
rect 26418 13880 26424 13892
rect 26476 13880 26482 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 27706 13920 27712 13932
rect 27203 13892 27712 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 27706 13880 27712 13892
rect 27764 13880 27770 13932
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13920 27859 13923
rect 28000 13920 28028 14028
rect 28902 14016 28908 14028
rect 28960 14016 28966 14068
rect 29730 14056 29736 14068
rect 29012 14028 29736 14056
rect 29012 13997 29040 14028
rect 29730 14016 29736 14028
rect 29788 14016 29794 14068
rect 30282 14016 30288 14068
rect 30340 14056 30346 14068
rect 30745 14059 30803 14065
rect 30745 14056 30757 14059
rect 30340 14028 30757 14056
rect 30340 14016 30346 14028
rect 30745 14025 30757 14028
rect 30791 14025 30803 14059
rect 30745 14019 30803 14025
rect 37182 14016 37188 14068
rect 37240 14056 37246 14068
rect 38105 14059 38163 14065
rect 38105 14056 38117 14059
rect 37240 14028 38117 14056
rect 37240 14016 37246 14028
rect 38105 14025 38117 14028
rect 38151 14025 38163 14059
rect 38105 14019 38163 14025
rect 28997 13991 29055 13997
rect 28997 13957 29009 13991
rect 29043 13957 29055 13991
rect 28997 13951 29055 13957
rect 29089 13991 29147 13997
rect 29089 13957 29101 13991
rect 29135 13988 29147 13991
rect 30466 13988 30472 14000
rect 29135 13960 30472 13988
rect 29135 13957 29147 13960
rect 29089 13951 29147 13957
rect 30466 13948 30472 13960
rect 30524 13948 30530 14000
rect 27847 13892 28028 13920
rect 30653 13923 30711 13929
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 30653 13889 30665 13923
rect 30699 13920 30711 13923
rect 37734 13920 37740 13932
rect 30699 13892 37740 13920
rect 30699 13889 30711 13892
rect 30653 13883 30711 13889
rect 37734 13880 37740 13892
rect 37792 13880 37798 13932
rect 38286 13920 38292 13932
rect 38247 13892 38292 13920
rect 38286 13880 38292 13892
rect 38344 13880 38350 13932
rect 23339 13824 23980 13852
rect 23339 13821 23351 13824
rect 23293 13815 23351 13821
rect 24302 13812 24308 13864
rect 24360 13852 24366 13864
rect 24949 13855 25007 13861
rect 24949 13852 24961 13855
rect 24360 13824 24961 13852
rect 24360 13812 24366 13824
rect 24949 13821 24961 13824
rect 24995 13852 25007 13855
rect 25406 13852 25412 13864
rect 24995 13824 25412 13852
rect 24995 13821 25007 13824
rect 24949 13815 25007 13821
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25866 13852 25872 13864
rect 25827 13824 25872 13852
rect 25866 13812 25872 13824
rect 25924 13852 25930 13864
rect 27062 13852 27068 13864
rect 25924 13824 27068 13852
rect 25924 13812 25930 13824
rect 27062 13812 27068 13824
rect 27120 13812 27126 13864
rect 29362 13852 29368 13864
rect 29323 13824 29368 13852
rect 29362 13812 29368 13824
rect 29420 13812 29426 13864
rect 23106 13744 23112 13796
rect 23164 13784 23170 13796
rect 23845 13787 23903 13793
rect 23845 13784 23857 13787
rect 23164 13756 23857 13784
rect 23164 13744 23170 13756
rect 23845 13753 23857 13756
rect 23891 13784 23903 13787
rect 24854 13784 24860 13796
rect 23891 13756 24860 13784
rect 23891 13753 23903 13756
rect 23845 13747 23903 13753
rect 24854 13744 24860 13756
rect 24912 13744 24918 13796
rect 30558 13784 30564 13796
rect 24964 13756 30564 13784
rect 22020 13688 22784 13716
rect 23934 13676 23940 13728
rect 23992 13716 23998 13728
rect 24964 13716 24992 13756
rect 30558 13744 30564 13756
rect 30616 13744 30622 13796
rect 27246 13716 27252 13728
rect 23992 13688 24992 13716
rect 27207 13688 27252 13716
rect 23992 13676 23998 13688
rect 27246 13676 27252 13688
rect 27304 13676 27310 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4798 13512 4804 13524
rect 3467 13484 4804 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 11146 13512 11152 13524
rect 5868 13484 11152 13512
rect 5868 13472 5874 13484
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 20806 13512 20812 13524
rect 11256 13484 20812 13512
rect 10594 13404 10600 13456
rect 10652 13444 10658 13456
rect 11256 13444 11284 13484
rect 20806 13472 20812 13484
rect 20864 13472 20870 13524
rect 20898 13472 20904 13524
rect 20956 13512 20962 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 20956 13484 21005 13512
rect 20956 13472 20962 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 21450 13472 21456 13524
rect 21508 13512 21514 13524
rect 23201 13515 23259 13521
rect 23201 13512 23213 13515
rect 21508 13484 23213 13512
rect 21508 13472 21514 13484
rect 23201 13481 23213 13484
rect 23247 13481 23259 13515
rect 23201 13475 23259 13481
rect 23382 13472 23388 13524
rect 23440 13512 23446 13524
rect 23845 13515 23903 13521
rect 23845 13512 23857 13515
rect 23440 13484 23857 13512
rect 23440 13472 23446 13484
rect 23845 13481 23857 13484
rect 23891 13481 23903 13515
rect 29362 13512 29368 13524
rect 23845 13475 23903 13481
rect 26436 13484 29368 13512
rect 10652 13416 11284 13444
rect 10652 13404 10658 13416
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 20530 13444 20536 13456
rect 13320 13416 20536 13444
rect 13320 13404 13326 13416
rect 20530 13404 20536 13416
rect 20588 13404 20594 13456
rect 20824 13444 20852 13472
rect 23658 13444 23664 13456
rect 20824 13416 23664 13444
rect 23658 13404 23664 13416
rect 23716 13404 23722 13456
rect 26436 13453 26464 13484
rect 29362 13472 29368 13484
rect 29420 13472 29426 13524
rect 26421 13447 26479 13453
rect 26421 13413 26433 13447
rect 26467 13413 26479 13447
rect 26421 13407 26479 13413
rect 26510 13404 26516 13456
rect 26568 13444 26574 13456
rect 27617 13447 27675 13453
rect 27617 13444 27629 13447
rect 26568 13416 27629 13444
rect 26568 13404 26574 13416
rect 27617 13413 27629 13416
rect 27663 13413 27675 13447
rect 27617 13407 27675 13413
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 2038 13376 2044 13388
rect 1719 13348 2044 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 2038 13336 2044 13348
rect 2096 13376 2102 13388
rect 2498 13376 2504 13388
rect 2096 13348 2504 13376
rect 2096 13336 2102 13348
rect 2498 13336 2504 13348
rect 2556 13376 2562 13388
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 2556 13348 4077 13376
rect 2556 13336 2562 13348
rect 4065 13345 4077 13348
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 8573 13379 8631 13385
rect 4387 13348 8524 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 6546 13308 6552 13320
rect 6507 13280 6552 13308
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 8496 13308 8524 13348
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 11422 13376 11428 13388
rect 8619 13348 11428 13376
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 11977 13379 12035 13385
rect 11977 13345 11989 13379
rect 12023 13376 12035 13379
rect 12618 13376 12624 13388
rect 12023 13348 12624 13376
rect 12023 13345 12035 13348
rect 11977 13339 12035 13345
rect 12618 13336 12624 13348
rect 12676 13376 12682 13388
rect 13170 13376 13176 13388
rect 12676 13348 13176 13376
rect 12676 13336 12682 13348
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 13630 13336 13636 13388
rect 13688 13376 13694 13388
rect 13725 13379 13783 13385
rect 13725 13376 13737 13379
rect 13688 13348 13737 13376
rect 13688 13336 13694 13348
rect 13725 13345 13737 13348
rect 13771 13376 13783 13379
rect 13814 13376 13820 13388
rect 13771 13348 13820 13376
rect 13771 13345 13783 13348
rect 13725 13339 13783 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13376 15439 13379
rect 15562 13376 15568 13388
rect 15427 13348 15568 13376
rect 15427 13345 15439 13348
rect 15381 13339 15439 13345
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15672 13348 16313 13376
rect 8938 13308 8944 13320
rect 8496 13280 8944 13308
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 9180 13280 9229 13308
rect 9180 13268 9186 13280
rect 9217 13277 9229 13280
rect 9263 13277 9275 13311
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 9217 13271 9275 13277
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 15672 13252 15700 13348
rect 16301 13345 16313 13348
rect 16347 13376 16359 13379
rect 16390 13376 16396 13388
rect 16347 13348 16396 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16666 13376 16672 13388
rect 16627 13348 16672 13376
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16758 13336 16764 13388
rect 16816 13376 16822 13388
rect 17218 13376 17224 13388
rect 16816 13348 17224 13376
rect 16816 13336 16822 13348
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 19150 13376 19156 13388
rect 17420 13348 19156 13376
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17420 13317 17448 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 20990 13376 20996 13388
rect 19300 13348 20208 13376
rect 19300 13336 19306 13348
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 17000 13280 17417 13308
rect 17000 13268 17006 13280
rect 17405 13277 17417 13280
rect 17451 13277 17463 13311
rect 17405 13271 17463 13277
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17552 13280 17597 13308
rect 17552 13268 17558 13280
rect 18874 13268 18880 13320
rect 18932 13308 18938 13320
rect 20180 13317 20208 13348
rect 20457 13348 20996 13376
rect 20165 13311 20223 13317
rect 18932 13280 18977 13308
rect 18932 13268 18938 13280
rect 20165 13277 20177 13311
rect 20211 13308 20223 13311
rect 20254 13308 20260 13320
rect 20211 13280 20260 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 1949 13243 2007 13249
rect 1949 13209 1961 13243
rect 1995 13209 2007 13243
rect 4430 13240 4436 13252
rect 3174 13212 4436 13240
rect 1949 13203 2007 13209
rect 1964 13172 1992 13203
rect 4430 13200 4436 13212
rect 4488 13200 4494 13252
rect 5810 13240 5816 13252
rect 5566 13212 5816 13240
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 6086 13240 6092 13252
rect 5999 13212 6092 13240
rect 6086 13200 6092 13212
rect 6144 13240 6150 13252
rect 6730 13240 6736 13252
rect 6144 13212 6736 13240
rect 6144 13200 6150 13212
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 6880 13212 6925 13240
rect 6880 13200 6886 13212
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 7156 13212 7314 13240
rect 7156 13200 7162 13212
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 9030 13240 9036 13252
rect 8444 13212 9036 13240
rect 8444 13200 8450 13212
rect 9030 13200 9036 13212
rect 9088 13240 9094 13252
rect 9493 13243 9551 13249
rect 9493 13240 9505 13243
rect 9088 13212 9505 13240
rect 9088 13200 9094 13212
rect 9493 13209 9505 13212
rect 9539 13209 9551 13243
rect 10870 13240 10876 13252
rect 10718 13212 10876 13240
rect 9493 13203 9551 13209
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 11241 13243 11299 13249
rect 11241 13209 11253 13243
rect 11287 13240 11299 13243
rect 12066 13240 12072 13252
rect 11287 13212 12072 13240
rect 11287 13209 11299 13212
rect 11241 13203 11299 13209
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 12986 13200 12992 13252
rect 13044 13200 13050 13252
rect 14369 13243 14427 13249
rect 14369 13209 14381 13243
rect 14415 13209 14427 13243
rect 14369 13203 14427 13209
rect 2958 13172 2964 13184
rect 1964 13144 2964 13172
rect 2958 13132 2964 13144
rect 3016 13172 3022 13184
rect 3510 13172 3516 13184
rect 3016 13144 3516 13172
rect 3016 13132 3022 13144
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 14274 13172 14280 13184
rect 5040 13144 14280 13172
rect 5040 13132 5046 13144
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14384 13172 14412 13203
rect 14458 13200 14464 13252
rect 14516 13240 14522 13252
rect 14516 13212 14561 13240
rect 14516 13200 14522 13212
rect 15654 13200 15660 13252
rect 15712 13200 15718 13252
rect 16390 13240 16396 13252
rect 16351 13212 16396 13240
rect 16390 13200 16396 13212
rect 16448 13200 16454 13252
rect 16666 13240 16672 13252
rect 16500 13212 16672 13240
rect 16022 13172 16028 13184
rect 14384 13144 16028 13172
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 16500 13172 16528 13212
rect 16666 13200 16672 13212
rect 16724 13240 16730 13252
rect 17954 13240 17960 13252
rect 16724 13212 17960 13240
rect 16724 13200 16730 13212
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 18230 13240 18236 13252
rect 18191 13212 18236 13240
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 18325 13243 18383 13249
rect 18325 13209 18337 13243
rect 18371 13240 18383 13243
rect 18598 13240 18604 13252
rect 18371 13212 18604 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 18598 13200 18604 13212
rect 18656 13200 18662 13252
rect 18690 13200 18696 13252
rect 18748 13240 18754 13252
rect 18966 13240 18972 13252
rect 18748 13212 18972 13240
rect 18748 13200 18754 13212
rect 18966 13200 18972 13212
rect 19024 13200 19030 13252
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 19334 13240 19340 13252
rect 19116 13212 19340 13240
rect 19116 13200 19122 13212
rect 19334 13200 19340 13212
rect 19392 13200 19398 13252
rect 19518 13240 19524 13252
rect 19479 13212 19524 13240
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13209 19671 13243
rect 19613 13203 19671 13209
rect 16356 13144 16528 13172
rect 16356 13132 16362 13144
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 19536 13172 19564 13200
rect 16632 13144 19564 13172
rect 19628 13172 19656 13203
rect 19886 13200 19892 13252
rect 19944 13240 19950 13252
rect 20457 13240 20485 13348
rect 20990 13336 20996 13348
rect 21048 13336 21054 13388
rect 21634 13376 21640 13388
rect 21547 13348 21640 13376
rect 21634 13336 21640 13348
rect 21692 13376 21698 13388
rect 22094 13376 22100 13388
rect 21692 13348 22100 13376
rect 21692 13336 21698 13348
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 22278 13336 22284 13388
rect 22336 13376 22342 13388
rect 23566 13376 23572 13388
rect 22336 13348 23572 13376
rect 22336 13336 22342 13348
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 23676 13376 23704 13404
rect 28261 13379 28319 13385
rect 28261 13376 28273 13379
rect 23676 13348 24624 13376
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 20901 13311 20959 13317
rect 20901 13308 20913 13311
rect 20864 13280 20913 13308
rect 20864 13268 20870 13280
rect 20901 13277 20913 13280
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 22738 13268 22744 13320
rect 22796 13308 22802 13320
rect 23109 13311 23167 13317
rect 23109 13308 23121 13311
rect 22796 13280 23121 13308
rect 22796 13268 22802 13280
rect 23109 13277 23121 13280
rect 23155 13308 23167 13311
rect 23753 13311 23811 13317
rect 23155 13280 23704 13308
rect 23155 13277 23167 13280
rect 23109 13271 23167 13277
rect 19944 13212 20485 13240
rect 19944 13200 19950 13212
rect 20530 13200 20536 13252
rect 20588 13240 20594 13252
rect 21729 13243 21787 13249
rect 20588 13212 21588 13240
rect 20588 13200 20594 13212
rect 20898 13172 20904 13184
rect 19628 13144 20904 13172
rect 16632 13132 16638 13144
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 21560 13172 21588 13212
rect 21729 13209 21741 13243
rect 21775 13240 21787 13243
rect 22554 13240 22560 13252
rect 21775 13212 22560 13240
rect 21775 13209 21787 13212
rect 21729 13203 21787 13209
rect 22554 13200 22560 13212
rect 22612 13200 22618 13252
rect 22649 13243 22707 13249
rect 22649 13209 22661 13243
rect 22695 13240 22707 13243
rect 23290 13240 23296 13252
rect 22695 13212 23296 13240
rect 22695 13209 22707 13212
rect 22649 13203 22707 13209
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 22462 13172 22468 13184
rect 21560 13144 22468 13172
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 23676 13172 23704 13280
rect 23753 13277 23765 13311
rect 23799 13308 23811 13311
rect 23842 13308 23848 13320
rect 23799 13280 23848 13308
rect 23799 13277 23811 13280
rect 23753 13271 23811 13277
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 24596 13317 24624 13348
rect 26620 13348 28273 13376
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 24670 13240 24676 13252
rect 24631 13212 24676 13240
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 25682 13200 25688 13252
rect 25740 13240 25746 13252
rect 25869 13243 25927 13249
rect 25869 13240 25881 13243
rect 25740 13212 25881 13240
rect 25740 13200 25746 13212
rect 25869 13209 25881 13212
rect 25915 13209 25927 13243
rect 25869 13203 25927 13209
rect 25961 13243 26019 13249
rect 25961 13209 25973 13243
rect 26007 13209 26019 13243
rect 25961 13203 26019 13209
rect 25498 13172 25504 13184
rect 23676 13144 25504 13172
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 25976 13172 26004 13203
rect 26620 13172 26648 13348
rect 28261 13345 28273 13348
rect 28307 13345 28319 13379
rect 28261 13339 28319 13345
rect 28166 13308 28172 13320
rect 28079 13280 28172 13308
rect 28166 13268 28172 13280
rect 28224 13308 28230 13320
rect 28442 13308 28448 13320
rect 28224 13280 28448 13308
rect 28224 13268 28230 13280
rect 28442 13268 28448 13280
rect 28500 13268 28506 13320
rect 28626 13268 28632 13320
rect 28684 13308 28690 13320
rect 28813 13311 28871 13317
rect 28813 13308 28825 13311
rect 28684 13280 28825 13308
rect 28684 13268 28690 13280
rect 28813 13277 28825 13280
rect 28859 13277 28871 13311
rect 29730 13308 29736 13320
rect 29643 13280 29736 13308
rect 28813 13271 28871 13277
rect 29730 13268 29736 13280
rect 29788 13308 29794 13320
rect 29914 13308 29920 13320
rect 29788 13280 29920 13308
rect 29788 13268 29794 13280
rect 29914 13268 29920 13280
rect 29972 13268 29978 13320
rect 27062 13240 27068 13252
rect 27023 13212 27068 13240
rect 27062 13200 27068 13212
rect 27120 13200 27126 13252
rect 27157 13243 27215 13249
rect 27157 13209 27169 13243
rect 27203 13209 27215 13243
rect 29825 13243 29883 13249
rect 29825 13240 29837 13243
rect 27157 13203 27215 13209
rect 27816 13212 29837 13240
rect 25976 13144 26648 13172
rect 27172 13172 27200 13203
rect 27816 13172 27844 13212
rect 29825 13209 29837 13212
rect 29871 13209 29883 13243
rect 29825 13203 29883 13209
rect 28902 13172 28908 13184
rect 27172 13144 27844 13172
rect 28863 13144 28908 13172
rect 28902 13132 28908 13144
rect 28960 13132 28966 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 8478 12968 8484 12980
rect 4488 12940 8484 12968
rect 4488 12928 4494 12940
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 11238 12968 11244 12980
rect 9140 12940 11244 12968
rect 934 12860 940 12912
rect 992 12900 998 12912
rect 2409 12903 2467 12909
rect 2409 12900 2421 12903
rect 992 12872 2421 12900
rect 992 12860 998 12872
rect 2409 12869 2421 12872
rect 2455 12869 2467 12903
rect 4154 12900 4160 12912
rect 4115 12872 4160 12900
rect 2409 12863 2467 12869
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 4801 12903 4859 12909
rect 4801 12900 4813 12903
rect 4540 12872 4813 12900
rect 4540 12844 4568 12872
rect 4801 12869 4813 12872
rect 4847 12869 4859 12903
rect 6914 12900 6920 12912
rect 6875 12872 6920 12900
rect 4801 12863 4859 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 8202 12900 8208 12912
rect 8142 12872 8208 12900
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2133 12835 2191 12841
rect 2133 12832 2145 12835
rect 2096 12804 2145 12832
rect 2096 12792 2102 12804
rect 2133 12801 2145 12804
rect 2179 12801 2191 12835
rect 2133 12795 2191 12801
rect 3528 12628 3556 12818
rect 4522 12792 4528 12844
rect 4580 12792 4586 12844
rect 5994 12832 6000 12844
rect 5736 12804 6000 12832
rect 3602 12724 3608 12776
rect 3660 12764 3666 12776
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 3660 12736 4721 12764
rect 3660 12724 3666 12736
rect 4709 12733 4721 12736
rect 4755 12764 4767 12767
rect 5534 12764 5540 12776
rect 4755 12736 5540 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5736 12773 5764 12804
rect 5994 12792 6000 12804
rect 6052 12792 6058 12844
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12832 8723 12835
rect 8938 12832 8944 12844
rect 8711 12804 8944 12832
rect 8711 12801 8723 12804
rect 8665 12795 8723 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 9140 12841 9168 12940
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 11940 12940 16344 12968
rect 11940 12928 11946 12940
rect 9401 12903 9459 12909
rect 9401 12869 9413 12903
rect 9447 12900 9459 12903
rect 9490 12900 9496 12912
rect 9447 12872 9496 12900
rect 9447 12869 9459 12872
rect 9401 12863 9459 12869
rect 9490 12860 9496 12872
rect 9548 12860 9554 12912
rect 10778 12900 10784 12912
rect 10626 12872 10784 12900
rect 10778 12860 10784 12872
rect 10836 12860 10842 12912
rect 13446 12860 13452 12912
rect 13504 12900 13510 12912
rect 13722 12900 13728 12912
rect 13504 12872 13728 12900
rect 13504 12860 13510 12872
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 14461 12903 14519 12909
rect 14461 12900 14473 12903
rect 14148 12872 14473 12900
rect 14148 12860 14154 12872
rect 14461 12869 14473 12872
rect 14507 12869 14519 12903
rect 14461 12863 14519 12869
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 15746 12900 15752 12912
rect 15427 12872 15752 12900
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 16316 12900 16344 12940
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 22278 12968 22284 12980
rect 16448 12940 22284 12968
rect 16448 12928 16454 12940
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 22554 12928 22560 12980
rect 22612 12968 22618 12980
rect 22612 12940 22876 12968
rect 22612 12928 22618 12940
rect 16758 12900 16764 12912
rect 16316 12872 16764 12900
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 17034 12900 17040 12912
rect 16995 12872 17040 12900
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 17129 12903 17187 12909
rect 17129 12869 17141 12903
rect 17175 12900 17187 12903
rect 17862 12900 17868 12912
rect 17175 12872 17868 12900
rect 17175 12869 17187 12872
rect 17129 12863 17187 12869
rect 17862 12860 17868 12872
rect 17920 12860 17926 12912
rect 18230 12900 18236 12912
rect 18064 12872 18236 12900
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 13170 12792 13176 12844
rect 13228 12792 13234 12844
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 15838 12832 15844 12844
rect 13412 12804 13860 12832
rect 15799 12804 15844 12832
rect 13412 12792 13418 12804
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 5810 12724 5816 12776
rect 5868 12764 5874 12776
rect 6546 12764 6552 12776
rect 5868 12736 6552 12764
rect 5868 12724 5874 12736
rect 6546 12724 6552 12736
rect 6604 12764 6610 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6604 12736 6653 12764
rect 6604 12724 6610 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 10594 12764 10600 12776
rect 6641 12727 6699 12733
rect 6748 12736 10600 12764
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 6748 12696 6776 12736
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10962 12724 10968 12776
rect 11020 12764 11026 12776
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 11020 12736 11161 12764
rect 11020 12724 11026 12736
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 11698 12764 11704 12776
rect 11296 12736 11704 12764
rect 11296 12724 11302 12736
rect 11698 12724 11704 12736
rect 11756 12764 11762 12776
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11756 12736 11805 12764
rect 11756 12724 11762 12736
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 13630 12764 13636 12776
rect 12115 12736 13636 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 13630 12724 13636 12736
rect 13688 12724 13694 12776
rect 13832 12773 13860 12804
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 16298 12832 16304 12844
rect 16040 12804 16304 12832
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12733 13875 12767
rect 13817 12727 13875 12733
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 14642 12764 14648 12776
rect 14415 12736 14648 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 14642 12724 14648 12736
rect 14700 12764 14706 12776
rect 16040 12764 16068 12804
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 18064 12832 18092 12872
rect 18230 12860 18236 12872
rect 18288 12860 18294 12912
rect 18325 12903 18383 12909
rect 18325 12869 18337 12903
rect 18371 12900 18383 12903
rect 20165 12903 20223 12909
rect 18371 12872 19921 12900
rect 18371 12869 18383 12872
rect 18325 12863 18383 12869
rect 17880 12804 18092 12832
rect 17880 12776 17908 12804
rect 14700 12736 16068 12764
rect 14700 12724 14706 12736
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 17034 12764 17040 12776
rect 16172 12736 17040 12764
rect 16172 12724 16178 12736
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17494 12764 17500 12776
rect 17455 12736 17500 12764
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 17862 12724 17868 12776
rect 17920 12724 17926 12776
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 18156 12736 18245 12764
rect 4120 12668 6776 12696
rect 4120 12656 4126 12668
rect 8478 12656 8484 12708
rect 8536 12696 8542 12708
rect 9030 12696 9036 12708
rect 8536 12668 9036 12696
rect 8536 12656 8542 12668
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 13078 12656 13084 12708
rect 13136 12696 13142 12708
rect 13722 12696 13728 12708
rect 13136 12668 13728 12696
rect 13136 12656 13142 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 16482 12656 16488 12708
rect 16540 12696 16546 12708
rect 18156 12696 18184 12736
rect 18233 12733 18245 12736
rect 18279 12764 18291 12767
rect 19058 12764 19064 12776
rect 18279 12736 18368 12764
rect 19019 12736 19064 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 16540 12668 18184 12696
rect 16540 12656 16546 12668
rect 18340 12640 18368 12736
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 19150 12724 19156 12776
rect 19208 12764 19214 12776
rect 19702 12764 19708 12776
rect 19208 12736 19708 12764
rect 19208 12724 19214 12736
rect 19702 12724 19708 12736
rect 19760 12724 19766 12776
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 18472 12668 18920 12696
rect 18472 12656 18478 12668
rect 11882 12628 11888 12640
rect 3528 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 16206 12628 16212 12640
rect 12492 12600 16212 12628
rect 12492 12588 12498 12600
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 18138 12628 18144 12640
rect 17092 12600 18144 12628
rect 17092 12588 17098 12600
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18322 12588 18328 12640
rect 18380 12588 18386 12640
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 18782 12628 18788 12640
rect 18656 12600 18788 12628
rect 18656 12588 18662 12600
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 18892 12628 18920 12668
rect 18966 12656 18972 12708
rect 19024 12696 19030 12708
rect 19794 12696 19800 12708
rect 19024 12668 19800 12696
rect 19024 12656 19030 12668
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 19893 12696 19921 12872
rect 20165 12869 20177 12903
rect 20211 12900 20223 12903
rect 20530 12900 20536 12912
rect 20211 12872 20536 12900
rect 20211 12869 20223 12872
rect 20165 12863 20223 12869
rect 20530 12860 20536 12872
rect 20588 12860 20594 12912
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 21085 12903 21143 12909
rect 21085 12900 21097 12903
rect 20680 12872 21097 12900
rect 20680 12860 20686 12872
rect 21085 12869 21097 12872
rect 21131 12900 21143 12903
rect 21450 12900 21456 12912
rect 21131 12872 21456 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 21450 12860 21456 12872
rect 21508 12860 21514 12912
rect 21910 12860 21916 12912
rect 21968 12900 21974 12912
rect 22097 12903 22155 12909
rect 22097 12900 22109 12903
rect 21968 12872 22109 12900
rect 21968 12860 21974 12872
rect 22097 12869 22109 12872
rect 22143 12869 22155 12903
rect 22097 12863 22155 12869
rect 22189 12903 22247 12909
rect 22189 12869 22201 12903
rect 22235 12900 22247 12903
rect 22738 12900 22744 12912
rect 22235 12872 22744 12900
rect 22235 12869 22247 12872
rect 22189 12863 22247 12869
rect 22738 12860 22744 12872
rect 22796 12860 22802 12912
rect 22848 12900 22876 12940
rect 23014 12928 23020 12980
rect 23072 12968 23078 12980
rect 23293 12971 23351 12977
rect 23293 12968 23305 12971
rect 23072 12940 23305 12968
rect 23072 12928 23078 12940
rect 23293 12937 23305 12940
rect 23339 12937 23351 12971
rect 23293 12931 23351 12937
rect 23937 12971 23995 12977
rect 23937 12937 23949 12971
rect 23983 12968 23995 12971
rect 24026 12968 24032 12980
rect 23983 12940 24032 12968
rect 23983 12937 23995 12940
rect 23937 12931 23995 12937
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 24578 12928 24584 12980
rect 24636 12968 24642 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 24636 12940 25237 12968
rect 24636 12928 24642 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 29178 12968 29184 12980
rect 25225 12931 25283 12937
rect 27724 12940 29184 12968
rect 26053 12903 26111 12909
rect 22848 12872 24900 12900
rect 24872 12844 24900 12872
rect 26053 12869 26065 12903
rect 26099 12900 26111 12903
rect 27249 12903 27307 12909
rect 27249 12900 27261 12903
rect 26099 12872 27261 12900
rect 26099 12869 26111 12872
rect 26053 12863 26111 12869
rect 27249 12869 27261 12872
rect 27295 12869 27307 12903
rect 27249 12863 27307 12869
rect 21726 12832 21732 12844
rect 21100 12804 21732 12832
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 21100 12764 21128 12804
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 23014 12792 23020 12844
rect 23072 12832 23078 12844
rect 23201 12835 23259 12841
rect 23201 12832 23213 12835
rect 23072 12804 23213 12832
rect 23072 12792 23078 12804
rect 23201 12801 23213 12804
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 20119 12736 21128 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 21174 12724 21180 12776
rect 21232 12764 21238 12776
rect 22370 12764 22376 12776
rect 21232 12736 22376 12764
rect 21232 12724 21238 12736
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 22741 12767 22799 12773
rect 22741 12733 22753 12767
rect 22787 12764 22799 12767
rect 22922 12764 22928 12776
rect 22787 12736 22928 12764
rect 22787 12733 22799 12736
rect 22741 12727 22799 12733
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 23216 12764 23244 12795
rect 23474 12792 23480 12844
rect 23532 12832 23538 12844
rect 23845 12835 23903 12841
rect 23845 12832 23857 12835
rect 23532 12804 23857 12832
rect 23532 12792 23538 12804
rect 23845 12801 23857 12804
rect 23891 12801 23903 12835
rect 23845 12795 23903 12801
rect 24489 12835 24547 12841
rect 24489 12801 24501 12835
rect 24535 12832 24547 12835
rect 24762 12832 24768 12844
rect 24535 12804 24768 12832
rect 24535 12801 24547 12804
rect 24489 12795 24547 12801
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 24854 12792 24860 12844
rect 24912 12792 24918 12844
rect 25133 12835 25191 12841
rect 25133 12801 25145 12835
rect 25179 12832 25191 12835
rect 25222 12832 25228 12844
rect 25179 12804 25228 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 25222 12792 25228 12804
rect 25280 12792 25286 12844
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12832 27215 12835
rect 27522 12832 27528 12844
rect 27203 12804 27528 12832
rect 27203 12801 27215 12804
rect 27157 12795 27215 12801
rect 27522 12792 27528 12804
rect 27580 12792 27586 12844
rect 25958 12764 25964 12776
rect 23216 12736 25820 12764
rect 25919 12736 25964 12764
rect 20714 12696 20720 12708
rect 19893 12668 20720 12696
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 21634 12696 21640 12708
rect 20864 12668 21640 12696
rect 20864 12656 20870 12668
rect 21634 12656 21640 12668
rect 21692 12656 21698 12708
rect 22278 12656 22284 12708
rect 22336 12696 22342 12708
rect 24581 12699 24639 12705
rect 24581 12696 24593 12699
rect 22336 12668 24593 12696
rect 22336 12656 22342 12668
rect 24581 12665 24593 12668
rect 24627 12696 24639 12699
rect 25682 12696 25688 12708
rect 24627 12668 25688 12696
rect 24627 12665 24639 12668
rect 24581 12659 24639 12665
rect 25682 12656 25688 12668
rect 25740 12656 25746 12708
rect 25792 12696 25820 12736
rect 25958 12724 25964 12736
rect 26016 12724 26022 12776
rect 26605 12767 26663 12773
rect 26605 12733 26617 12767
rect 26651 12764 26663 12767
rect 27724 12764 27752 12940
rect 29178 12928 29184 12940
rect 29236 12928 29242 12980
rect 30374 12928 30380 12980
rect 30432 12968 30438 12980
rect 32401 12971 32459 12977
rect 32401 12968 32413 12971
rect 30432 12940 32413 12968
rect 30432 12928 30438 12940
rect 32401 12937 32413 12940
rect 32447 12937 32459 12971
rect 32401 12931 32459 12937
rect 27982 12900 27988 12912
rect 27943 12872 27988 12900
rect 27982 12860 27988 12872
rect 28040 12860 28046 12912
rect 30834 12900 30840 12912
rect 30795 12872 30840 12900
rect 30834 12860 30840 12872
rect 30892 12860 30898 12912
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12832 32367 12835
rect 33962 12832 33968 12844
rect 32355 12804 33968 12832
rect 32355 12801 32367 12804
rect 32309 12795 32367 12801
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 36446 12792 36452 12844
rect 36504 12832 36510 12844
rect 38013 12835 38071 12841
rect 38013 12832 38025 12835
rect 36504 12804 38025 12832
rect 36504 12792 36510 12804
rect 38013 12801 38025 12804
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 26651 12736 27752 12764
rect 27893 12767 27951 12773
rect 26651 12733 26663 12736
rect 26605 12727 26663 12733
rect 27893 12733 27905 12767
rect 27939 12733 27951 12767
rect 27893 12727 27951 12733
rect 26234 12696 26240 12708
rect 25792 12668 26240 12696
rect 26234 12656 26240 12668
rect 26292 12656 26298 12708
rect 27908 12696 27936 12727
rect 28074 12724 28080 12776
rect 28132 12764 28138 12776
rect 28169 12767 28227 12773
rect 28169 12764 28181 12767
rect 28132 12736 28181 12764
rect 28132 12724 28138 12736
rect 28169 12733 28181 12736
rect 28215 12733 28227 12767
rect 30742 12764 30748 12776
rect 30703 12736 30748 12764
rect 28169 12727 28227 12733
rect 30742 12724 30748 12736
rect 30800 12724 30806 12776
rect 31662 12764 31668 12776
rect 31623 12736 31668 12764
rect 31662 12724 31668 12736
rect 31720 12724 31726 12776
rect 31018 12696 31024 12708
rect 27908 12668 31024 12696
rect 31018 12656 31024 12668
rect 31076 12656 31082 12708
rect 26142 12628 26148 12640
rect 18892 12600 26148 12628
rect 26142 12588 26148 12600
rect 26200 12628 26206 12640
rect 27062 12628 27068 12640
rect 26200 12600 27068 12628
rect 26200 12588 26206 12600
rect 27062 12588 27068 12600
rect 27120 12588 27126 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1936 12427 1994 12433
rect 1936 12393 1948 12427
rect 1982 12424 1994 12427
rect 1982 12396 3832 12424
rect 1982 12393 1994 12396
rect 1936 12387 1994 12393
rect 3804 12356 3832 12396
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4062 12424 4068 12436
rect 3936 12396 4068 12424
rect 3936 12384 3942 12396
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8478 12424 8484 12436
rect 8352 12396 8484 12424
rect 8352 12384 8358 12396
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 23474 12424 23480 12436
rect 8956 12396 13952 12424
rect 5736 12356 5764 12384
rect 3804 12328 5764 12356
rect 7834 12316 7840 12368
rect 7892 12356 7898 12368
rect 8956 12356 8984 12396
rect 13924 12368 13952 12396
rect 14016 12396 23480 12424
rect 7892 12328 8984 12356
rect 7892 12316 7898 12328
rect 9030 12316 9036 12368
rect 9088 12356 9094 12368
rect 10778 12356 10784 12368
rect 9088 12328 10784 12356
rect 9088 12316 9094 12328
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 12894 12316 12900 12368
rect 12952 12356 12958 12368
rect 13078 12356 13084 12368
rect 12952 12328 13084 12356
rect 12952 12316 12958 12328
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 13906 12316 13912 12368
rect 13964 12316 13970 12368
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 1673 12291 1731 12297
rect 1673 12288 1685 12291
rect 1636 12260 1685 12288
rect 1636 12248 1642 12260
rect 1673 12257 1685 12260
rect 1719 12288 1731 12291
rect 2038 12288 2044 12300
rect 1719 12260 2044 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 5077 12291 5135 12297
rect 3896 12260 5028 12288
rect 3896 12220 3924 12260
rect 3082 12192 3924 12220
rect 5000 12220 5028 12260
rect 5077 12257 5089 12291
rect 5123 12288 5135 12291
rect 5166 12288 5172 12300
rect 5123 12260 5172 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12288 5779 12291
rect 6730 12288 6736 12300
rect 5767 12260 6736 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 5626 12220 5632 12232
rect 5000 12192 5632 12220
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 3602 12112 3608 12164
rect 3660 12152 3666 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 3660 12124 4077 12152
rect 3660 12112 3666 12124
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4065 12115 4123 12121
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4212 12124 4257 12152
rect 4212 12112 4218 12124
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 4890 12152 4896 12164
rect 4764 12124 4896 12152
rect 4764 12112 4770 12124
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 2866 12084 2872 12096
rect 1912 12056 2872 12084
rect 1912 12044 1918 12056
rect 2866 12044 2872 12056
rect 2924 12084 2930 12096
rect 3421 12087 3479 12093
rect 3421 12084 3433 12087
rect 2924 12056 3433 12084
rect 2924 12044 2930 12056
rect 3421 12053 3433 12056
rect 3467 12053 3479 12087
rect 5736 12084 5764 12251
rect 6730 12248 6736 12260
rect 6788 12288 6794 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 6788 12260 9873 12288
rect 6788 12248 6794 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 9861 12251 9919 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11514 12288 11520 12300
rect 11475 12260 11520 12288
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14016 12288 14044 12396
rect 23474 12384 23480 12396
rect 23532 12384 23538 12436
rect 26142 12384 26148 12436
rect 26200 12424 26206 12436
rect 27433 12427 27491 12433
rect 27433 12424 27445 12427
rect 26200 12396 27445 12424
rect 26200 12384 26206 12396
rect 27433 12393 27445 12396
rect 27479 12393 27491 12427
rect 27433 12387 27491 12393
rect 34885 12427 34943 12433
rect 34885 12393 34897 12427
rect 34931 12424 34943 12427
rect 36446 12424 36452 12436
rect 34931 12396 36452 12424
rect 34931 12393 34943 12396
rect 34885 12387 34943 12393
rect 36446 12384 36452 12396
rect 36504 12384 36510 12436
rect 14550 12316 14556 12368
rect 14608 12356 14614 12368
rect 14734 12356 14740 12368
rect 14608 12328 14740 12356
rect 14608 12316 14614 12328
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 17678 12356 17684 12368
rect 15528 12328 17684 12356
rect 15528 12316 15534 12328
rect 17678 12316 17684 12328
rect 17736 12316 17742 12368
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 20625 12359 20683 12365
rect 20625 12356 20637 12359
rect 17920 12328 20637 12356
rect 17920 12316 17926 12328
rect 13872 12260 14044 12288
rect 13872 12248 13878 12260
rect 15286 12248 15292 12300
rect 15344 12288 15350 12300
rect 15344 12260 15700 12288
rect 15344 12248 15350 12260
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8294 12220 8300 12232
rect 7791 12192 8300 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8570 12220 8576 12232
rect 8531 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9582 12220 9588 12232
rect 9272 12192 9588 12220
rect 9272 12180 9278 12192
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 15672 12229 15700 12260
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16632 12260 16865 12288
rect 16632 12248 16638 12260
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 16853 12251 16911 12257
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17972 12288 18000 12328
rect 20625 12325 20637 12328
rect 20671 12325 20683 12359
rect 20625 12319 20683 12325
rect 20898 12316 20904 12368
rect 20956 12356 20962 12368
rect 21174 12356 21180 12368
rect 20956 12328 21180 12356
rect 20956 12316 20962 12328
rect 21174 12316 21180 12328
rect 21232 12316 21238 12368
rect 21269 12359 21327 12365
rect 21269 12325 21281 12359
rect 21315 12356 21327 12359
rect 24673 12359 24731 12365
rect 21315 12328 22416 12356
rect 21315 12325 21327 12328
rect 21269 12319 21327 12325
rect 17092 12260 18000 12288
rect 17092 12248 17098 12260
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 20073 12291 20131 12297
rect 18104 12260 18736 12288
rect 18104 12248 18110 12260
rect 10505 12223 10563 12229
rect 10505 12220 10517 12223
rect 10284 12192 10517 12220
rect 10284 12180 10290 12192
rect 10505 12189 10517 12192
rect 10551 12189 10563 12223
rect 15657 12223 15715 12229
rect 12650 12192 15608 12220
rect 10505 12183 10563 12189
rect 5997 12155 6055 12161
rect 5997 12121 6009 12155
rect 6043 12121 6055 12155
rect 8110 12152 8116 12164
rect 7222 12124 8116 12152
rect 5997 12115 6055 12121
rect 5810 12084 5816 12096
rect 5736 12056 5816 12084
rect 3421 12047 3479 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6012 12084 6040 12115
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 8386 12152 8392 12164
rect 8347 12124 8392 12152
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 9125 12155 9183 12161
rect 9125 12121 9137 12155
rect 9171 12152 9183 12155
rect 9674 12152 9680 12164
rect 9171 12124 9680 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9674 12112 9680 12124
rect 9732 12152 9738 12164
rect 10134 12152 10140 12164
rect 9732 12124 10140 12152
rect 9732 12112 9738 12124
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 13265 12155 13323 12161
rect 13265 12121 13277 12155
rect 13311 12152 13323 12155
rect 13354 12152 13360 12164
rect 13311 12124 13360 12152
rect 13311 12121 13323 12124
rect 13265 12115 13323 12121
rect 13354 12112 13360 12124
rect 13412 12112 13418 12164
rect 14274 12152 14280 12164
rect 14235 12124 14280 12152
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 15010 12152 15016 12164
rect 14971 12124 15016 12152
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 15580 12152 15608 12192
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 16390 12220 16396 12232
rect 15703 12192 16396 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17862 12220 17868 12232
rect 17543 12192 17868 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 16945 12155 17003 12161
rect 15580 12124 15884 12152
rect 7282 12084 7288 12096
rect 6012 12056 7288 12084
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10284 12056 10609 12084
rect 10284 12044 10290 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 10836 12056 15761 12084
rect 10836 12044 10842 12056
rect 15749 12053 15761 12056
rect 15795 12053 15807 12087
rect 15856 12084 15884 12124
rect 16945 12121 16957 12155
rect 16991 12152 17003 12155
rect 17310 12152 17316 12164
rect 16991 12124 17316 12152
rect 16991 12121 17003 12124
rect 16945 12115 17003 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 17678 12112 17684 12164
rect 17736 12152 17742 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 17736 12124 18061 12152
rect 17736 12112 17742 12124
rect 18049 12121 18061 12124
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 18141 12155 18199 12161
rect 18141 12121 18153 12155
rect 18187 12152 18199 12155
rect 18506 12152 18512 12164
rect 18187 12124 18512 12152
rect 18187 12121 18199 12124
rect 18141 12115 18199 12121
rect 18506 12112 18512 12124
rect 18564 12112 18570 12164
rect 18708 12161 18736 12260
rect 20073 12257 20085 12291
rect 20119 12288 20131 12291
rect 22278 12288 22284 12300
rect 20119 12260 22284 12288
rect 20119 12257 20131 12260
rect 20073 12251 20131 12257
rect 22278 12248 22284 12260
rect 22336 12248 22342 12300
rect 22388 12288 22416 12328
rect 24673 12325 24685 12359
rect 24719 12356 24731 12359
rect 27982 12356 27988 12368
rect 24719 12328 27988 12356
rect 24719 12325 24731 12328
rect 24673 12319 24731 12325
rect 27982 12316 27988 12328
rect 28040 12316 28046 12368
rect 28629 12359 28687 12365
rect 28629 12325 28641 12359
rect 28675 12356 28687 12359
rect 37274 12356 37280 12368
rect 28675 12328 37280 12356
rect 28675 12325 28687 12328
rect 28629 12319 28687 12325
rect 37274 12316 37280 12328
rect 37332 12316 37338 12368
rect 22388 12260 23336 12288
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 21358 12220 21364 12232
rect 21223 12192 21364 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 18693 12155 18751 12161
rect 18693 12121 18705 12155
rect 18739 12152 18751 12155
rect 18782 12152 18788 12164
rect 18739 12124 18788 12152
rect 18739 12121 18751 12124
rect 18693 12115 18751 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 20165 12155 20223 12161
rect 20165 12121 20177 12155
rect 20211 12152 20223 12155
rect 20898 12152 20904 12164
rect 20211 12124 20904 12152
rect 20211 12121 20223 12124
rect 20165 12115 20223 12121
rect 20898 12112 20904 12124
rect 20956 12112 20962 12164
rect 22002 12112 22008 12164
rect 22060 12152 22066 12164
rect 22189 12155 22247 12161
rect 22189 12152 22201 12155
rect 22060 12124 22201 12152
rect 22060 12112 22066 12124
rect 22189 12121 22201 12124
rect 22235 12121 22247 12155
rect 22189 12115 22247 12121
rect 22281 12155 22339 12161
rect 22281 12121 22293 12155
rect 22327 12152 22339 12155
rect 23014 12152 23020 12164
rect 22327 12124 23020 12152
rect 22327 12121 22339 12124
rect 22281 12115 22339 12121
rect 23014 12112 23020 12124
rect 23072 12112 23078 12164
rect 23198 12152 23204 12164
rect 23159 12124 23204 12152
rect 23198 12112 23204 12124
rect 23256 12112 23262 12164
rect 23308 12152 23336 12260
rect 23768 12272 23848 12300
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12220 23719 12223
rect 23768 12220 23796 12272
rect 23842 12248 23848 12272
rect 23900 12248 23906 12300
rect 24946 12248 24952 12300
rect 25004 12288 25010 12300
rect 25869 12291 25927 12297
rect 25869 12288 25881 12291
rect 25004 12260 25881 12288
rect 25004 12248 25010 12260
rect 25869 12257 25881 12260
rect 25915 12257 25927 12291
rect 25869 12251 25927 12257
rect 26050 12248 26056 12300
rect 26108 12288 26114 12300
rect 26145 12291 26203 12297
rect 26145 12288 26157 12291
rect 26108 12260 26157 12288
rect 26108 12248 26114 12260
rect 26145 12257 26157 12260
rect 26191 12288 26203 12291
rect 26191 12260 30696 12288
rect 26191 12257 26203 12260
rect 26145 12251 26203 12257
rect 24302 12220 24308 12232
rect 23707 12192 24308 12220
rect 23707 12189 23719 12192
rect 23661 12183 23719 12189
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 24578 12220 24584 12232
rect 24539 12192 24584 12220
rect 24578 12180 24584 12192
rect 24636 12180 24642 12232
rect 24670 12180 24676 12232
rect 24728 12220 24734 12232
rect 27338 12220 27344 12232
rect 24728 12192 25268 12220
rect 27299 12192 27344 12220
rect 24728 12180 24734 12192
rect 25130 12152 25136 12164
rect 23308 12124 25136 12152
rect 25130 12112 25136 12124
rect 25188 12112 25194 12164
rect 25240 12152 25268 12192
rect 27338 12180 27344 12192
rect 27396 12180 27402 12232
rect 30668 12220 30696 12260
rect 30742 12248 30748 12300
rect 30800 12288 30806 12300
rect 30929 12291 30987 12297
rect 30929 12288 30941 12291
rect 30800 12260 30941 12288
rect 30800 12248 30806 12260
rect 30929 12257 30941 12260
rect 30975 12257 30987 12291
rect 30929 12251 30987 12257
rect 31662 12220 31668 12232
rect 30668 12192 31668 12220
rect 31662 12180 31668 12192
rect 31720 12180 31726 12232
rect 34054 12180 34060 12232
rect 34112 12220 34118 12232
rect 35069 12223 35127 12229
rect 35069 12220 35081 12223
rect 34112 12192 35081 12220
rect 34112 12180 34118 12192
rect 35069 12189 35081 12192
rect 35115 12189 35127 12223
rect 35069 12183 35127 12189
rect 25961 12155 26019 12161
rect 25961 12152 25973 12155
rect 25240 12124 25973 12152
rect 25961 12121 25973 12124
rect 26007 12121 26019 12155
rect 25961 12115 26019 12121
rect 26418 12112 26424 12164
rect 26476 12152 26482 12164
rect 26970 12152 26976 12164
rect 26476 12124 26976 12152
rect 26476 12112 26482 12124
rect 26970 12112 26976 12124
rect 27028 12112 27034 12164
rect 28445 12155 28503 12161
rect 28445 12121 28457 12155
rect 28491 12121 28503 12155
rect 28445 12115 28503 12121
rect 21910 12084 21916 12096
rect 15856 12056 21916 12084
rect 15749 12047 15807 12053
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 23750 12084 23756 12096
rect 23711 12056 23756 12084
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 27154 12084 27160 12096
rect 23992 12056 27160 12084
rect 23992 12044 23998 12056
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 27706 12044 27712 12096
rect 27764 12084 27770 12096
rect 28460 12084 28488 12115
rect 27764 12056 28488 12084
rect 27764 12044 27770 12056
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 750 11840 756 11892
rect 808 11880 814 11892
rect 808 11852 3188 11880
rect 808 11840 814 11852
rect 2406 11772 2412 11824
rect 2464 11772 2470 11824
rect 3160 11812 3188 11852
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3329 11883 3387 11889
rect 3329 11880 3341 11883
rect 3292 11852 3341 11880
rect 3292 11840 3298 11852
rect 3329 11849 3341 11852
rect 3375 11849 3387 11883
rect 3329 11843 3387 11849
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3786 11880 3792 11892
rect 3568 11852 3792 11880
rect 3568 11840 3574 11852
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 5166 11880 5172 11892
rect 3936 11852 5172 11880
rect 3936 11840 3942 11852
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 6822 11880 6828 11892
rect 6012 11852 6828 11880
rect 4154 11812 4160 11824
rect 3160 11784 4160 11812
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 6012 11821 6040 11852
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 8481 11883 8539 11889
rect 8481 11849 8493 11883
rect 8527 11880 8539 11883
rect 8662 11880 8668 11892
rect 8527 11852 8668 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 8849 11883 8907 11889
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 9306 11880 9312 11892
rect 8895 11852 9312 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9306 11840 9312 11852
rect 9364 11880 9370 11892
rect 9364 11852 16804 11880
rect 9364 11840 9370 11852
rect 5997 11815 6055 11821
rect 5997 11781 6009 11815
rect 6043 11781 6055 11815
rect 9030 11812 9036 11824
rect 8234 11784 9036 11812
rect 5997 11775 6055 11781
rect 9030 11772 9036 11784
rect 9088 11772 9094 11824
rect 9416 11821 9444 11852
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11781 9459 11815
rect 9401 11775 9459 11781
rect 11514 11772 11520 11824
rect 11572 11812 11578 11824
rect 11572 11784 12650 11812
rect 11572 11772 11578 11784
rect 13446 11772 13452 11824
rect 13504 11772 13510 11824
rect 14550 11812 14556 11824
rect 14511 11784 14556 11812
rect 14550 11772 14556 11784
rect 14608 11772 14614 11824
rect 15105 11815 15163 11821
rect 15105 11781 15117 11815
rect 15151 11812 15163 11815
rect 15378 11812 15384 11824
rect 15151 11784 15384 11812
rect 15151 11781 15163 11784
rect 15105 11775 15163 11781
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 15749 11815 15807 11821
rect 15749 11781 15761 11815
rect 15795 11812 15807 11815
rect 15795 11784 16712 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 1578 11744 1584 11756
rect 1539 11716 1584 11744
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 6454 11744 6460 11756
rect 5382 11716 6460 11744
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 6730 11744 6736 11756
rect 6691 11716 6736 11744
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 10836 11716 11161 11744
rect 10836 11704 10842 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11882 11744 11888 11756
rect 11296 11716 11888 11744
rect 11296 11704 11302 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2866 11676 2872 11688
rect 1903 11648 2872 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2866 11636 2872 11648
rect 2924 11676 2930 11688
rect 3786 11676 3792 11688
rect 2924 11648 3792 11676
rect 2924 11636 2930 11648
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11676 4307 11679
rect 4890 11676 4896 11688
rect 4295 11648 4896 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 3988 11540 4016 11639
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 6178 11676 6184 11688
rect 5684 11648 6184 11676
rect 5684 11636 5690 11648
rect 6178 11636 6184 11648
rect 6236 11636 6242 11688
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 9122 11676 9128 11688
rect 7055 11648 8984 11676
rect 9083 11648 9128 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 5258 11568 5264 11620
rect 5316 11608 5322 11620
rect 8956 11608 8984 11648
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 11698 11676 11704 11688
rect 9232 11648 11704 11676
rect 9232 11608 9260 11648
rect 11256 11620 11284 11648
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11676 12219 11679
rect 13464 11676 13492 11772
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 13814 11744 13820 11756
rect 13596 11716 13820 11744
rect 13596 11704 13602 11716
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 13906 11676 13912 11688
rect 12207 11648 13492 11676
rect 13867 11648 13912 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 14458 11676 14464 11688
rect 14419 11648 14464 11676
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 16482 11676 16488 11688
rect 15703 11648 16488 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 5316 11580 5948 11608
rect 8956 11580 9260 11608
rect 5316 11568 5322 11580
rect 4062 11540 4068 11552
rect 3975 11512 4068 11540
rect 4062 11500 4068 11512
rect 4120 11540 4126 11552
rect 5810 11540 5816 11552
rect 4120 11512 5816 11540
rect 4120 11500 4126 11512
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 5920 11540 5948 11580
rect 10778 11568 10784 11620
rect 10836 11608 10842 11620
rect 10836 11580 11192 11608
rect 10836 11568 10842 11580
rect 11054 11540 11060 11552
rect 5920 11512 11060 11540
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11164 11540 11192 11580
rect 11238 11568 11244 11620
rect 11296 11568 11302 11620
rect 13262 11568 13268 11620
rect 13320 11608 13326 11620
rect 14550 11608 14556 11620
rect 13320 11580 14556 11608
rect 13320 11568 13326 11580
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 15378 11568 15384 11620
rect 15436 11608 15442 11620
rect 15838 11608 15844 11620
rect 15436 11580 15844 11608
rect 15436 11568 15442 11580
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 16209 11611 16267 11617
rect 16209 11577 16221 11611
rect 16255 11577 16267 11611
rect 16209 11571 16267 11577
rect 14826 11540 14832 11552
rect 11164 11512 14832 11540
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 16224 11540 16252 11571
rect 16482 11540 16488 11552
rect 15160 11512 16488 11540
rect 15160 11500 15166 11512
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16684 11540 16712 11784
rect 16776 11608 16804 11852
rect 16850 11840 16856 11892
rect 16908 11880 16914 11892
rect 16908 11852 16988 11880
rect 16908 11840 16914 11852
rect 16960 11821 16988 11852
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17552 11852 18084 11880
rect 17552 11840 17558 11852
rect 16945 11815 17003 11821
rect 16945 11781 16957 11815
rect 16991 11781 17003 11815
rect 16945 11775 17003 11781
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 17954 11812 17960 11824
rect 17083 11784 17960 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 17586 11636 17592 11688
rect 17644 11676 17650 11688
rect 18056 11676 18084 11852
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18966 11880 18972 11892
rect 18380 11852 18972 11880
rect 18380 11840 18386 11852
rect 18966 11840 18972 11852
rect 19024 11840 19030 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19610 11880 19616 11892
rect 19116 11852 19616 11880
rect 19116 11840 19122 11852
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 20220 11852 20361 11880
rect 20220 11840 20226 11852
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20990 11880 20996 11892
rect 20951 11852 20996 11880
rect 20349 11843 20407 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 24026 11880 24032 11892
rect 21968 11852 24032 11880
rect 21968 11840 21974 11852
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 28813 11883 28871 11889
rect 28813 11880 28825 11883
rect 24320 11852 28825 11880
rect 18509 11815 18567 11821
rect 18509 11812 18521 11815
rect 18340 11784 18521 11812
rect 18340 11756 18368 11784
rect 18509 11781 18521 11784
rect 18555 11781 18567 11815
rect 18509 11775 18567 11781
rect 18601 11815 18659 11821
rect 18601 11781 18613 11815
rect 18647 11812 18659 11815
rect 18647 11784 19288 11812
rect 18647 11781 18659 11784
rect 18601 11775 18659 11781
rect 18322 11704 18328 11756
rect 18380 11704 18386 11756
rect 19260 11744 19288 11784
rect 19334 11772 19340 11824
rect 19392 11812 19398 11824
rect 19705 11815 19763 11821
rect 19705 11812 19717 11815
rect 19392 11784 19717 11812
rect 19392 11772 19398 11784
rect 19705 11781 19717 11784
rect 19751 11781 19763 11815
rect 19705 11775 19763 11781
rect 19794 11772 19800 11824
rect 19852 11812 19858 11824
rect 21082 11812 21088 11824
rect 19852 11784 21088 11812
rect 19852 11772 19858 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 22094 11812 22100 11824
rect 22055 11784 22100 11812
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22925 11815 22983 11821
rect 22925 11812 22937 11815
rect 22336 11784 22937 11812
rect 22336 11772 22342 11784
rect 22925 11781 22937 11784
rect 22971 11781 22983 11815
rect 22925 11775 22983 11781
rect 23474 11772 23480 11824
rect 23532 11812 23538 11824
rect 23934 11812 23940 11824
rect 23532 11784 23940 11812
rect 23532 11772 23538 11784
rect 23934 11772 23940 11784
rect 23992 11772 23998 11824
rect 24320 11821 24348 11852
rect 28813 11849 28825 11852
rect 28859 11849 28871 11883
rect 34054 11880 34060 11892
rect 34015 11852 34060 11880
rect 28813 11843 28871 11849
rect 34054 11840 34060 11852
rect 34112 11840 34118 11892
rect 24305 11815 24363 11821
rect 24305 11812 24317 11815
rect 24044 11784 24317 11812
rect 19518 11744 19524 11756
rect 19260 11716 19524 11744
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 19610 11704 19616 11756
rect 19668 11744 19674 11756
rect 20257 11747 20315 11753
rect 19668 11716 19713 11744
rect 19668 11704 19674 11716
rect 20257 11713 20269 11747
rect 20303 11742 20315 11747
rect 20622 11744 20628 11756
rect 20364 11742 20628 11744
rect 20303 11716 20628 11742
rect 20303 11714 20392 11716
rect 20303 11713 20315 11714
rect 20257 11707 20315 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 20901 11747 20959 11753
rect 20901 11713 20913 11747
rect 20947 11744 20959 11747
rect 21726 11744 21732 11756
rect 20947 11716 21732 11744
rect 20947 11713 20959 11716
rect 20901 11707 20959 11713
rect 21726 11704 21732 11716
rect 21784 11704 21790 11756
rect 21910 11704 21916 11756
rect 21968 11744 21974 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21968 11716 22017 11744
rect 21968 11704 21974 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 24044 11744 24072 11784
rect 24305 11781 24317 11784
rect 24351 11781 24363 11815
rect 24305 11775 24363 11781
rect 24397 11815 24455 11821
rect 24397 11781 24409 11815
rect 24443 11812 24455 11815
rect 25314 11812 25320 11824
rect 24443 11784 25320 11812
rect 24443 11781 24455 11784
rect 24397 11775 24455 11781
rect 25314 11772 25320 11784
rect 25372 11772 25378 11824
rect 25682 11772 25688 11824
rect 25740 11812 25746 11824
rect 25869 11815 25927 11821
rect 25869 11812 25881 11815
rect 25740 11784 25881 11812
rect 25740 11772 25746 11784
rect 25869 11781 25881 11784
rect 25915 11781 25927 11815
rect 25869 11775 25927 11781
rect 25961 11815 26019 11821
rect 25961 11781 25973 11815
rect 26007 11812 26019 11815
rect 27062 11812 27068 11824
rect 26007 11784 27068 11812
rect 26007 11781 26019 11784
rect 25961 11775 26019 11781
rect 27062 11772 27068 11784
rect 27120 11772 27126 11824
rect 34790 11812 34796 11824
rect 31726 11784 34796 11812
rect 22005 11707 22063 11713
rect 23492 11716 24072 11744
rect 18230 11676 18236 11688
rect 17644 11648 17689 11676
rect 18056 11648 18236 11676
rect 17644 11636 17650 11648
rect 18230 11636 18236 11648
rect 18288 11676 18294 11688
rect 18785 11679 18843 11685
rect 18785 11676 18797 11679
rect 18288 11648 18797 11676
rect 18288 11636 18294 11648
rect 18785 11645 18797 11648
rect 18831 11645 18843 11679
rect 22462 11676 22468 11688
rect 18785 11639 18843 11645
rect 18892 11664 19932 11676
rect 20169 11664 22468 11676
rect 18892 11648 22468 11664
rect 18892 11608 18920 11648
rect 19904 11636 20197 11648
rect 22462 11636 22468 11648
rect 22520 11636 22526 11688
rect 22833 11679 22891 11685
rect 22833 11645 22845 11679
rect 22879 11676 22891 11679
rect 22922 11676 22928 11688
rect 22879 11648 22928 11676
rect 22879 11645 22891 11648
rect 22833 11639 22891 11645
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 23106 11676 23112 11688
rect 23067 11648 23112 11676
rect 23106 11636 23112 11648
rect 23164 11636 23170 11688
rect 23492 11676 23520 11716
rect 26694 11704 26700 11756
rect 26752 11744 26758 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26752 11716 27169 11744
rect 26752 11704 26758 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27246 11704 27252 11756
rect 27304 11744 27310 11756
rect 27801 11747 27859 11753
rect 27801 11744 27813 11747
rect 27304 11716 27813 11744
rect 27304 11704 27310 11716
rect 27801 11713 27813 11716
rect 27847 11713 27859 11747
rect 27801 11707 27859 11713
rect 28721 11747 28779 11753
rect 28721 11713 28733 11747
rect 28767 11744 28779 11747
rect 31726 11744 31754 11784
rect 34790 11772 34796 11784
rect 34848 11772 34854 11824
rect 28767 11716 31754 11744
rect 33965 11747 34023 11753
rect 28767 11713 28779 11716
rect 28721 11707 28779 11713
rect 33965 11713 33977 11747
rect 34011 11713 34023 11747
rect 33965 11707 34023 11713
rect 24578 11676 24584 11688
rect 23216 11648 23520 11676
rect 24539 11648 24584 11676
rect 16776 11580 18920 11608
rect 18966 11568 18972 11620
rect 19024 11608 19030 11620
rect 23216 11608 23244 11648
rect 24578 11636 24584 11648
rect 24636 11676 24642 11688
rect 24636 11648 24854 11676
rect 24636 11636 24642 11648
rect 19024 11580 23244 11608
rect 24826 11608 24854 11648
rect 25130 11636 25136 11688
rect 25188 11676 25194 11688
rect 26237 11679 26295 11685
rect 26237 11676 26249 11679
rect 25188 11648 26249 11676
rect 25188 11636 25194 11648
rect 26237 11645 26249 11648
rect 26283 11676 26295 11679
rect 26326 11676 26332 11688
rect 26283 11648 26332 11676
rect 26283 11645 26295 11648
rect 26237 11639 26295 11645
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 31662 11636 31668 11688
rect 31720 11676 31726 11688
rect 33980 11676 34008 11707
rect 37458 11676 37464 11688
rect 31720 11648 34008 11676
rect 37419 11648 37464 11676
rect 31720 11636 31726 11648
rect 37458 11636 37464 11648
rect 37516 11636 37522 11688
rect 37737 11679 37795 11685
rect 37737 11645 37749 11679
rect 37783 11645 37795 11679
rect 37737 11639 37795 11645
rect 26970 11608 26976 11620
rect 24826 11580 26976 11608
rect 19024 11568 19030 11580
rect 26970 11568 26976 11580
rect 27028 11568 27034 11620
rect 27154 11568 27160 11620
rect 27212 11608 27218 11620
rect 27249 11611 27307 11617
rect 27249 11608 27261 11611
rect 27212 11580 27261 11608
rect 27212 11568 27218 11580
rect 27249 11577 27261 11580
rect 27295 11577 27307 11611
rect 27249 11571 27307 11577
rect 28534 11568 28540 11620
rect 28592 11608 28598 11620
rect 37752 11608 37780 11639
rect 28592 11580 37780 11608
rect 28592 11568 28598 11580
rect 18138 11540 18144 11552
rect 16684 11512 18144 11540
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 23750 11540 23756 11552
rect 18472 11512 23756 11540
rect 18472 11500 18478 11512
rect 23750 11500 23756 11512
rect 23808 11500 23814 11552
rect 24026 11500 24032 11552
rect 24084 11540 24090 11552
rect 27893 11543 27951 11549
rect 27893 11540 27905 11543
rect 24084 11512 27905 11540
rect 24084 11500 24090 11512
rect 27893 11509 27905 11512
rect 27939 11509 27951 11543
rect 27893 11503 27951 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 14274 11336 14280 11348
rect 9732 11308 14280 11336
rect 9732 11296 9738 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 15102 11336 15108 11348
rect 14384 11308 15108 11336
rect 3418 11268 3424 11280
rect 3379 11240 3424 11268
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 4065 11271 4123 11277
rect 4065 11237 4077 11271
rect 4111 11268 4123 11271
rect 5258 11268 5264 11280
rect 4111 11240 5264 11268
rect 4111 11237 4123 11240
rect 4065 11231 4123 11237
rect 1578 11160 1584 11212
rect 1636 11200 1642 11212
rect 1673 11203 1731 11209
rect 1673 11200 1685 11203
rect 1636 11172 1685 11200
rect 1636 11160 1642 11172
rect 1673 11169 1685 11172
rect 1719 11169 1731 11203
rect 1673 11163 1731 11169
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 4080 11200 4108 11231
rect 5258 11228 5264 11240
rect 5316 11228 5322 11280
rect 10134 11268 10140 11280
rect 8128 11240 10140 11268
rect 1995 11172 4108 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 5537 11203 5595 11209
rect 4856 11172 5304 11200
rect 4856 11160 4862 11172
rect 5276 11144 5304 11172
rect 5537 11169 5549 11203
rect 5583 11200 5595 11203
rect 5810 11200 5816 11212
rect 5583 11172 5816 11200
rect 5583 11169 5595 11172
rect 5537 11163 5595 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 6822 11200 6828 11212
rect 6328 11172 6828 11200
rect 6328 11160 6334 11172
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7926 11200 7932 11212
rect 7524 11172 7932 11200
rect 7524 11160 7530 11172
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 3970 11092 3976 11144
rect 4028 11132 4034 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4028 11104 4905 11132
rect 4028 11092 4034 11104
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5258 11092 5264 11144
rect 5316 11092 5322 11144
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 8128 11141 8156 11240
rect 10134 11228 10140 11240
rect 10192 11228 10198 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 12526 11268 12532 11280
rect 12308 11240 12532 11268
rect 12308 11228 12314 11240
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 12676 11240 13645 11268
rect 12676 11228 12682 11240
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 13906 11228 13912 11280
rect 13964 11268 13970 11280
rect 14384 11268 14412 11308
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 16298 11336 16304 11348
rect 15344 11308 16304 11336
rect 15344 11296 15350 11308
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 19334 11336 19340 11348
rect 16632 11308 19340 11336
rect 16632 11296 16638 11308
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 19521 11339 19579 11345
rect 19521 11305 19533 11339
rect 19567 11336 19579 11339
rect 19702 11336 19708 11348
rect 19567 11308 19708 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 19702 11296 19708 11308
rect 19760 11296 19766 11348
rect 20898 11336 20904 11348
rect 19904 11308 20904 11336
rect 13964 11240 14412 11268
rect 13964 11228 13970 11240
rect 15746 11228 15752 11280
rect 15804 11268 15810 11280
rect 16758 11268 16764 11280
rect 15804 11240 16764 11268
rect 15804 11228 15810 11240
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 19794 11268 19800 11280
rect 16868 11240 19800 11268
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9861 11203 9919 11209
rect 9861 11200 9873 11203
rect 9180 11172 9873 11200
rect 9180 11160 9186 11172
rect 9861 11169 9873 11172
rect 9907 11200 9919 11203
rect 10873 11203 10931 11209
rect 10873 11200 10885 11203
rect 9907 11172 10885 11200
rect 9907 11169 9919 11172
rect 9861 11163 9919 11169
rect 10873 11169 10885 11172
rect 10919 11169 10931 11203
rect 10873 11163 10931 11169
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 14277 11203 14335 11209
rect 14277 11200 14289 11203
rect 11940 11172 14289 11200
rect 11940 11160 11946 11172
rect 14277 11169 14289 11172
rect 14323 11200 14335 11203
rect 15010 11200 15016 11212
rect 14323 11172 15016 11200
rect 14323 11169 14335 11172
rect 14277 11163 14335 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 15838 11160 15844 11212
rect 15896 11200 15902 11212
rect 16868 11209 16896 11240
rect 19794 11228 19800 11240
rect 19852 11228 19858 11280
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15896 11172 16037 11200
rect 15896 11160 15902 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 16853 11203 16911 11209
rect 16853 11169 16865 11203
rect 16899 11169 16911 11203
rect 16853 11163 16911 11169
rect 17034 11160 17040 11212
rect 17092 11200 17098 11212
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 17092 11172 17141 11200
rect 17092 11160 17098 11172
rect 17129 11169 17141 11172
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 19904 11200 19932 11308
rect 20898 11296 20904 11308
rect 20956 11296 20962 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21729 11339 21787 11345
rect 21729 11336 21741 11339
rect 21232 11308 21741 11336
rect 21232 11296 21238 11308
rect 21729 11305 21741 11308
rect 21775 11305 21787 11339
rect 21729 11299 21787 11305
rect 22186 11296 22192 11348
rect 22244 11336 22250 11348
rect 22373 11339 22431 11345
rect 22373 11336 22385 11339
rect 22244 11308 22385 11336
rect 22244 11296 22250 11308
rect 22373 11305 22385 11308
rect 22419 11305 22431 11339
rect 22373 11299 22431 11305
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25317 11339 25375 11345
rect 25317 11336 25329 11339
rect 24912 11308 25329 11336
rect 24912 11296 24918 11308
rect 25317 11305 25329 11308
rect 25363 11305 25375 11339
rect 25317 11299 25375 11305
rect 25406 11296 25412 11348
rect 25464 11336 25470 11348
rect 25961 11339 26019 11345
rect 25961 11336 25973 11339
rect 25464 11308 25973 11336
rect 25464 11296 25470 11308
rect 25961 11305 25973 11308
rect 26007 11305 26019 11339
rect 26602 11336 26608 11348
rect 26563 11308 26608 11336
rect 25961 11299 26019 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 27062 11296 27068 11348
rect 27120 11336 27126 11348
rect 27249 11339 27307 11345
rect 27249 11336 27261 11339
rect 27120 11308 27261 11336
rect 27120 11296 27126 11308
rect 27249 11305 27261 11308
rect 27295 11305 27307 11339
rect 27249 11299 27307 11305
rect 19978 11228 19984 11280
rect 20036 11268 20042 11280
rect 22554 11268 22560 11280
rect 20036 11240 22560 11268
rect 20036 11228 20042 11240
rect 22554 11228 22560 11240
rect 22612 11268 22618 11280
rect 22612 11240 23428 11268
rect 22612 11228 22618 11240
rect 20622 11200 20628 11212
rect 17368 11172 19932 11200
rect 19989 11172 20628 11200
rect 17368 11160 17374 11172
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11101 8171 11135
rect 9674 11132 9680 11144
rect 8113 11095 8171 11101
rect 9140 11104 9680 11132
rect 4157 11067 4215 11073
rect 3174 11036 4108 11064
rect 4080 10996 4108 11036
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4614 11064 4620 11076
rect 4203 11036 4620 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4614 11024 4620 11036
rect 4672 11064 4678 11076
rect 4798 11064 4804 11076
rect 4672 11036 4804 11064
rect 4672 11024 4678 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 5810 11064 5816 11076
rect 4908 11036 5672 11064
rect 5771 11036 5816 11064
rect 4908 10996 4936 11036
rect 4080 10968 4936 10996
rect 5644 10996 5672 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 7561 11067 7619 11073
rect 7561 11064 7573 11067
rect 7432 11036 7573 11064
rect 7432 11024 7438 11036
rect 7561 11033 7573 11036
rect 7607 11033 7619 11067
rect 8386 11064 8392 11076
rect 8347 11036 8392 11064
rect 7561 11027 7619 11033
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 9140 11073 9168 11104
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12897 11135 12955 11141
rect 12897 11132 12909 11135
rect 12492 11104 12909 11132
rect 12492 11092 12498 11104
rect 12897 11101 12909 11104
rect 12943 11132 12955 11135
rect 13262 11132 13268 11144
rect 12943 11104 13268 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 13814 11132 13820 11144
rect 13587 11104 13820 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 18693 11135 18751 11141
rect 18693 11101 18705 11135
rect 18739 11132 18751 11135
rect 18782 11132 18788 11144
rect 18739 11104 18788 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 19242 11092 19248 11144
rect 19300 11132 19306 11144
rect 19429 11135 19487 11141
rect 19429 11132 19441 11135
rect 19300 11104 19441 11132
rect 19300 11092 19306 11104
rect 19429 11101 19441 11104
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19610 11092 19616 11144
rect 19668 11132 19674 11144
rect 19989 11132 20017 11172
rect 20622 11160 20628 11172
rect 20680 11160 20686 11212
rect 23400 11209 23428 11240
rect 23750 11228 23756 11280
rect 23808 11268 23814 11280
rect 23808 11240 27844 11268
rect 23808 11228 23814 11240
rect 21177 11203 21235 11209
rect 21177 11169 21189 11203
rect 21223 11200 21235 11203
rect 23385 11203 23443 11209
rect 21223 11172 22416 11200
rect 21223 11169 21235 11172
rect 21177 11163 21235 11169
rect 19668 11104 20017 11132
rect 19668 11092 19674 11104
rect 21358 11092 21364 11144
rect 21416 11132 21422 11144
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21416 11104 21649 11132
rect 21416 11092 21422 11104
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 22281 11135 22339 11141
rect 22281 11132 22293 11135
rect 22244 11104 22293 11132
rect 22244 11092 22250 11104
rect 22281 11101 22293 11104
rect 22327 11101 22339 11135
rect 22388 11132 22416 11172
rect 23385 11169 23397 11203
rect 23431 11169 23443 11203
rect 23658 11200 23664 11212
rect 23619 11172 23664 11200
rect 23385 11163 23443 11169
rect 23658 11160 23664 11172
rect 23716 11200 23722 11212
rect 25130 11200 25136 11212
rect 23716 11172 25136 11200
rect 23716 11160 23722 11172
rect 25130 11160 25136 11172
rect 25188 11160 25194 11212
rect 27706 11200 27712 11212
rect 26068 11172 27712 11200
rect 26068 11144 26096 11172
rect 27706 11160 27712 11172
rect 27764 11160 27770 11212
rect 23198 11132 23204 11144
rect 22388 11104 23204 11132
rect 22281 11095 22339 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 24118 11092 24124 11144
rect 24176 11132 24182 11144
rect 24578 11132 24584 11144
rect 24176 11104 24584 11132
rect 24176 11092 24182 11104
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 24762 11132 24768 11144
rect 24723 11104 24768 11132
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 25225 11135 25283 11141
rect 25225 11101 25237 11135
rect 25271 11132 25283 11135
rect 25406 11132 25412 11144
rect 25271 11104 25412 11132
rect 25271 11101 25283 11104
rect 25225 11095 25283 11101
rect 25406 11092 25412 11104
rect 25464 11092 25470 11144
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11132 25927 11135
rect 26050 11132 26056 11144
rect 25915 11104 26056 11132
rect 25915 11101 25927 11104
rect 25869 11095 25927 11101
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 26510 11132 26516 11144
rect 26471 11104 26516 11132
rect 26510 11092 26516 11104
rect 26568 11092 26574 11144
rect 27154 11132 27160 11144
rect 27115 11104 27160 11132
rect 27154 11092 27160 11104
rect 27212 11132 27218 11144
rect 27816 11141 27844 11240
rect 27801 11135 27859 11141
rect 27212 11104 27614 11132
rect 27212 11092 27218 11104
rect 9125 11067 9183 11073
rect 9125 11064 9137 11067
rect 8720 11036 9137 11064
rect 8720 11024 8726 11036
rect 9125 11033 9137 11036
rect 9171 11033 9183 11067
rect 9125 11027 9183 11033
rect 9416 11036 11008 11064
rect 7282 10996 7288 11008
rect 5644 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9416 10996 9444 11036
rect 9364 10968 9444 10996
rect 9364 10956 9370 10968
rect 9490 10956 9496 11008
rect 9548 10996 9554 11008
rect 10410 10996 10416 11008
rect 9548 10968 10416 10996
rect 9548 10956 9554 10968
rect 10410 10956 10416 10968
rect 10468 10956 10474 11008
rect 10980 10996 11008 11036
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11149 11067 11207 11073
rect 11149 11064 11161 11067
rect 11112 11036 11161 11064
rect 11112 11024 11118 11036
rect 11149 11033 11161 11036
rect 11195 11033 11207 11067
rect 12802 11064 12808 11076
rect 12374 11036 12808 11064
rect 11149 11027 11207 11033
rect 12802 11024 12808 11036
rect 12860 11024 12866 11076
rect 13998 11064 14004 11076
rect 13464 11036 14004 11064
rect 13464 10996 13492 11036
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14550 11064 14556 11076
rect 14511 11036 14556 11064
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 14884 11036 15042 11064
rect 14884 11024 14890 11036
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16574 11064 16580 11076
rect 15896 11036 16580 11064
rect 15896 11024 15902 11036
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 16945 11067 17003 11073
rect 16945 11033 16957 11067
rect 16991 11064 17003 11067
rect 17494 11064 17500 11076
rect 16991 11036 17500 11064
rect 16991 11033 17003 11036
rect 16945 11027 17003 11033
rect 17494 11024 17500 11036
rect 17552 11024 17558 11076
rect 18046 11064 18052 11076
rect 18007 11036 18052 11064
rect 18046 11024 18052 11036
rect 18104 11024 18110 11076
rect 18141 11067 18199 11073
rect 18141 11033 18153 11067
rect 18187 11064 18199 11067
rect 18230 11064 18236 11076
rect 18187 11036 18236 11064
rect 18187 11033 18199 11036
rect 18141 11027 18199 11033
rect 18230 11024 18236 11036
rect 18288 11024 18294 11076
rect 18966 11064 18972 11076
rect 18432 11036 18972 11064
rect 10980 10968 13492 10996
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 18432 10996 18460 11036
rect 18966 11024 18972 11036
rect 19024 11024 19030 11076
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 19978 11064 19984 11076
rect 19576 11036 19984 11064
rect 19576 11024 19582 11036
rect 19978 11024 19984 11036
rect 20036 11024 20042 11076
rect 20162 11064 20168 11076
rect 20123 11036 20168 11064
rect 20162 11024 20168 11036
rect 20220 11024 20226 11076
rect 20254 11024 20260 11076
rect 20312 11064 20318 11076
rect 20312 11036 20357 11064
rect 20312 11024 20318 11036
rect 20714 11024 20720 11076
rect 20772 11064 20778 11076
rect 23106 11064 23112 11076
rect 20772 11036 23112 11064
rect 20772 11024 20778 11036
rect 23106 11024 23112 11036
rect 23164 11024 23170 11076
rect 23474 11024 23480 11076
rect 23532 11064 23538 11076
rect 27586 11064 27614 11104
rect 27801 11101 27813 11135
rect 27847 11101 27859 11135
rect 27801 11095 27859 11101
rect 28350 11064 28356 11076
rect 23532 11036 23577 11064
rect 27586 11036 28356 11064
rect 23532 11024 23538 11036
rect 28350 11024 28356 11036
rect 28408 11024 28414 11076
rect 34790 11024 34796 11076
rect 34848 11064 34854 11076
rect 35894 11064 35900 11076
rect 34848 11036 35900 11064
rect 34848 11024 34854 11036
rect 35894 11024 35900 11036
rect 35952 11024 35958 11076
rect 13596 10968 18460 10996
rect 13596 10956 13602 10968
rect 18506 10956 18512 11008
rect 18564 10996 18570 11008
rect 22002 10996 22008 11008
rect 18564 10968 22008 10996
rect 18564 10956 18570 10968
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 24578 10996 24584 11008
rect 24539 10968 24584 10996
rect 24578 10956 24584 10968
rect 24636 10956 24642 11008
rect 24854 10956 24860 11008
rect 24912 10996 24918 11008
rect 25866 10996 25872 11008
rect 24912 10968 25872 10996
rect 24912 10956 24918 10968
rect 25866 10956 25872 10968
rect 25924 10956 25930 11008
rect 27890 10996 27896 11008
rect 27851 10968 27896 10996
rect 27890 10956 27896 10968
rect 27948 10956 27954 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 3970 10792 3976 10804
rect 1636 10764 3976 10792
rect 1636 10752 1642 10764
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 6638 10792 6644 10804
rect 4632 10764 6644 10792
rect 1857 10727 1915 10733
rect 1857 10693 1869 10727
rect 1903 10724 1915 10727
rect 1946 10724 1952 10736
rect 1903 10696 1952 10724
rect 1903 10693 1915 10696
rect 1857 10687 1915 10693
rect 1946 10684 1952 10696
rect 2004 10684 2010 10736
rect 3602 10684 3608 10736
rect 3660 10724 3666 10736
rect 4632 10724 4660 10764
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 13538 10792 13544 10804
rect 6932 10764 13544 10792
rect 6932 10733 6960 10764
rect 13538 10752 13544 10764
rect 13596 10752 13602 10804
rect 17678 10792 17684 10804
rect 14568 10764 17684 10792
rect 3660 10696 4660 10724
rect 5997 10727 6055 10733
rect 3660 10684 3666 10696
rect 5997 10693 6009 10727
rect 6043 10724 6055 10727
rect 6917 10727 6975 10733
rect 6917 10724 6929 10727
rect 6043 10696 6929 10724
rect 6043 10693 6055 10696
rect 5997 10687 6055 10693
rect 6917 10693 6929 10696
rect 6963 10693 6975 10727
rect 9306 10724 9312 10736
rect 6917 10687 6975 10693
rect 8680 10696 9312 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 3970 10656 3976 10668
rect 2990 10628 3740 10656
rect 3931 10628 3976 10656
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3712 10461 3740 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4614 10588 4620 10600
rect 4295 10560 4620 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 5368 10520 5396 10642
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 8294 10616 8300 10668
rect 8352 10656 8358 10668
rect 8680 10665 8708 10696
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9401 10727 9459 10733
rect 9401 10693 9413 10727
rect 9447 10724 9459 10727
rect 9674 10724 9680 10736
rect 9447 10696 9680 10724
rect 9447 10693 9459 10696
rect 9401 10687 9459 10693
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 11698 10724 11704 10736
rect 10626 10696 11704 10724
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 12124 10696 12173 10724
rect 12124 10684 12130 10696
rect 12161 10693 12173 10696
rect 12207 10693 12219 10727
rect 12161 10687 12219 10693
rect 12618 10684 12624 10736
rect 12676 10684 12682 10736
rect 13722 10684 13728 10736
rect 13780 10724 13786 10736
rect 13909 10727 13967 10733
rect 13909 10724 13921 10727
rect 13780 10696 13921 10724
rect 13780 10684 13786 10696
rect 13909 10693 13921 10696
rect 13955 10693 13967 10727
rect 14458 10724 14464 10736
rect 14419 10696 14464 10724
rect 13909 10687 13967 10693
rect 14458 10684 14464 10696
rect 14516 10684 14522 10736
rect 14568 10733 14596 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 17920 10764 18460 10792
rect 17920 10752 17926 10764
rect 14553 10727 14611 10733
rect 14553 10693 14565 10727
rect 14599 10693 14611 10727
rect 14553 10687 14611 10693
rect 15105 10727 15163 10733
rect 15105 10693 15117 10727
rect 15151 10724 15163 10727
rect 15194 10724 15200 10736
rect 15151 10696 15200 10724
rect 15151 10693 15163 10696
rect 15105 10687 15163 10693
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 15470 10684 15476 10736
rect 15528 10724 15534 10736
rect 15657 10727 15715 10733
rect 15657 10724 15669 10727
rect 15528 10696 15669 10724
rect 15528 10684 15534 10696
rect 15657 10693 15669 10696
rect 15703 10693 15715 10727
rect 15657 10687 15715 10693
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10724 15807 10727
rect 15838 10724 15844 10736
rect 15795 10696 15844 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 16298 10724 16304 10736
rect 16259 10696 16304 10724
rect 16298 10684 16304 10696
rect 16356 10684 16362 10736
rect 16942 10724 16948 10736
rect 16903 10696 16948 10724
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 17037 10727 17095 10733
rect 17037 10693 17049 10727
rect 17083 10724 17095 10727
rect 18432 10724 18460 10764
rect 18506 10752 18512 10804
rect 18564 10792 18570 10804
rect 18564 10764 21680 10792
rect 18564 10752 18570 10764
rect 18874 10724 18880 10736
rect 17083 10696 18368 10724
rect 18432 10696 18880 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 18340 10668 18368 10696
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 19153 10727 19211 10733
rect 19153 10693 19165 10727
rect 19199 10724 19211 10727
rect 19242 10724 19248 10736
rect 19199 10696 19248 10724
rect 19199 10693 19211 10696
rect 19153 10687 19211 10693
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 19334 10684 19340 10736
rect 19392 10724 19398 10736
rect 20162 10724 20168 10736
rect 19392 10696 20168 10724
rect 19392 10684 19398 10696
rect 20162 10684 20168 10696
rect 20220 10684 20226 10736
rect 20714 10724 20720 10736
rect 20272 10696 20720 10724
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8352 10628 8677 10656
rect 8352 10616 8358 10628
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10962 10656 10968 10668
rect 10836 10628 10968 10656
rect 10836 10616 10842 10628
rect 10962 10616 10968 10628
rect 11020 10656 11026 10668
rect 11882 10656 11888 10668
rect 11020 10628 11284 10656
rect 11843 10628 11888 10656
rect 11020 10616 11026 10628
rect 6638 10588 6644 10600
rect 6599 10560 6644 10588
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 9122 10588 9128 10600
rect 6748 10560 8984 10588
rect 9083 10560 9128 10588
rect 6748 10520 6776 10560
rect 5368 10492 6776 10520
rect 8956 10520 8984 10560
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 10042 10588 10048 10600
rect 9232 10560 10048 10588
rect 9232 10520 9260 10560
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10557 11207 10591
rect 11256 10588 11284 10628
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18230 10656 18236 10668
rect 18012 10628 18236 10656
rect 18012 10616 18018 10628
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 18322 10616 18328 10668
rect 18380 10616 18386 10668
rect 20272 10656 20300 10696
rect 20714 10684 20720 10696
rect 20772 10684 20778 10736
rect 20901 10727 20959 10733
rect 20901 10693 20913 10727
rect 20947 10724 20959 10727
rect 21542 10724 21548 10736
rect 20947 10696 21548 10724
rect 20947 10693 20959 10696
rect 20901 10687 20959 10693
rect 21542 10684 21548 10696
rect 21600 10684 21606 10736
rect 21652 10724 21680 10764
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 22097 10795 22155 10801
rect 22097 10792 22109 10795
rect 22060 10764 22109 10792
rect 22060 10752 22066 10764
rect 22097 10761 22109 10764
rect 22143 10761 22155 10795
rect 22097 10755 22155 10761
rect 22738 10752 22744 10804
rect 22796 10792 22802 10804
rect 23385 10795 23443 10801
rect 23385 10792 23397 10795
rect 22796 10764 23397 10792
rect 22796 10752 22802 10764
rect 23385 10761 23397 10764
rect 23431 10761 23443 10795
rect 23385 10755 23443 10761
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 24029 10795 24087 10801
rect 24029 10792 24041 10795
rect 23532 10764 24041 10792
rect 23532 10752 23538 10764
rect 24029 10761 24041 10764
rect 24075 10761 24087 10795
rect 26142 10792 26148 10804
rect 24029 10755 24087 10761
rect 24872 10764 25176 10792
rect 26103 10764 26148 10792
rect 24872 10724 24900 10764
rect 25038 10724 25044 10736
rect 21652 10696 24900 10724
rect 24999 10696 25044 10724
rect 19996 10628 20300 10656
rect 19996 10600 20024 10628
rect 20346 10616 20352 10668
rect 20404 10656 20410 10668
rect 20801 10659 20859 10665
rect 20801 10656 20813 10659
rect 20404 10628 20449 10656
rect 20640 10628 20813 10656
rect 20404 10616 20410 10628
rect 20640 10600 20668 10628
rect 20801 10625 20813 10628
rect 20847 10625 20859 10659
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 20801 10619 20859 10625
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22462 10616 22468 10668
rect 22520 10656 22526 10668
rect 22649 10659 22707 10665
rect 22649 10656 22661 10659
rect 22520 10628 22661 10656
rect 22520 10616 22526 10628
rect 22649 10625 22661 10628
rect 22695 10656 22707 10659
rect 22695 10628 22876 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 17218 10588 17224 10600
rect 11256 10560 16813 10588
rect 17179 10560 17224 10588
rect 11149 10551 11207 10557
rect 8956 10492 9260 10520
rect 11164 10520 11192 10551
rect 11698 10520 11704 10532
rect 11164 10492 11704 10520
rect 11698 10480 11704 10492
rect 11756 10520 11762 10532
rect 11882 10520 11888 10532
rect 11756 10492 11888 10520
rect 11756 10480 11762 10492
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 16574 10520 16580 10532
rect 14108 10492 16580 10520
rect 3697 10455 3755 10461
rect 3697 10421 3709 10455
rect 3743 10452 3755 10455
rect 14108 10452 14136 10492
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 16785 10520 16813 10560
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17310 10548 17316 10600
rect 17368 10588 17374 10600
rect 18414 10588 18420 10600
rect 17368 10560 18420 10588
rect 17368 10548 17374 10560
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18506 10548 18512 10600
rect 18564 10548 18570 10600
rect 19058 10588 19064 10600
rect 19019 10560 19064 10588
rect 19058 10548 19064 10560
rect 19116 10548 19122 10600
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 19978 10588 19984 10600
rect 19751 10560 19984 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 20622 10548 20628 10600
rect 20680 10548 20686 10600
rect 20990 10548 20996 10600
rect 21048 10588 21054 10600
rect 22741 10591 22799 10597
rect 22741 10588 22753 10591
rect 21048 10560 22753 10588
rect 21048 10548 21054 10560
rect 22741 10557 22753 10560
rect 22787 10557 22799 10591
rect 22848 10588 22876 10628
rect 23106 10616 23112 10668
rect 23164 10656 23170 10668
rect 23952 10665 23980 10696
rect 25038 10684 25044 10696
rect 25096 10684 25102 10736
rect 25148 10724 25176 10764
rect 26142 10752 26148 10764
rect 26200 10752 26206 10804
rect 28166 10724 28172 10736
rect 25148 10696 28172 10724
rect 28166 10684 28172 10696
rect 28224 10684 28230 10736
rect 38289 10727 38347 10733
rect 38289 10693 38301 10727
rect 38335 10724 38347 10727
rect 38378 10724 38384 10736
rect 38335 10696 38384 10724
rect 38335 10693 38347 10696
rect 38289 10687 38347 10693
rect 38378 10684 38384 10696
rect 38436 10684 38442 10736
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 23164 10628 23305 10656
rect 23164 10616 23170 10628
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 23937 10659 23995 10665
rect 23937 10625 23949 10659
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 25682 10616 25688 10668
rect 25740 10656 25746 10668
rect 26053 10659 26111 10665
rect 26053 10656 26065 10659
rect 25740 10628 26065 10656
rect 25740 10616 25746 10628
rect 26053 10625 26065 10628
rect 26099 10656 26111 10659
rect 26694 10656 26700 10668
rect 26099 10628 26700 10656
rect 26099 10625 26111 10628
rect 26053 10619 26111 10625
rect 26694 10616 26700 10628
rect 26752 10656 26758 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 26752 10628 27169 10656
rect 26752 10616 26758 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 38102 10656 38108 10668
rect 38063 10628 38108 10656
rect 27157 10619 27215 10625
rect 38102 10616 38108 10628
rect 38160 10616 38166 10668
rect 24026 10588 24032 10600
rect 22848 10560 24032 10588
rect 22741 10551 22799 10557
rect 24026 10548 24032 10560
rect 24084 10548 24090 10600
rect 24946 10588 24952 10600
rect 24907 10560 24952 10588
rect 24946 10548 24952 10560
rect 25004 10548 25010 10600
rect 25130 10548 25136 10600
rect 25188 10588 25194 10600
rect 25225 10591 25283 10597
rect 25225 10588 25237 10591
rect 25188 10560 25237 10588
rect 25188 10548 25194 10560
rect 25225 10557 25237 10560
rect 25271 10557 25283 10591
rect 25225 10551 25283 10557
rect 25406 10548 25412 10600
rect 25464 10588 25470 10600
rect 26142 10588 26148 10600
rect 25464 10560 26148 10588
rect 25464 10548 25470 10560
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 18524 10520 18552 10548
rect 25866 10520 25872 10532
rect 16785 10492 18552 10520
rect 19996 10492 25872 10520
rect 3743 10424 14136 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 19996 10452 20024 10492
rect 25866 10480 25872 10492
rect 25924 10520 25930 10532
rect 27154 10520 27160 10532
rect 25924 10492 27160 10520
rect 25924 10480 25930 10492
rect 27154 10480 27160 10492
rect 27212 10480 27218 10532
rect 14240 10424 20024 10452
rect 20165 10455 20223 10461
rect 14240 10412 14246 10424
rect 20165 10421 20177 10455
rect 20211 10452 20223 10455
rect 20346 10452 20352 10464
rect 20211 10424 20352 10452
rect 20211 10421 20223 10424
rect 20165 10415 20223 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 22462 10412 22468 10464
rect 22520 10452 22526 10464
rect 27249 10455 27307 10461
rect 27249 10452 27261 10455
rect 22520 10424 27261 10452
rect 22520 10412 22526 10424
rect 27249 10421 27261 10424
rect 27295 10421 27307 10455
rect 27249 10415 27307 10421
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 2188 10220 3433 10248
rect 2188 10208 2194 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 3421 10211 3479 10217
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 3936 10220 4537 10248
rect 3936 10208 3942 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 7098 10248 7104 10260
rect 4672 10220 7104 10248
rect 4672 10208 4678 10220
rect 7098 10208 7104 10220
rect 7156 10248 7162 10260
rect 14826 10248 14832 10260
rect 7156 10220 14832 10248
rect 7156 10208 7162 10220
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 17218 10248 17224 10260
rect 14976 10220 17224 10248
rect 14976 10208 14982 10220
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 17678 10248 17684 10260
rect 17328 10220 17684 10248
rect 8481 10183 8539 10189
rect 6656 10152 8432 10180
rect 6656 10124 6684 10152
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 1673 10115 1731 10121
rect 1673 10112 1685 10115
rect 1636 10084 1685 10112
rect 1636 10072 1642 10084
rect 1673 10081 1685 10084
rect 1719 10081 1731 10115
rect 1673 10075 1731 10081
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 3234 10112 3240 10124
rect 1995 10084 3240 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 4065 10115 4123 10121
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4614 10112 4620 10124
rect 4111 10084 4620 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4080 10044 4108 10075
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 6638 10112 6644 10124
rect 5123 10084 6644 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 7098 10112 7104 10124
rect 7059 10084 7104 10112
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 8404 10112 8432 10152
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 8754 10180 8760 10192
rect 8527 10152 8760 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 10502 10140 10508 10192
rect 10560 10180 10566 10192
rect 11054 10180 11060 10192
rect 10560 10152 11060 10180
rect 10560 10140 10566 10152
rect 11054 10140 11060 10152
rect 11112 10180 11118 10192
rect 11514 10180 11520 10192
rect 11112 10152 11520 10180
rect 11112 10140 11118 10152
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 13170 10140 13176 10192
rect 13228 10180 13234 10192
rect 13228 10152 13860 10180
rect 13228 10140 13234 10152
rect 9122 10112 9128 10124
rect 8404 10084 9128 10112
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 12434 10112 12440 10124
rect 9447 10084 12440 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 12434 10072 12440 10084
rect 12492 10072 12498 10124
rect 12710 10072 12716 10124
rect 12768 10112 12774 10124
rect 13538 10112 13544 10124
rect 12768 10084 13544 10112
rect 12768 10072 12774 10084
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13832 10112 13860 10152
rect 13906 10140 13912 10192
rect 13964 10180 13970 10192
rect 14182 10180 14188 10192
rect 13964 10152 14188 10180
rect 13964 10140 13970 10152
rect 14182 10140 14188 10152
rect 14240 10140 14246 10192
rect 15654 10140 15660 10192
rect 15712 10180 15718 10192
rect 17328 10180 17356 10220
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 17954 10248 17960 10260
rect 17828 10220 17960 10248
rect 17828 10208 17834 10220
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 20809 10251 20867 10257
rect 20809 10248 20821 10251
rect 18288 10220 20821 10248
rect 18288 10208 18294 10220
rect 20809 10217 20821 10220
rect 20855 10217 20867 10251
rect 20809 10211 20867 10217
rect 21453 10251 21511 10257
rect 21453 10217 21465 10251
rect 21499 10248 21511 10251
rect 21634 10248 21640 10260
rect 21499 10220 21640 10248
rect 21499 10217 21511 10220
rect 21453 10211 21511 10217
rect 21634 10208 21640 10220
rect 21692 10208 21698 10260
rect 22370 10208 22376 10260
rect 22428 10248 22434 10260
rect 22741 10251 22799 10257
rect 22741 10248 22753 10251
rect 22428 10220 22753 10248
rect 22428 10208 22434 10220
rect 22741 10217 22753 10220
rect 22787 10217 22799 10251
rect 22741 10211 22799 10217
rect 23014 10208 23020 10260
rect 23072 10248 23078 10260
rect 24673 10251 24731 10257
rect 24673 10248 24685 10251
rect 23072 10220 24685 10248
rect 23072 10208 23078 10220
rect 24673 10217 24685 10220
rect 24719 10217 24731 10251
rect 25314 10248 25320 10260
rect 25275 10220 25320 10248
rect 24673 10211 24731 10217
rect 25314 10208 25320 10220
rect 25372 10208 25378 10260
rect 30098 10208 30104 10260
rect 30156 10248 30162 10260
rect 32861 10251 32919 10257
rect 32861 10248 32873 10251
rect 30156 10220 32873 10248
rect 30156 10208 30162 10220
rect 32861 10217 32873 10220
rect 32907 10217 32919 10251
rect 32861 10211 32919 10217
rect 15712 10152 17356 10180
rect 15712 10140 15718 10152
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 17460 10152 19012 10180
rect 17460 10140 17466 10152
rect 14826 10112 14832 10124
rect 13832 10084 14832 10112
rect 14826 10072 14832 10084
rect 14884 10072 14890 10124
rect 15473 10115 15531 10121
rect 15473 10081 15485 10115
rect 15519 10112 15531 10115
rect 16298 10112 16304 10124
rect 15519 10084 16304 10112
rect 15519 10081 15531 10084
rect 15473 10075 15531 10081
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 16482 10072 16488 10124
rect 16540 10112 16546 10124
rect 16945 10115 17003 10121
rect 16945 10112 16957 10115
rect 16540 10084 16957 10112
rect 16540 10072 16546 10084
rect 16945 10081 16957 10084
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 18506 10112 18512 10124
rect 17828 10084 18512 10112
rect 17828 10072 17834 10084
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 18984 10112 19012 10152
rect 19058 10140 19064 10192
rect 19116 10180 19122 10192
rect 23198 10180 23204 10192
rect 19116 10152 23204 10180
rect 19116 10140 19122 10152
rect 23198 10140 23204 10152
rect 23256 10140 23262 10192
rect 23934 10180 23940 10192
rect 23895 10152 23940 10180
rect 23934 10140 23940 10152
rect 23992 10140 23998 10192
rect 27798 10140 27804 10192
rect 27856 10140 27862 10192
rect 19150 10112 19156 10124
rect 18984 10084 19156 10112
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 20438 10112 20444 10124
rect 19444 10084 20444 10112
rect 3082 10016 4108 10044
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10013 4399 10047
rect 11514 10044 11520 10056
rect 10534 10016 11520 10044
rect 4341 10007 4399 10013
rect 4356 9908 4384 10007
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11698 10044 11704 10056
rect 11659 10016 11704 10044
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 14458 10044 14464 10056
rect 14419 10016 14464 10044
rect 14458 10004 14464 10016
rect 14516 10044 14522 10056
rect 15286 10044 15292 10056
rect 14516 10016 15292 10044
rect 14516 10004 14522 10016
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 17494 10004 17500 10056
rect 17552 10044 17558 10056
rect 18877 10047 18935 10053
rect 17552 10016 18084 10044
rect 17552 10004 17558 10016
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 5626 9976 5632 9988
rect 5399 9948 5632 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 7466 9976 7472 9988
rect 6578 9948 7472 9976
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 7926 9976 7932 9988
rect 7887 9948 7932 9976
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9976 8079 9979
rect 8110 9976 8116 9988
rect 8067 9948 8116 9976
rect 8067 9945 8079 9948
rect 8021 9939 8079 9945
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 11149 9979 11207 9985
rect 11149 9976 11161 9979
rect 11112 9948 11161 9976
rect 11112 9936 11118 9948
rect 11149 9945 11161 9948
rect 11195 9945 11207 9979
rect 11149 9939 11207 9945
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 11977 9979 12035 9985
rect 11977 9976 11989 9979
rect 11664 9948 11989 9976
rect 11664 9936 11670 9948
rect 11977 9945 11989 9948
rect 12023 9945 12035 9979
rect 11977 9939 12035 9945
rect 12250 9936 12256 9988
rect 12308 9976 12314 9988
rect 13722 9976 13728 9988
rect 12308 9948 12466 9976
rect 13683 9948 13728 9976
rect 12308 9936 12314 9948
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 14366 9936 14372 9988
rect 14424 9976 14430 9988
rect 14737 9979 14795 9985
rect 14737 9976 14749 9979
rect 14424 9948 14749 9976
rect 14424 9936 14430 9948
rect 14737 9945 14749 9948
rect 14783 9976 14795 9979
rect 15194 9976 15200 9988
rect 14783 9948 15200 9976
rect 14783 9945 14795 9948
rect 14737 9939 14795 9945
rect 15194 9936 15200 9948
rect 15252 9936 15258 9988
rect 15565 9979 15623 9985
rect 15565 9945 15577 9979
rect 15611 9976 15623 9979
rect 15930 9976 15936 9988
rect 15611 9948 15936 9976
rect 15611 9945 15623 9948
rect 15565 9939 15623 9945
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 16117 9979 16175 9985
rect 16117 9945 16129 9979
rect 16163 9976 16175 9979
rect 16298 9976 16304 9988
rect 16163 9948 16304 9976
rect 16163 9945 16175 9948
rect 16117 9939 16175 9945
rect 16298 9936 16304 9948
rect 16356 9936 16362 9988
rect 16666 9976 16672 9988
rect 16627 9948 16672 9976
rect 16666 9936 16672 9948
rect 16724 9936 16730 9988
rect 16761 9979 16819 9985
rect 16761 9945 16773 9979
rect 16807 9976 16819 9979
rect 17328 9976 17356 10004
rect 16807 9948 17356 9976
rect 18056 9976 18084 10016
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19444 10044 19472 10084
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 22097 10115 22155 10121
rect 22097 10112 22109 10115
rect 20548 10084 22109 10112
rect 18923 10016 19472 10044
rect 19521 10047 19579 10053
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19521 10013 19533 10047
rect 19567 10044 19579 10047
rect 19567 10016 19840 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 18233 9979 18291 9985
rect 18233 9976 18245 9979
rect 18056 9948 18245 9976
rect 16807 9945 16819 9948
rect 16761 9939 16819 9945
rect 18233 9945 18245 9948
rect 18279 9945 18291 9979
rect 18233 9939 18291 9945
rect 18325 9979 18383 9985
rect 18325 9945 18337 9979
rect 18371 9945 18383 9979
rect 18325 9939 18383 9945
rect 16022 9908 16028 9920
rect 4356 9880 16028 9908
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 16206 9868 16212 9920
rect 16264 9908 16270 9920
rect 17218 9908 17224 9920
rect 16264 9880 17224 9908
rect 16264 9868 16270 9880
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 17402 9868 17408 9920
rect 17460 9908 17466 9920
rect 17954 9908 17960 9920
rect 17460 9880 17960 9908
rect 17460 9868 17466 9880
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18340 9908 18368 9939
rect 18506 9936 18512 9988
rect 18564 9976 18570 9988
rect 19705 9979 19763 9985
rect 19705 9976 19717 9979
rect 18564 9948 19717 9976
rect 18564 9936 18570 9948
rect 19705 9945 19717 9948
rect 19751 9945 19763 9979
rect 19812 9976 19840 10016
rect 19886 10004 19892 10056
rect 19944 10044 19950 10056
rect 20548 10044 20576 10084
rect 22097 10081 22109 10084
rect 22143 10081 22155 10115
rect 22097 10075 22155 10081
rect 22278 10072 22284 10124
rect 22336 10112 22342 10124
rect 27065 10115 27123 10121
rect 22336 10084 24624 10112
rect 22336 10072 22342 10084
rect 19944 10016 20576 10044
rect 20717 10047 20775 10053
rect 19944 10004 19950 10016
rect 20717 10013 20729 10047
rect 20763 10044 20775 10047
rect 20806 10044 20812 10056
rect 20763 10016 20812 10044
rect 20763 10013 20775 10016
rect 20717 10007 20775 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 21082 10004 21088 10056
rect 21140 10044 21146 10056
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 21140 10016 21373 10044
rect 21140 10004 21146 10016
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 22002 10044 22008 10056
rect 21963 10016 22008 10044
rect 21361 10007 21419 10013
rect 22002 10004 22008 10016
rect 22060 10004 22066 10056
rect 22370 10004 22376 10056
rect 22428 10044 22434 10056
rect 24596 10053 24624 10084
rect 27065 10081 27077 10115
rect 27111 10112 27123 10115
rect 27246 10112 27252 10124
rect 27111 10084 27252 10112
rect 27111 10081 27123 10084
rect 27065 10075 27123 10081
rect 27246 10072 27252 10084
rect 27304 10072 27310 10124
rect 27816 10112 27844 10140
rect 27893 10115 27951 10121
rect 27893 10112 27905 10115
rect 27816 10084 27905 10112
rect 27893 10081 27905 10084
rect 27939 10081 27951 10115
rect 27893 10075 27951 10081
rect 22649 10047 22707 10053
rect 22649 10044 22661 10047
rect 22428 10016 22661 10044
rect 22428 10004 22434 10016
rect 22649 10013 22661 10016
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10013 24639 10047
rect 24581 10007 24639 10013
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10044 25283 10047
rect 25498 10044 25504 10056
rect 25271 10016 25504 10044
rect 25271 10013 25283 10016
rect 25225 10007 25283 10013
rect 25498 10004 25504 10016
rect 25556 10004 25562 10056
rect 25866 10044 25872 10056
rect 25827 10016 25872 10044
rect 25866 10004 25872 10016
rect 25924 10004 25930 10056
rect 32769 10047 32827 10053
rect 32769 10013 32781 10047
rect 32815 10044 32827 10047
rect 34422 10044 34428 10056
rect 32815 10016 34428 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 34422 10004 34428 10016
rect 34480 10004 34486 10056
rect 37182 10004 37188 10056
rect 37240 10044 37246 10056
rect 37461 10047 37519 10053
rect 37461 10044 37473 10047
rect 37240 10016 37473 10044
rect 37240 10004 37246 10016
rect 37461 10013 37473 10016
rect 37507 10013 37519 10047
rect 37734 10044 37740 10056
rect 37695 10016 37740 10044
rect 37461 10007 37519 10013
rect 37734 10004 37740 10016
rect 37792 10004 37798 10056
rect 21818 9976 21824 9988
rect 19812 9948 21824 9976
rect 19705 9939 19763 9945
rect 21818 9936 21824 9948
rect 21876 9936 21882 9988
rect 23385 9979 23443 9985
rect 23385 9945 23397 9979
rect 23431 9945 23443 9979
rect 23385 9939 23443 9945
rect 23477 9979 23535 9985
rect 23477 9945 23489 9979
rect 23523 9976 23535 9979
rect 24026 9976 24032 9988
rect 23523 9948 24032 9976
rect 23523 9945 23535 9948
rect 23477 9939 23535 9945
rect 18104 9880 18368 9908
rect 18104 9868 18110 9880
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 21174 9908 21180 9920
rect 19208 9880 21180 9908
rect 19208 9868 19214 9880
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 23400 9908 23428 9939
rect 24026 9936 24032 9948
rect 24084 9936 24090 9988
rect 27157 9979 27215 9985
rect 27157 9945 27169 9979
rect 27203 9976 27215 9979
rect 27890 9976 27896 9988
rect 27203 9948 27896 9976
rect 27203 9945 27215 9948
rect 27157 9939 27215 9945
rect 27890 9936 27896 9948
rect 27948 9936 27954 9988
rect 23348 9880 23428 9908
rect 23348 9868 23354 9880
rect 25406 9868 25412 9920
rect 25464 9908 25470 9920
rect 25961 9911 26019 9917
rect 25961 9908 25973 9911
rect 25464 9880 25973 9908
rect 25464 9868 25470 9880
rect 25961 9877 25973 9880
rect 26007 9877 26019 9911
rect 25961 9871 26019 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 13722 9704 13728 9716
rect 3844 9676 4108 9704
rect 3844 9664 3850 9676
rect 1394 9596 1400 9648
rect 1452 9636 1458 9648
rect 1857 9639 1915 9645
rect 1857 9636 1869 9639
rect 1452 9608 1869 9636
rect 1452 9596 1458 9608
rect 1857 9605 1869 9608
rect 1903 9636 1915 9639
rect 2130 9636 2136 9648
rect 1903 9608 2136 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 3970 9636 3976 9648
rect 3082 9608 3976 9636
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 4080 9636 4108 9676
rect 4724 9676 5672 9704
rect 4724 9636 4752 9676
rect 4080 9608 4752 9636
rect 5644 9636 5672 9676
rect 7208 9676 8156 9704
rect 7208 9636 7236 9676
rect 5644 9608 7236 9636
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 4062 9568 4068 9580
rect 4023 9540 4068 9568
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 6270 9568 6276 9580
rect 5474 9540 6276 9568
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 8128 9568 8156 9676
rect 9692 9676 13728 9704
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 9692 9645 9720 9676
rect 13722 9664 13728 9676
rect 13780 9704 13786 9716
rect 24670 9704 24676 9716
rect 13780 9676 24676 9704
rect 13780 9664 13786 9676
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 25038 9664 25044 9716
rect 25096 9704 25102 9716
rect 26053 9707 26111 9713
rect 26053 9704 26065 9707
rect 25096 9676 26065 9704
rect 25096 9664 25102 9676
rect 26053 9673 26065 9676
rect 26099 9673 26111 9707
rect 26053 9667 26111 9673
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 8536 9608 8861 9636
rect 8536 9596 8542 9608
rect 8849 9605 8861 9608
rect 8895 9605 8907 9639
rect 8849 9599 8907 9605
rect 9677 9639 9735 9645
rect 9677 9605 9689 9639
rect 9723 9636 9735 9639
rect 9723 9608 9757 9636
rect 9723 9605 9735 9608
rect 9677 9599 9735 9605
rect 10410 9596 10416 9648
rect 10468 9596 10474 9648
rect 12250 9596 12256 9648
rect 12308 9636 12314 9648
rect 12308 9608 12650 9636
rect 12308 9596 12314 9608
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13688 9608 13921 9636
rect 13688 9596 13694 9608
rect 13909 9605 13921 9608
rect 13955 9605 13967 9639
rect 14553 9639 14611 9645
rect 14553 9636 14565 9639
rect 13909 9599 13967 9605
rect 14016 9608 14565 9636
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4430 9500 4436 9512
rect 3651 9472 4436 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 4764 9472 5825 9500
rect 4764 9460 4770 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7834 9500 7840 9512
rect 6871 9472 7840 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 2498 9364 2504 9376
rect 2280 9336 2504 9364
rect 2280 9324 2286 9336
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 4328 9367 4386 9373
rect 4328 9333 4340 9367
rect 4374 9364 4386 9367
rect 6086 9364 6092 9376
rect 4374 9336 6092 9364
rect 4374 9333 4386 9336
rect 4328 9327 4386 9333
rect 6086 9324 6092 9336
rect 6144 9324 6150 9376
rect 6564 9364 6592 9463
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 7944 9500 7972 9554
rect 8128 9540 8769 9568
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 9180 9540 9413 9568
rect 9180 9528 9186 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 10134 9500 10140 9512
rect 7944 9472 10140 9500
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10226 9460 10232 9512
rect 10284 9500 10290 9512
rect 10284 9472 11652 9500
rect 10284 9460 10290 9472
rect 9122 9432 9128 9444
rect 8220 9404 9128 9432
rect 8220 9364 8248 9404
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 11624 9432 11652 9472
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11756 9472 11897 9500
rect 11756 9460 11762 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 14016 9500 14044 9608
rect 14553 9605 14565 9608
rect 14599 9605 14611 9639
rect 14553 9599 14611 9605
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 15657 9639 15715 9645
rect 15657 9636 15669 9639
rect 14700 9608 15148 9636
rect 14700 9596 14706 9608
rect 15120 9577 15148 9608
rect 15212 9608 15669 9636
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 11885 9463 11943 9469
rect 11992 9472 14044 9500
rect 14461 9503 14519 9509
rect 11992 9432 12020 9472
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14507 9472 15056 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 10704 9404 11284 9432
rect 11624 9404 12020 9432
rect 6564 9336 8248 9364
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8570 9364 8576 9376
rect 8352 9336 8576 9364
rect 8352 9324 8358 9336
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 10704 9364 10732 9404
rect 11146 9364 11152 9376
rect 8720 9336 10732 9364
rect 11107 9336 11152 9364
rect 8720 9324 8726 9336
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11256 9364 11284 9404
rect 11974 9364 11980 9376
rect 11256 9336 11980 9364
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12148 9367 12206 9373
rect 12148 9333 12160 9367
rect 12194 9364 12206 9367
rect 12342 9364 12348 9376
rect 12194 9336 12348 9364
rect 12194 9333 12206 9336
rect 12148 9327 12206 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 14366 9364 14372 9376
rect 12584 9336 14372 9364
rect 12584 9324 12590 9336
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15028 9364 15056 9472
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 15212 9432 15240 9608
rect 15657 9605 15669 9608
rect 15703 9605 15715 9639
rect 15657 9599 15715 9605
rect 15749 9639 15807 9645
rect 15749 9605 15761 9639
rect 15795 9636 15807 9639
rect 16022 9636 16028 9648
rect 15795 9608 16028 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 16298 9636 16304 9648
rect 16259 9608 16304 9636
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 17394 9639 17452 9645
rect 17394 9636 17406 9639
rect 16816 9608 17406 9636
rect 16816 9596 16822 9608
rect 17394 9605 17406 9608
rect 17440 9605 17452 9639
rect 17394 9599 17452 9605
rect 17490 9639 17548 9645
rect 17490 9605 17502 9639
rect 17536 9636 17548 9639
rect 18230 9636 18236 9648
rect 17536 9608 18236 9636
rect 17536 9605 17548 9608
rect 17490 9599 17548 9605
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 18322 9596 18328 9648
rect 18380 9636 18386 9648
rect 19242 9636 19248 9648
rect 18380 9608 19248 9636
rect 18380 9596 18386 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 19334 9596 19340 9648
rect 19392 9636 19398 9648
rect 19702 9636 19708 9648
rect 19392 9608 19708 9636
rect 19392 9596 19398 9608
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 19812 9608 20660 9636
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16540 9540 16804 9568
rect 16540 9528 16546 9540
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 16022 9500 16028 9512
rect 15712 9472 16028 9500
rect 15712 9460 15718 9472
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 16776 9500 16804 9540
rect 16850 9528 16856 9580
rect 16908 9568 16914 9580
rect 17218 9568 17224 9580
rect 16908 9540 17224 9568
rect 16908 9528 16914 9540
rect 17218 9528 17224 9540
rect 17276 9528 17282 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18064 9540 18521 9568
rect 17681 9503 17739 9509
rect 17681 9500 17693 9503
rect 16776 9472 17693 9500
rect 17681 9469 17693 9472
rect 17727 9469 17739 9503
rect 17681 9463 17739 9469
rect 15160 9404 15240 9432
rect 15160 9392 15166 9404
rect 15286 9392 15292 9444
rect 15344 9432 15350 9444
rect 18064 9432 18092 9540
rect 18509 9537 18521 9540
rect 18555 9568 18567 9571
rect 18800 9568 19012 9574
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 18555 9546 19441 9568
rect 18555 9540 18828 9546
rect 18984 9540 19441 9546
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19812 9568 19840 9608
rect 19429 9531 19487 9537
rect 19628 9540 19840 9568
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18414 9500 18420 9512
rect 18288 9472 18420 9500
rect 18288 9460 18294 9472
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 18656 9472 18705 9500
rect 18656 9460 18662 9472
rect 18693 9469 18705 9472
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19628 9500 19656 9540
rect 18932 9472 19656 9500
rect 18932 9460 18938 9472
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 19760 9472 19805 9500
rect 20548 9488 20576 9608
rect 20632 9577 20660 9608
rect 21174 9596 21180 9648
rect 21232 9636 21238 9648
rect 21361 9639 21419 9645
rect 21232 9608 21312 9636
rect 21232 9596 21238 9608
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 20717 9571 20775 9577
rect 20717 9537 20729 9571
rect 20763 9558 20775 9571
rect 20898 9558 20904 9580
rect 20763 9537 20904 9558
rect 20717 9531 20904 9537
rect 20732 9530 20904 9531
rect 20898 9528 20904 9530
rect 20956 9528 20962 9580
rect 21284 9577 21312 9608
rect 21361 9605 21373 9639
rect 21407 9636 21419 9639
rect 21542 9636 21548 9648
rect 21407 9608 21548 9636
rect 21407 9605 21419 9608
rect 21361 9599 21419 9605
rect 21542 9596 21548 9608
rect 21600 9596 21606 9648
rect 21910 9596 21916 9648
rect 21968 9636 21974 9648
rect 22189 9639 22247 9645
rect 22189 9636 22201 9639
rect 21968 9608 22201 9636
rect 21968 9596 21974 9608
rect 22189 9605 22201 9608
rect 22235 9605 22247 9639
rect 22189 9599 22247 9605
rect 22278 9596 22284 9648
rect 22336 9636 22342 9648
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 22336 9608 22753 9636
rect 22336 9596 22342 9608
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 23845 9639 23903 9645
rect 23845 9605 23857 9639
rect 23891 9636 23903 9639
rect 25406 9636 25412 9648
rect 23891 9608 25412 9636
rect 23891 9605 23903 9608
rect 23845 9599 23903 9605
rect 25406 9596 25412 9608
rect 25464 9596 25470 9648
rect 27893 9639 27951 9645
rect 27893 9605 27905 9639
rect 27939 9636 27951 9639
rect 28718 9636 28724 9648
rect 27939 9608 28724 9636
rect 27939 9605 27951 9608
rect 27893 9599 27951 9605
rect 28718 9596 28724 9608
rect 28776 9596 28782 9648
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 21634 9568 21640 9580
rect 21315 9540 21640 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 24857 9571 24915 9577
rect 24857 9537 24869 9571
rect 24903 9568 24915 9571
rect 25590 9568 25596 9580
rect 24903 9540 25596 9568
rect 24903 9537 24915 9540
rect 24857 9531 24915 9537
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25961 9571 26019 9577
rect 25961 9537 25973 9571
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27801 9571 27859 9577
rect 27801 9537 27813 9571
rect 27847 9568 27859 9571
rect 28810 9568 28816 9580
rect 27847 9540 28816 9568
rect 27847 9537 27859 9540
rect 27801 9531 27859 9537
rect 21542 9500 21548 9512
rect 20686 9488 20852 9500
rect 20916 9488 21548 9500
rect 20548 9472 21548 9488
rect 19760 9460 19766 9472
rect 20548 9460 20714 9472
rect 20824 9460 20944 9472
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9500 22155 9503
rect 23753 9503 23811 9509
rect 23753 9500 23765 9503
rect 22143 9472 23765 9500
rect 22143 9469 22155 9472
rect 22097 9463 22155 9469
rect 23753 9469 23765 9472
rect 23799 9500 23811 9503
rect 24486 9500 24492 9512
rect 23799 9472 24492 9500
rect 23799 9469 23811 9472
rect 23753 9463 23811 9469
rect 24486 9460 24492 9472
rect 24544 9460 24550 9512
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 25976 9500 26004 9531
rect 24728 9472 26004 9500
rect 24728 9460 24734 9472
rect 15344 9404 18092 9432
rect 15344 9392 15350 9404
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 19610 9432 19616 9444
rect 18380 9404 19616 9432
rect 18380 9392 18386 9404
rect 19610 9392 19616 9404
rect 19668 9392 19674 9444
rect 19794 9392 19800 9444
rect 19852 9432 19858 9444
rect 22278 9432 22284 9444
rect 19852 9404 22284 9432
rect 19852 9392 19858 9404
rect 22278 9392 22284 9404
rect 22336 9392 22342 9444
rect 23198 9392 23204 9444
rect 23256 9432 23262 9444
rect 24305 9435 24363 9441
rect 24305 9432 24317 9435
rect 23256 9404 24317 9432
rect 23256 9392 23262 9404
rect 24305 9401 24317 9404
rect 24351 9432 24363 9435
rect 24578 9432 24584 9444
rect 24351 9404 24584 9432
rect 24351 9401 24363 9404
rect 24305 9395 24363 9401
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 25976 9432 26004 9472
rect 26142 9460 26148 9512
rect 26200 9500 26206 9512
rect 27172 9500 27200 9531
rect 28810 9528 28816 9540
rect 28868 9528 28874 9580
rect 29730 9500 29736 9512
rect 26200 9472 27200 9500
rect 27586 9472 29736 9500
rect 26200 9460 26206 9472
rect 27586 9432 27614 9472
rect 29730 9460 29736 9472
rect 29788 9460 29794 9512
rect 25976 9404 27614 9432
rect 20898 9364 20904 9376
rect 15028 9336 20904 9364
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 21542 9324 21548 9376
rect 21600 9364 21606 9376
rect 22186 9364 22192 9376
rect 21600 9336 22192 9364
rect 21600 9324 21606 9336
rect 22186 9324 22192 9336
rect 22244 9324 22250 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 24949 9367 25007 9373
rect 24949 9364 24961 9367
rect 22704 9336 24961 9364
rect 22704 9324 22710 9336
rect 24949 9333 24961 9336
rect 24995 9333 25007 9367
rect 24949 9327 25007 9333
rect 27249 9367 27307 9373
rect 27249 9333 27261 9367
rect 27295 9364 27307 9367
rect 27338 9364 27344 9376
rect 27295 9336 27344 9364
rect 27295 9333 27307 9336
rect 27249 9327 27307 9333
rect 27338 9324 27344 9336
rect 27396 9324 27402 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9120 1676 9172
rect 1728 9160 1734 9172
rect 8294 9160 8300 9172
rect 1728 9132 8300 9160
rect 1728 9120 1734 9132
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 12618 9160 12624 9172
rect 10735 9132 12624 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 13630 9160 13636 9172
rect 12860 9132 13636 9160
rect 12860 9120 12866 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14550 9160 14556 9172
rect 13964 9132 14556 9160
rect 13964 9120 13970 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 15654 9160 15660 9172
rect 14792 9132 15660 9160
rect 14792 9120 14798 9132
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 17144 9132 18460 9160
rect 3050 9052 3056 9104
rect 3108 9092 3114 9104
rect 3329 9095 3387 9101
rect 3329 9092 3341 9095
rect 3108 9064 3341 9092
rect 3108 9052 3114 9064
rect 3329 9061 3341 9064
rect 3375 9092 3387 9095
rect 3694 9092 3700 9104
rect 3375 9064 3700 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 3694 9052 3700 9064
rect 3752 9052 3758 9104
rect 5534 9052 5540 9104
rect 5592 9092 5598 9104
rect 6822 9092 6828 9104
rect 5592 9064 6828 9092
rect 5592 9052 5598 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 8573 9095 8631 9101
rect 8573 9061 8585 9095
rect 8619 9092 8631 9095
rect 10778 9092 10784 9104
rect 8619 9064 10784 9092
rect 8619 9061 8631 9064
rect 8573 9055 8631 9061
rect 10778 9052 10784 9064
rect 10836 9052 10842 9104
rect 17144 9092 17172 9132
rect 17402 9092 17408 9104
rect 10888 9064 11376 9092
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 1596 8996 3985 9024
rect 1596 8968 1624 8996
rect 3973 8993 3985 8996
rect 4019 9024 4031 9027
rect 4246 9024 4252 9036
rect 4019 8996 4252 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 7558 9024 7564 9036
rect 5368 8996 7564 9024
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 5368 8942 5396 8996
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9490 9024 9496 9036
rect 9263 8996 9496 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 9024 9919 9027
rect 10686 9024 10692 9036
rect 9907 8996 10692 9024
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 6822 8956 6828 8968
rect 6783 8928 6828 8956
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 1854 8888 1860 8900
rect 1815 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 3970 8888 3976 8900
rect 3082 8860 3976 8888
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 4154 8848 4160 8900
rect 4212 8888 4218 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 4212 8860 4261 8888
rect 4212 8848 4218 8860
rect 4249 8857 4261 8860
rect 4295 8888 4307 8891
rect 4338 8888 4344 8900
rect 4295 8860 4344 8888
rect 4295 8857 4307 8860
rect 4249 8851 4307 8857
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 5994 8888 6000 8900
rect 5955 8860 6000 8888
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 7101 8891 7159 8897
rect 7101 8857 7113 8891
rect 7147 8857 7159 8891
rect 7101 8851 7159 8857
rect 7116 8820 7144 8851
rect 7558 8848 7564 8900
rect 7616 8848 7622 8900
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 9364 8860 9409 8888
rect 9364 8848 9370 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 10888 8888 10916 9064
rect 11238 9024 11244 9036
rect 11199 8996 11244 9024
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11348 9024 11376 9064
rect 13280 9064 17172 9092
rect 17315 9064 17408 9092
rect 13280 9036 13308 9064
rect 13262 9024 13268 9036
rect 11348 8996 12572 9024
rect 13175 8996 13268 9024
rect 12544 8968 12572 8996
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13906 8984 13912 9036
rect 13964 9024 14228 9036
rect 14292 9024 14504 9036
rect 14734 9024 14740 9036
rect 13964 9008 14740 9024
rect 13964 8984 13970 9008
rect 14200 8996 14320 9008
rect 14476 8996 14740 9008
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 9024 16359 9027
rect 16758 9024 16764 9036
rect 16347 8996 16764 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 16758 8984 16764 8996
rect 16816 9024 16822 9036
rect 17328 9033 17356 9064
rect 17402 9052 17408 9064
rect 17460 9092 17466 9104
rect 18322 9092 18328 9104
rect 17460 9064 18328 9092
rect 17460 9052 17466 9064
rect 18322 9052 18328 9064
rect 18380 9052 18386 9104
rect 18432 9092 18460 9132
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 19521 9163 19579 9169
rect 19521 9160 19533 9163
rect 18748 9132 19533 9160
rect 18748 9120 18754 9132
rect 19521 9129 19533 9132
rect 19567 9129 19579 9163
rect 19521 9123 19579 9129
rect 19610 9120 19616 9172
rect 19668 9160 19674 9172
rect 20622 9160 20628 9172
rect 19668 9132 20628 9160
rect 19668 9120 19674 9132
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 21174 9160 21180 9172
rect 20772 9132 21180 9160
rect 20772 9120 20778 9132
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 21361 9163 21419 9169
rect 21361 9129 21373 9163
rect 21407 9160 21419 9163
rect 21910 9160 21916 9172
rect 21407 9132 21916 9160
rect 21407 9129 21419 9132
rect 21361 9123 21419 9129
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 22186 9120 22192 9172
rect 22244 9160 22250 9172
rect 22244 9132 25544 9160
rect 22244 9120 22250 9132
rect 21542 9092 21548 9104
rect 18432 9064 21548 9092
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 24673 9095 24731 9101
rect 24673 9092 24685 9095
rect 21652 9064 24685 9092
rect 17313 9027 17371 9033
rect 16816 8996 17172 9024
rect 16816 8984 16822 8996
rect 12526 8916 12532 8968
rect 12584 8916 12590 8968
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 15470 8956 15476 8968
rect 13136 8928 15476 8956
rect 13136 8916 13142 8928
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 17144 8956 17172 8996
rect 17313 8993 17325 9027
rect 17359 8993 17371 9027
rect 17586 9024 17592 9036
rect 17313 8987 17371 8993
rect 17420 8996 17592 9024
rect 17420 8956 17448 8996
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 17696 8996 18728 9024
rect 17696 8956 17724 8996
rect 17144 8928 17448 8956
rect 17604 8928 17724 8956
rect 18700 8956 18728 8996
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 18840 8996 18885 9024
rect 18840 8984 18846 8996
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 21652 9024 21680 9064
rect 24673 9061 24685 9064
rect 24719 9061 24731 9095
rect 24673 9055 24731 9061
rect 22833 9027 22891 9033
rect 22833 9024 22845 9027
rect 19024 8996 21680 9024
rect 21744 8996 22845 9024
rect 19024 8984 19030 8996
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18700 8928 19441 8956
rect 11514 8888 11520 8900
rect 9548 8860 10916 8888
rect 11475 8860 11520 8888
rect 9548 8848 9554 8860
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 12066 8848 12072 8900
rect 12124 8848 12130 8900
rect 14265 8891 14323 8897
rect 14265 8857 14277 8891
rect 14311 8888 14323 8891
rect 14366 8888 14372 8900
rect 14311 8860 14372 8888
rect 14311 8857 14323 8860
rect 14265 8851 14323 8857
rect 14366 8848 14372 8860
rect 14424 8848 14430 8900
rect 14734 8848 14740 8900
rect 14792 8888 14798 8900
rect 15105 8891 15163 8897
rect 15105 8888 15117 8891
rect 14792 8860 15117 8888
rect 14792 8848 14798 8860
rect 15105 8857 15117 8860
rect 15151 8857 15163 8891
rect 15105 8851 15163 8857
rect 16393 8891 16451 8897
rect 16393 8857 16405 8891
rect 16439 8857 16451 8891
rect 16393 8851 16451 8857
rect 8110 8820 8116 8832
rect 7116 8792 8116 8820
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 16114 8820 16120 8832
rect 8628 8792 16120 8820
rect 8628 8780 8634 8792
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 16408 8820 16436 8851
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 17604 8888 17632 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 19978 8956 19984 8968
rect 19576 8928 19984 8956
rect 19576 8916 19582 8928
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8956 21327 8959
rect 21358 8956 21364 8968
rect 21315 8928 21364 8956
rect 21315 8925 21327 8928
rect 21269 8919 21327 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 16540 8860 17632 8888
rect 16540 8848 16546 8860
rect 17678 8848 17684 8900
rect 17736 8888 17742 8900
rect 17865 8891 17923 8897
rect 17865 8888 17877 8891
rect 17736 8860 17877 8888
rect 17736 8848 17742 8860
rect 17865 8857 17877 8860
rect 17911 8857 17923 8891
rect 17865 8851 17923 8857
rect 17957 8891 18015 8897
rect 17957 8857 17969 8891
rect 18003 8888 18015 8891
rect 18966 8888 18972 8900
rect 18003 8860 18972 8888
rect 18003 8857 18015 8860
rect 17957 8851 18015 8857
rect 18966 8848 18972 8860
rect 19024 8848 19030 8900
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 19334 8888 19340 8900
rect 19116 8860 19340 8888
rect 19116 8848 19122 8860
rect 19334 8848 19340 8860
rect 19392 8888 19398 8900
rect 20165 8891 20223 8897
rect 20165 8888 20177 8891
rect 19392 8860 20177 8888
rect 19392 8848 19398 8860
rect 20165 8857 20177 8860
rect 20211 8857 20223 8891
rect 20165 8851 20223 8857
rect 20254 8848 20260 8900
rect 20312 8888 20318 8900
rect 20806 8888 20812 8900
rect 20312 8860 20357 8888
rect 20767 8860 20812 8888
rect 20312 8848 20318 8860
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 21744 8888 21772 8996
rect 22833 8993 22845 8996
rect 22879 8993 22891 9027
rect 22833 8987 22891 8993
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 25516 8965 25544 9132
rect 25774 9052 25780 9104
rect 25832 9092 25838 9104
rect 37550 9092 37556 9104
rect 25832 9064 37556 9092
rect 25832 9052 25838 9064
rect 37550 9052 37556 9064
rect 37608 9052 37614 9104
rect 26970 8984 26976 9036
rect 27028 9024 27034 9036
rect 27525 9027 27583 9033
rect 27525 9024 27537 9027
rect 27028 8996 27537 9024
rect 27028 8984 27034 8996
rect 27525 8993 27537 8996
rect 27571 8993 27583 9027
rect 27525 8987 27583 8993
rect 23661 8959 23719 8965
rect 23661 8956 23673 8959
rect 23256 8928 23673 8956
rect 23256 8916 23262 8928
rect 23661 8925 23673 8928
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 25501 8959 25559 8965
rect 25501 8925 25513 8959
rect 25547 8925 25559 8959
rect 38010 8956 38016 8968
rect 37971 8928 38016 8956
rect 25501 8919 25559 8925
rect 22554 8888 22560 8900
rect 21232 8860 21772 8888
rect 22515 8860 22560 8888
rect 21232 8848 21238 8860
rect 22554 8848 22560 8860
rect 22612 8848 22618 8900
rect 22646 8848 22652 8900
rect 22704 8888 22710 8900
rect 24596 8888 24624 8919
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 27246 8888 27252 8900
rect 22704 8860 22749 8888
rect 23584 8860 24624 8888
rect 27207 8860 27252 8888
rect 22704 8848 22710 8860
rect 21358 8820 21364 8832
rect 16408 8792 21364 8820
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 21634 8780 21640 8832
rect 21692 8820 21698 8832
rect 23584 8820 23612 8860
rect 27246 8848 27252 8860
rect 27304 8848 27310 8900
rect 27338 8848 27344 8900
rect 27396 8888 27402 8900
rect 27396 8860 27441 8888
rect 27396 8848 27402 8860
rect 23750 8820 23756 8832
rect 21692 8792 23612 8820
rect 23711 8792 23756 8820
rect 21692 8780 21698 8792
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 25590 8820 25596 8832
rect 25551 8792 25596 8820
rect 25590 8780 25596 8792
rect 25648 8780 25654 8832
rect 25682 8780 25688 8832
rect 25740 8820 25746 8832
rect 27614 8820 27620 8832
rect 25740 8792 27620 8820
rect 25740 8780 25746 8792
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 5997 8619 6055 8625
rect 4172 8588 5948 8616
rect 4172 8548 4200 8588
rect 4614 8548 4620 8560
rect 3082 8520 4200 8548
rect 4264 8520 4620 8548
rect 4264 8492 4292 8520
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5920 8548 5948 8588
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 9214 8616 9220 8628
rect 6043 8588 9220 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 13262 8616 13268 8628
rect 9416 8588 13268 8616
rect 7190 8548 7196 8560
rect 5920 8520 7196 8548
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 8570 8548 8576 8560
rect 8418 8520 8576 8548
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 9416 8557 9444 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14826 8616 14832 8628
rect 14056 8588 14832 8616
rect 14056 8576 14062 8588
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 16482 8616 16488 8628
rect 15396 8588 16488 8616
rect 9401 8551 9459 8557
rect 9401 8517 9413 8551
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 10042 8508 10048 8560
rect 10100 8508 10106 8560
rect 11882 8548 11888 8560
rect 10980 8520 11888 8548
rect 4246 8480 4252 8492
rect 4207 8452 4252 8480
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 9122 8480 9128 8492
rect 9083 8452 9128 8480
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8412 1915 8415
rect 3605 8415 3663 8421
rect 1903 8384 3556 8412
rect 1903 8381 1915 8384
rect 1857 8375 1915 8381
rect 3528 8344 3556 8384
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 4154 8412 4160 8424
rect 3651 8384 4160 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 6914 8412 6920 8424
rect 4571 8384 6776 8412
rect 6875 8384 6920 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 4062 8344 4068 8356
rect 3528 8316 4068 8344
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 6748 8344 6776 8384
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 7193 8415 7251 8421
rect 7193 8381 7205 8415
rect 7239 8412 7251 8415
rect 10980 8412 11008 8520
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 12526 8508 12532 8560
rect 12584 8508 12590 8560
rect 15286 8548 15292 8560
rect 13280 8520 15292 8548
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 13280 8480 13308 8520
rect 15286 8508 15292 8520
rect 15344 8508 15350 8560
rect 15396 8557 15424 8588
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17184 8588 19196 8616
rect 17184 8576 17190 8588
rect 15381 8551 15439 8557
rect 15381 8517 15393 8551
rect 15427 8517 15439 8551
rect 15381 8511 15439 8517
rect 15470 8508 15476 8560
rect 15528 8548 15534 8560
rect 16934 8551 16992 8557
rect 16934 8548 16946 8551
rect 15528 8520 16946 8548
rect 15528 8508 15534 8520
rect 16934 8517 16946 8520
rect 16980 8517 16992 8551
rect 16934 8511 16992 8517
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17310 8548 17316 8560
rect 17083 8520 17316 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 18230 8548 18236 8560
rect 18191 8520 18236 8548
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 18325 8551 18383 8557
rect 18325 8517 18337 8551
rect 18371 8548 18383 8551
rect 18506 8548 18512 8560
rect 18371 8520 18512 8548
rect 18371 8517 18383 8520
rect 18325 8511 18383 8517
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 19168 8548 19196 8588
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 19300 8588 20085 8616
rect 19300 8576 19306 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20073 8579 20131 8585
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 21085 8619 21143 8625
rect 21085 8616 21097 8619
rect 20312 8588 21097 8616
rect 20312 8576 20318 8588
rect 21085 8585 21097 8588
rect 21131 8585 21143 8619
rect 21085 8579 21143 8585
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 21416 8588 25145 8616
rect 21416 8576 21422 8588
rect 25133 8585 25145 8588
rect 25179 8585 25191 8619
rect 28994 8616 29000 8628
rect 28955 8588 29000 8616
rect 25133 8579 25191 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 20346 8548 20352 8560
rect 19168 8520 20352 8548
rect 20346 8508 20352 8520
rect 20404 8508 20410 8560
rect 20456 8520 22048 8548
rect 13188 8452 13308 8480
rect 7239 8384 11008 8412
rect 11149 8415 11207 8421
rect 7239 8381 7251 8384
rect 7193 8375 7251 8381
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 8665 8347 8723 8353
rect 5684 8316 6684 8344
rect 6748 8316 7052 8344
rect 5684 8304 5690 8316
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4982 8276 4988 8288
rect 3936 8248 4988 8276
rect 3936 8236 3942 8248
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 6656 8276 6684 8316
rect 6822 8276 6828 8288
rect 6656 8248 6828 8276
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 7024 8276 7052 8316
rect 8665 8313 8677 8347
rect 8711 8344 8723 8347
rect 8711 8316 9260 8344
rect 8711 8313 8723 8316
rect 8665 8307 8723 8313
rect 7742 8276 7748 8288
rect 7024 8248 7748 8276
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 9232 8276 9260 8316
rect 9858 8276 9864 8288
rect 9232 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10870 8276 10876 8288
rect 10192 8248 10876 8276
rect 10192 8236 10198 8248
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11164 8276 11192 8375
rect 11348 8344 11376 8440
rect 11698 8412 11704 8424
rect 11659 8384 11704 8412
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 11808 8384 11989 8412
rect 11808 8344 11836 8384
rect 11977 8381 11989 8384
rect 12023 8412 12035 8415
rect 13188 8412 13216 8452
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13998 8480 14004 8492
rect 13412 8452 14004 8480
rect 13412 8440 13418 8452
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 14332 8452 14381 8480
rect 14332 8440 14338 8452
rect 14369 8449 14381 8452
rect 14415 8480 14427 8483
rect 14458 8480 14464 8492
rect 14415 8452 14464 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19076 8452 19993 8480
rect 19076 8424 19104 8452
rect 19981 8449 19993 8452
rect 20027 8480 20039 8483
rect 20456 8480 20484 8520
rect 20027 8452 20484 8480
rect 20027 8449 20039 8452
rect 20173 8450 20209 8452
rect 19981 8443 20039 8449
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20864 8452 21005 8480
rect 20864 8440 20870 8452
rect 20993 8449 21005 8452
rect 21039 8480 21051 8483
rect 21910 8480 21916 8492
rect 21039 8452 21916 8480
rect 21039 8449 21051 8452
rect 20993 8443 21051 8449
rect 21910 8440 21916 8452
rect 21968 8440 21974 8492
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 12023 8384 13216 8412
rect 13556 8384 13737 8412
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 11348 8316 11836 8344
rect 12986 8304 12992 8356
rect 13044 8344 13050 8356
rect 13556 8344 13584 8384
rect 13725 8381 13737 8384
rect 13771 8412 13783 8415
rect 15289 8415 15347 8421
rect 13771 8384 15240 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 13044 8316 13584 8344
rect 13044 8304 13050 8316
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 15212 8344 15240 8384
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15838 8412 15844 8424
rect 15335 8384 15844 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8400 16359 8415
rect 16390 8400 16396 8424
rect 16347 8381 16396 8400
rect 16301 8375 16396 8381
rect 16316 8372 16396 8375
rect 16448 8372 16454 8424
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17310 8412 17316 8424
rect 16632 8384 17316 8412
rect 16632 8372 16638 8384
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 17420 8384 17816 8412
rect 17420 8344 17448 8384
rect 13688 8316 14964 8344
rect 15212 8316 17448 8344
rect 17497 8347 17555 8353
rect 13688 8304 13694 8316
rect 14182 8276 14188 8288
rect 11164 8248 14188 8276
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 14645 8279 14703 8285
rect 14645 8245 14657 8279
rect 14691 8276 14703 8279
rect 14826 8276 14832 8288
rect 14691 8248 14832 8276
rect 14691 8245 14703 8248
rect 14645 8239 14703 8245
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 14936 8276 14964 8316
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 17586 8344 17592 8356
rect 17543 8316 17592 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 17586 8304 17592 8316
rect 17644 8304 17650 8356
rect 17788 8344 17816 8384
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18690 8412 18696 8424
rect 17920 8384 18696 8412
rect 17920 8372 17926 8384
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19058 8372 19064 8424
rect 19116 8372 19122 8424
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8412 19303 8415
rect 21542 8412 21548 8424
rect 19291 8384 21548 8412
rect 19291 8381 19303 8384
rect 19245 8375 19303 8381
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 22020 8412 22048 8520
rect 22370 8508 22376 8560
rect 22428 8548 22434 8560
rect 22474 8551 22532 8557
rect 22474 8548 22486 8551
rect 22428 8520 22486 8548
rect 22428 8508 22434 8520
rect 22474 8517 22486 8520
rect 22520 8517 22532 8551
rect 22474 8511 22532 8517
rect 23014 8508 23020 8560
rect 23072 8548 23078 8560
rect 23566 8548 23572 8560
rect 23072 8520 23572 8548
rect 23072 8508 23078 8520
rect 23566 8508 23572 8520
rect 23624 8508 23630 8560
rect 23937 8551 23995 8557
rect 23937 8548 23949 8551
rect 23768 8520 23949 8548
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 23768 8480 23796 8520
rect 23937 8517 23949 8520
rect 23983 8517 23995 8551
rect 23937 8511 23995 8517
rect 23716 8452 23796 8480
rect 23716 8440 23722 8452
rect 23842 8440 23848 8492
rect 23900 8480 23906 8492
rect 24489 8483 24547 8489
rect 23900 8452 23945 8480
rect 23900 8440 23906 8452
rect 24489 8449 24501 8483
rect 24535 8480 24547 8483
rect 24578 8480 24584 8492
rect 24535 8452 24584 8480
rect 24535 8449 24547 8452
rect 24489 8443 24547 8449
rect 24578 8440 24584 8452
rect 24636 8440 24642 8492
rect 25038 8480 25044 8492
rect 24999 8452 25044 8480
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 25498 8480 25504 8492
rect 25459 8452 25504 8480
rect 25498 8440 25504 8452
rect 25556 8480 25562 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 25556 8452 26065 8480
rect 25556 8440 25562 8452
rect 26053 8449 26065 8452
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 28905 8483 28963 8489
rect 28905 8449 28917 8483
rect 28951 8480 28963 8483
rect 29730 8480 29736 8492
rect 28951 8452 29736 8480
rect 28951 8449 28963 8452
rect 28905 8443 28963 8449
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 22373 8415 22431 8421
rect 22020 8384 22324 8412
rect 17788 8316 19748 8344
rect 18506 8276 18512 8288
rect 14936 8248 18512 8276
rect 18506 8236 18512 8248
rect 18564 8236 18570 8288
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 19334 8276 19340 8288
rect 18748 8248 19340 8276
rect 18748 8236 18754 8248
rect 19334 8236 19340 8248
rect 19392 8236 19398 8288
rect 19720 8276 19748 8316
rect 19794 8304 19800 8356
rect 19852 8344 19858 8356
rect 22186 8344 22192 8356
rect 19852 8316 22192 8344
rect 19852 8304 19858 8316
rect 22186 8304 22192 8316
rect 22244 8304 22250 8356
rect 21082 8276 21088 8288
rect 19720 8248 21088 8276
rect 21082 8236 21088 8248
rect 21140 8236 21146 8288
rect 22296 8276 22324 8384
rect 22373 8381 22385 8415
rect 22419 8412 22431 8415
rect 22738 8412 22744 8424
rect 22419 8384 22744 8412
rect 22419 8381 22431 8384
rect 22373 8375 22431 8381
rect 22738 8372 22744 8384
rect 22796 8372 22802 8424
rect 23382 8412 23388 8424
rect 23343 8384 23388 8412
rect 23382 8372 23388 8384
rect 23440 8372 23446 8424
rect 23474 8372 23480 8424
rect 23532 8412 23538 8424
rect 23532 8400 23704 8412
rect 24044 8400 25912 8412
rect 23532 8384 25912 8400
rect 23532 8372 23538 8384
rect 23676 8372 24072 8384
rect 22756 8344 22784 8372
rect 23106 8344 23112 8356
rect 22756 8316 23112 8344
rect 23106 8304 23112 8316
rect 23164 8304 23170 8356
rect 24581 8347 24639 8353
rect 24581 8313 24593 8347
rect 24627 8344 24639 8347
rect 24670 8344 24676 8356
rect 24627 8316 24676 8344
rect 24627 8313 24639 8316
rect 24581 8307 24639 8313
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 25884 8353 25912 8384
rect 25869 8347 25927 8353
rect 25869 8313 25881 8347
rect 25915 8313 25927 8347
rect 25869 8307 25927 8313
rect 23382 8276 23388 8288
rect 22296 8248 23388 8276
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 30834 8276 30840 8288
rect 23624 8248 30840 8276
rect 23624 8236 23630 8248
rect 30834 8236 30840 8248
rect 30892 8236 30898 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 3200 8044 3341 8072
rect 3200 8032 3206 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 3329 8035 3387 8041
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 8662 8072 8668 8084
rect 8527 8044 8668 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 11698 8032 11704 8084
rect 11756 8032 11762 8084
rect 11872 8075 11930 8081
rect 11872 8041 11884 8075
rect 11918 8072 11930 8075
rect 13170 8072 13176 8084
rect 11918 8044 13176 8072
rect 11918 8041 11930 8044
rect 11872 8035 11930 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14366 8072 14372 8084
rect 13780 8044 14372 8072
rect 13780 8032 13786 8044
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 14700 8044 16037 8072
rect 14700 8032 14706 8044
rect 16025 8041 16037 8044
rect 16071 8072 16083 8075
rect 17770 8072 17776 8084
rect 16071 8044 17776 8072
rect 16071 8041 16083 8044
rect 16025 8035 16083 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18472 8044 18828 8072
rect 18472 8032 18478 8044
rect 3694 7964 3700 8016
rect 3752 8004 3758 8016
rect 4982 8004 4988 8016
rect 3752 7976 4988 8004
rect 3752 7964 3758 7976
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 6914 7964 6920 8016
rect 6972 8004 6978 8016
rect 7098 8004 7104 8016
rect 6972 7976 7104 8004
rect 6972 7964 6978 7976
rect 7098 7964 7104 7976
rect 7156 7964 7162 8016
rect 11149 8007 11207 8013
rect 8404 7976 9536 8004
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 3326 7936 3332 7948
rect 1903 7908 3332 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 3326 7896 3332 7908
rect 3384 7936 3390 7948
rect 3878 7936 3884 7948
rect 3384 7908 3884 7936
rect 3384 7896 3390 7908
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 4614 7896 4620 7948
rect 4672 7936 4678 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4672 7908 4721 7936
rect 4672 7896 4678 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 4709 7899 4767 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 7374 7936 7380 7948
rect 6328 7908 7380 7936
rect 6328 7896 6334 7908
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 7742 7936 7748 7948
rect 7607 7908 7748 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7828 1642 7880
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4798 7868 4804 7880
rect 4019 7840 4804 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 8404 7877 8432 7976
rect 9508 7936 9536 7976
rect 11149 7973 11161 8007
rect 11195 8004 11207 8007
rect 11606 8004 11612 8016
rect 11195 7976 11612 8004
rect 11195 7973 11207 7976
rect 11149 7967 11207 7973
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 11330 7936 11336 7948
rect 9508 7908 11336 7936
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 11716 7936 11744 8032
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 16942 8004 16948 8016
rect 12952 7976 13492 8004
rect 12952 7964 12958 7976
rect 13464 7948 13492 7976
rect 15580 7976 16948 8004
rect 11624 7908 11744 7936
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5500 7840 5549 7868
rect 5500 7828 5506 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 11624 7877 11652 7908
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 13188 7936 13400 7948
rect 11940 7920 13400 7936
rect 11940 7908 13216 7920
rect 11940 7896 11946 7908
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9180 7840 9413 7868
rect 9180 7828 9186 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 13372 7868 13400 7920
rect 13446 7896 13452 7948
rect 13504 7936 13510 7948
rect 15580 7936 15608 7976
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 17402 7964 17408 8016
rect 17460 8004 17466 8016
rect 17460 7976 18460 8004
rect 17460 7964 17466 7976
rect 13504 7908 15608 7936
rect 16577 7939 16635 7945
rect 13504 7896 13510 7908
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 16666 7936 16672 7948
rect 16623 7908 16672 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 16850 7896 16856 7948
rect 16908 7936 16914 7948
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 16908 7908 17601 7936
rect 16908 7896 16914 7908
rect 17589 7905 17601 7908
rect 17635 7936 17647 7939
rect 17954 7936 17960 7948
rect 17635 7908 17960 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18432 7945 18460 7976
rect 18506 7964 18512 8016
rect 18564 7964 18570 8016
rect 18800 8004 18828 8044
rect 18874 8032 18880 8084
rect 18932 8072 18938 8084
rect 21453 8075 21511 8081
rect 21453 8072 21465 8075
rect 18932 8044 21465 8072
rect 18932 8032 18938 8044
rect 21453 8041 21465 8044
rect 21499 8041 21511 8075
rect 21453 8035 21511 8041
rect 22462 8032 22468 8084
rect 22520 8072 22526 8084
rect 23385 8075 23443 8081
rect 23385 8072 23397 8075
rect 22520 8044 23397 8072
rect 22520 8032 22526 8044
rect 23385 8041 23397 8044
rect 23431 8041 23443 8075
rect 26234 8072 26240 8084
rect 26195 8044 26240 8072
rect 23385 8035 23443 8041
rect 26234 8032 26240 8044
rect 26292 8032 26298 8084
rect 33962 8032 33968 8084
rect 34020 8072 34026 8084
rect 38105 8075 38163 8081
rect 38105 8072 38117 8075
rect 34020 8044 38117 8072
rect 34020 8032 34026 8044
rect 38105 8041 38117 8044
rect 38151 8041 38163 8075
rect 38105 8035 38163 8041
rect 20254 8004 20260 8016
rect 18800 7976 20260 8004
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 20714 8004 20720 8016
rect 20364 7976 20720 8004
rect 18417 7939 18475 7945
rect 18417 7905 18429 7939
rect 18463 7905 18475 7939
rect 18524 7936 18552 7964
rect 19521 7939 19579 7945
rect 18524 7908 19380 7936
rect 18417 7899 18475 7905
rect 13372 7840 13768 7868
rect 11609 7831 11667 7837
rect 4614 7800 4620 7812
rect 3082 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4816 7800 4844 7828
rect 5718 7800 5724 7812
rect 4816 7772 5724 7800
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 5828 7772 6302 7800
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 5828 7732 5856 7772
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 9732 7772 9777 7800
rect 9732 7760 9738 7772
rect 10134 7760 10140 7812
rect 10192 7760 10198 7812
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 11020 7772 12304 7800
rect 11020 7760 11026 7772
rect 2832 7704 5856 7732
rect 2832 7692 2838 7704
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 8754 7732 8760 7744
rect 6052 7704 8760 7732
rect 6052 7692 6058 7704
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 11882 7732 11888 7744
rect 9272 7704 11888 7732
rect 9272 7692 9278 7704
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12276 7732 12304 7772
rect 12894 7760 12900 7812
rect 12952 7760 12958 7812
rect 13262 7760 13268 7812
rect 13320 7800 13326 7812
rect 13630 7800 13636 7812
rect 13320 7772 13636 7800
rect 13320 7760 13326 7772
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 13740 7800 13768 7840
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13964 7840 14289 7868
rect 13964 7828 13970 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 17552 7840 17993 7868
rect 17552 7828 17558 7840
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 13740 7772 14565 7800
rect 14553 7769 14565 7772
rect 14599 7800 14611 7803
rect 14642 7800 14648 7812
rect 14599 7772 14648 7800
rect 14599 7769 14611 7772
rect 14553 7763 14611 7769
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 15778 7772 16620 7800
rect 13170 7732 13176 7744
rect 12276 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 14734 7732 14740 7744
rect 13872 7704 14740 7732
rect 13872 7692 13878 7704
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14826 7692 14832 7744
rect 14884 7732 14890 7744
rect 16298 7732 16304 7744
rect 14884 7704 16304 7732
rect 14884 7692 14890 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16592 7732 16620 7772
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 17965 7800 17993 7840
rect 19352 7862 19380 7908
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 19886 7936 19892 7948
rect 19567 7908 19892 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20364 7936 20392 7976
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 24210 8004 24216 8016
rect 21376 7976 24216 8004
rect 20180 7908 20392 7936
rect 20441 7939 20499 7945
rect 19429 7871 19487 7877
rect 19429 7862 19441 7871
rect 19352 7837 19441 7862
rect 19475 7837 19487 7871
rect 20180 7868 20208 7908
rect 20441 7905 20453 7939
rect 20487 7936 20499 7939
rect 21174 7936 21180 7948
rect 20487 7908 21180 7936
rect 20487 7905 20499 7908
rect 20441 7899 20499 7905
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 19352 7834 19487 7837
rect 19429 7831 19487 7834
rect 19536 7840 20208 7868
rect 20349 7871 20407 7877
rect 18141 7803 18199 7809
rect 18141 7800 18153 7803
rect 16724 7772 16769 7800
rect 17965 7772 18153 7800
rect 16724 7760 16730 7772
rect 18141 7769 18153 7772
rect 18187 7769 18199 7803
rect 18141 7763 18199 7769
rect 18233 7803 18291 7809
rect 18233 7769 18245 7803
rect 18279 7800 18291 7803
rect 19536 7800 19564 7840
rect 20349 7837 20361 7871
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 18279 7772 19564 7800
rect 18279 7769 18291 7772
rect 18233 7763 18291 7769
rect 17770 7732 17776 7744
rect 16592 7704 17776 7732
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 18156 7732 18184 7763
rect 19610 7760 19616 7812
rect 19668 7800 19674 7812
rect 20364 7800 20392 7831
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21376 7877 21404 7976
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 26418 8004 26424 8016
rect 24320 7976 26424 8004
rect 22741 7939 22799 7945
rect 22741 7936 22753 7939
rect 21744 7908 22753 7936
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 21140 7840 21373 7868
rect 21140 7828 21146 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21542 7828 21548 7880
rect 21600 7868 21606 7880
rect 21744 7868 21772 7908
rect 22741 7905 22753 7908
rect 22787 7905 22799 7939
rect 24320 7936 24348 7976
rect 26418 7964 26424 7976
rect 26476 7964 26482 8016
rect 22741 7899 22799 7905
rect 23400 7908 24348 7936
rect 23400 7880 23428 7908
rect 24670 7896 24676 7948
rect 24728 7936 24734 7948
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24728 7908 24961 7936
rect 24728 7896 24734 7908
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 22002 7868 22008 7880
rect 21600 7840 21772 7868
rect 21963 7840 22008 7868
rect 21600 7828 21606 7840
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 22094 7828 22100 7880
rect 22152 7868 22158 7880
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 22152 7840 22661 7868
rect 22152 7828 22158 7840
rect 22649 7837 22661 7840
rect 22695 7868 22707 7871
rect 23198 7868 23204 7880
rect 22695 7840 23204 7868
rect 22695 7837 22707 7840
rect 22649 7831 22707 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7868 23351 7871
rect 23382 7868 23388 7880
rect 23339 7840 23388 7868
rect 23339 7837 23351 7840
rect 23293 7831 23351 7837
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 26142 7868 26148 7880
rect 26103 7840 26148 7868
rect 26142 7828 26148 7840
rect 26200 7828 26206 7880
rect 38286 7868 38292 7880
rect 38247 7840 38292 7868
rect 38286 7828 38292 7840
rect 38344 7828 38350 7880
rect 19668 7772 20392 7800
rect 19668 7760 19674 7772
rect 21174 7760 21180 7812
rect 21232 7800 21238 7812
rect 23566 7800 23572 7812
rect 21232 7772 23572 7800
rect 21232 7760 21238 7772
rect 23566 7760 23572 7772
rect 23624 7760 23630 7812
rect 24673 7803 24731 7809
rect 24673 7769 24685 7803
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 24765 7803 24823 7809
rect 24765 7769 24777 7803
rect 24811 7800 24823 7803
rect 25590 7800 25596 7812
rect 24811 7772 25596 7800
rect 24811 7769 24823 7772
rect 24765 7763 24823 7769
rect 19978 7732 19984 7744
rect 18156 7704 19984 7732
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20990 7692 20996 7744
rect 21048 7732 21054 7744
rect 22097 7735 22155 7741
rect 22097 7732 22109 7735
rect 21048 7704 22109 7732
rect 21048 7692 21054 7704
rect 22097 7701 22109 7704
rect 22143 7701 22155 7735
rect 24688 7732 24716 7763
rect 25590 7760 25596 7772
rect 25648 7760 25654 7812
rect 24946 7732 24952 7744
rect 24688 7704 24952 7732
rect 22097 7695 22155 7701
rect 24946 7692 24952 7704
rect 25004 7692 25010 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1762 7528 1768 7540
rect 1723 7500 1768 7528
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 5776 7500 10180 7528
rect 5776 7488 5782 7500
rect 4522 7460 4528 7472
rect 3910 7432 4528 7460
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5166 7460 5172 7472
rect 5031 7432 5172 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5166 7420 5172 7432
rect 5224 7420 5230 7472
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 6362 7460 6368 7472
rect 5951 7432 6368 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 6362 7420 6368 7432
rect 6420 7420 6426 7472
rect 6546 7420 6552 7472
rect 6604 7460 6610 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 6604 7432 6837 7460
rect 6604 7420 6610 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 7374 7420 7380 7472
rect 7432 7460 7438 7472
rect 7926 7460 7932 7472
rect 7432 7432 7932 7460
rect 7432 7420 7438 7432
rect 7926 7420 7932 7432
rect 7984 7420 7990 7472
rect 9858 7460 9864 7472
rect 9154 7432 9864 7460
rect 9858 7420 9864 7432
rect 9916 7420 9922 7472
rect 10152 7469 10180 7500
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 12066 7528 12072 7540
rect 10284 7500 12072 7528
rect 10284 7488 10290 7500
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 12176 7500 13860 7528
rect 10137 7463 10195 7469
rect 10137 7429 10149 7463
rect 10183 7429 10195 7463
rect 10137 7423 10195 7429
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 11238 7460 11244 7472
rect 10928 7432 11244 7460
rect 10928 7420 10934 7432
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 11330 7420 11336 7472
rect 11388 7460 11394 7472
rect 12176 7460 12204 7500
rect 13538 7460 13544 7472
rect 11388 7432 12204 7460
rect 13202 7432 13544 7460
rect 11388 7420 11394 7432
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 13832 7460 13860 7500
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15252 7500 16221 7528
rect 15252 7488 15258 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 16209 7491 16267 7497
rect 16482 7488 16488 7540
rect 16540 7528 16546 7540
rect 16850 7528 16856 7540
rect 16540 7500 16856 7528
rect 16540 7488 16546 7500
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 18506 7528 18512 7540
rect 17000 7500 18512 7528
rect 17000 7488 17006 7500
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 18782 7488 18788 7540
rect 18840 7528 18846 7540
rect 22097 7531 22155 7537
rect 22097 7528 22109 7531
rect 18840 7500 22109 7528
rect 18840 7488 18846 7500
rect 22097 7497 22109 7500
rect 22143 7497 22155 7531
rect 22097 7491 22155 7497
rect 23106 7488 23112 7540
rect 23164 7528 23170 7540
rect 23385 7531 23443 7537
rect 23385 7528 23397 7531
rect 23164 7500 23397 7528
rect 23164 7488 23170 7500
rect 23385 7497 23397 7500
rect 23431 7497 23443 7531
rect 24486 7528 24492 7540
rect 24447 7500 24492 7528
rect 23385 7491 23443 7497
rect 24486 7488 24492 7500
rect 24544 7488 24550 7540
rect 24854 7528 24860 7540
rect 24815 7500 24860 7528
rect 24854 7488 24860 7500
rect 24912 7528 24918 7540
rect 25225 7531 25283 7537
rect 25225 7528 25237 7531
rect 24912 7500 25237 7528
rect 24912 7488 24918 7500
rect 25225 7497 25237 7500
rect 25271 7497 25283 7531
rect 25225 7491 25283 7497
rect 37458 7488 37464 7540
rect 37516 7528 37522 7540
rect 38197 7531 38255 7537
rect 38197 7528 38209 7531
rect 37516 7500 38209 7528
rect 37516 7488 37522 7500
rect 38197 7497 38209 7500
rect 38243 7497 38255 7531
rect 38197 7491 38255 7497
rect 17037 7463 17095 7469
rect 13832 7432 14674 7460
rect 17037 7429 17049 7463
rect 17083 7460 17095 7463
rect 17862 7460 17868 7472
rect 17083 7432 17868 7460
rect 17083 7429 17095 7432
rect 17037 7423 17095 7429
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 18138 7420 18144 7472
rect 18196 7460 18202 7472
rect 19521 7463 19579 7469
rect 19521 7460 19533 7463
rect 18196 7432 19533 7460
rect 18196 7420 18202 7432
rect 19521 7429 19533 7432
rect 19567 7429 19579 7463
rect 20806 7460 20812 7472
rect 19521 7423 19579 7429
rect 19621 7432 20812 7460
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 1596 7188 1624 7355
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5813 7395 5871 7401
rect 4856 7364 5672 7392
rect 4856 7352 4862 7364
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 1728 7296 2421 7324
rect 1728 7284 1734 7296
rect 2409 7293 2421 7296
rect 2455 7293 2467 7327
rect 2409 7287 2467 7293
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 3326 7324 3332 7336
rect 2731 7296 3332 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4212 7296 4445 7324
rect 4212 7284 4218 7296
rect 4433 7293 4445 7296
rect 4479 7324 4491 7327
rect 5258 7324 5264 7336
rect 4479 7296 5264 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 5258 7284 5264 7296
rect 5316 7324 5322 7336
rect 5534 7324 5540 7336
rect 5316 7296 5540 7324
rect 5316 7284 5322 7296
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5644 7324 5672 7364
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 5859 7364 6745 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6270 7324 6276 7336
rect 5644 7296 6276 7324
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 5994 7256 6000 7268
rect 4448 7228 6000 7256
rect 4448 7188 4476 7228
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6748 7256 6776 7355
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9677 7395 9735 7401
rect 9272 7364 9628 7392
rect 9272 7352 9278 7364
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7653 7327 7711 7333
rect 7653 7324 7665 7327
rect 7156 7296 7665 7324
rect 7156 7284 7162 7296
rect 7653 7293 7665 7296
rect 7699 7293 7711 7327
rect 9306 7324 9312 7336
rect 7653 7287 7711 7293
rect 7760 7296 9312 7324
rect 7760 7256 7788 7296
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 9600 7324 9628 7364
rect 9677 7361 9689 7395
rect 9723 7392 9735 7395
rect 10502 7392 10508 7404
rect 9723 7364 10508 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 11146 7392 11152 7404
rect 10796 7364 11152 7392
rect 10796 7324 10824 7364
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 13906 7392 13912 7404
rect 13867 7364 13912 7392
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 15838 7392 15844 7404
rect 15528 7364 15844 7392
rect 15528 7352 15534 7364
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 18506 7392 18512 7404
rect 17788 7364 18512 7392
rect 9600 7296 10824 7324
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11701 7327 11759 7333
rect 11701 7324 11713 7327
rect 10919 7296 11713 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11701 7293 11713 7296
rect 11747 7293 11759 7327
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11701 7287 11759 7293
rect 11808 7296 11989 7324
rect 6748 7228 7788 7256
rect 10502 7216 10508 7268
rect 10560 7256 10566 7268
rect 10888 7256 10916 7287
rect 10560 7228 10916 7256
rect 10560 7216 10566 7228
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 11808 7256 11836 7296
rect 11977 7293 11989 7296
rect 12023 7324 12035 7327
rect 14182 7324 14188 7336
rect 12023 7296 14044 7324
rect 14143 7296 14188 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 13446 7256 13452 7268
rect 11664 7228 11836 7256
rect 13407 7228 13452 7256
rect 11664 7216 11670 7228
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 1596 7160 4476 7188
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 11054 7188 11060 7200
rect 4580 7160 11060 7188
rect 4580 7148 4586 7160
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 12342 7188 12348 7200
rect 11848 7160 12348 7188
rect 11848 7148 11854 7160
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 13906 7188 13912 7200
rect 12584 7160 13912 7188
rect 12584 7148 12590 7160
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14016 7188 14044 7296
rect 14182 7284 14188 7296
rect 14240 7324 14246 7336
rect 16945 7327 17003 7333
rect 14240 7296 16896 7324
rect 14240 7284 14246 7296
rect 16868 7256 16896 7296
rect 16945 7293 16957 7327
rect 16991 7324 17003 7327
rect 17034 7324 17040 7336
rect 16991 7296 17040 7324
rect 16991 7293 17003 7296
rect 16945 7287 17003 7293
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 17788 7324 17816 7364
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18656 7364 18797 7392
rect 18656 7352 18662 7364
rect 18785 7361 18797 7364
rect 18831 7361 18843 7395
rect 18785 7355 18843 7361
rect 19058 7352 19064 7404
rect 19116 7392 19122 7404
rect 19429 7395 19487 7401
rect 19429 7392 19441 7395
rect 19116 7364 19441 7392
rect 19116 7352 19122 7364
rect 19429 7361 19441 7364
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 17954 7324 17960 7336
rect 17144 7296 17816 7324
rect 17915 7296 17960 7324
rect 17144 7256 17172 7296
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 18877 7327 18935 7333
rect 18877 7324 18889 7327
rect 18288 7296 18889 7324
rect 18288 7284 18294 7296
rect 18877 7293 18889 7296
rect 18923 7293 18935 7327
rect 18877 7287 18935 7293
rect 18138 7256 18144 7268
rect 15212 7228 16344 7256
rect 16868 7228 17172 7256
rect 17236 7228 18144 7256
rect 15212 7188 15240 7228
rect 14016 7160 15240 7188
rect 15657 7191 15715 7197
rect 15657 7157 15669 7191
rect 15703 7188 15715 7191
rect 16206 7188 16212 7200
rect 15703 7160 16212 7188
rect 15703 7157 15715 7160
rect 15657 7151 15715 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16316 7188 16344 7228
rect 17236 7188 17264 7228
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 19621 7256 19649 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 20901 7463 20959 7469
rect 20901 7429 20913 7463
rect 20947 7460 20959 7463
rect 21542 7460 21548 7472
rect 20947 7432 21548 7460
rect 20947 7429 20959 7432
rect 20901 7423 20959 7429
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 22830 7420 22836 7472
rect 22888 7460 22894 7472
rect 24029 7463 24087 7469
rect 22888 7432 23980 7460
rect 22888 7420 22894 7432
rect 20070 7392 20076 7404
rect 20031 7364 20076 7392
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21692 7364 22017 7392
rect 21692 7352 21698 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7324 20867 7327
rect 22664 7324 22692 7355
rect 23198 7352 23204 7404
rect 23256 7392 23262 7404
rect 23952 7401 23980 7432
rect 24029 7429 24041 7463
rect 24075 7460 24087 7463
rect 25958 7460 25964 7472
rect 24075 7432 25964 7460
rect 24075 7429 24087 7432
rect 24029 7423 24087 7429
rect 25958 7420 25964 7432
rect 26016 7420 26022 7472
rect 23293 7395 23351 7401
rect 23293 7392 23305 7395
rect 23256 7364 23305 7392
rect 23256 7352 23262 7364
rect 23293 7361 23305 7364
rect 23339 7361 23351 7395
rect 23293 7355 23351 7361
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7392 24455 7395
rect 26602 7392 26608 7404
rect 24443 7364 26608 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 26602 7352 26608 7364
rect 26660 7352 26666 7404
rect 38102 7392 38108 7404
rect 38063 7364 38108 7392
rect 38102 7352 38108 7364
rect 38160 7352 38166 7404
rect 24578 7324 24584 7336
rect 20855 7296 22094 7324
rect 22664 7296 24584 7324
rect 20855 7293 20867 7296
rect 20809 7287 20867 7293
rect 20165 7259 20223 7265
rect 20165 7256 20177 7259
rect 18564 7228 19649 7256
rect 19720 7228 20177 7256
rect 18564 7216 18570 7228
rect 16316 7160 17264 7188
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18782 7188 18788 7200
rect 17920 7160 18788 7188
rect 17920 7148 17926 7160
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 18874 7148 18880 7200
rect 18932 7188 18938 7200
rect 19720 7188 19748 7228
rect 20165 7225 20177 7228
rect 20211 7225 20223 7259
rect 20165 7219 20223 7225
rect 20622 7216 20628 7268
rect 20680 7256 20686 7268
rect 21082 7256 21088 7268
rect 20680 7228 21088 7256
rect 20680 7216 20686 7228
rect 21082 7216 21088 7228
rect 21140 7216 21146 7268
rect 21358 7256 21364 7268
rect 21319 7228 21364 7256
rect 21358 7216 21364 7228
rect 21416 7216 21422 7268
rect 22066 7256 22094 7296
rect 24578 7284 24584 7296
rect 24636 7284 24642 7336
rect 24486 7256 24492 7268
rect 22066 7228 24492 7256
rect 24486 7216 24492 7228
rect 24544 7216 24550 7268
rect 18932 7160 19748 7188
rect 18932 7148 18938 7160
rect 19978 7148 19984 7200
rect 20036 7188 20042 7200
rect 22002 7188 22008 7200
rect 20036 7160 22008 7188
rect 20036 7148 20042 7160
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 22738 7188 22744 7200
rect 22699 7160 22744 7188
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1936 6987 1994 6993
rect 1936 6953 1948 6987
rect 1982 6984 1994 6987
rect 3510 6984 3516 6996
rect 1982 6956 3516 6984
rect 1982 6953 1994 6956
rect 1936 6947 1994 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 4614 6944 4620 6996
rect 4672 6984 4678 6996
rect 9030 6984 9036 6996
rect 4672 6956 9036 6984
rect 4672 6944 4678 6956
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9232 6956 11744 6984
rect 6273 6919 6331 6925
rect 6273 6885 6285 6919
rect 6319 6916 6331 6919
rect 6362 6916 6368 6928
rect 6319 6888 6368 6916
rect 6319 6885 6331 6888
rect 6273 6879 6331 6885
rect 6362 6876 6368 6888
rect 6420 6876 6426 6928
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 9122 6916 9128 6928
rect 8168 6888 9128 6916
rect 8168 6876 8174 6888
rect 9122 6876 9128 6888
rect 9180 6876 9186 6928
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1673 6851 1731 6857
rect 1673 6848 1685 6851
rect 1636 6820 1685 6848
rect 1636 6808 1642 6820
rect 1673 6817 1685 6820
rect 1719 6817 1731 6851
rect 1673 6811 1731 6817
rect 3234 6808 3240 6860
rect 3292 6848 3298 6860
rect 3421 6851 3479 6857
rect 3421 6848 3433 6851
rect 3292 6820 3433 6848
rect 3292 6808 3298 6820
rect 3421 6817 3433 6820
rect 3467 6817 3479 6851
rect 4522 6848 4528 6860
rect 4435 6820 4528 6848
rect 3421 6811 3479 6817
rect 4522 6808 4528 6820
rect 4580 6848 4586 6860
rect 5442 6848 5448 6860
rect 4580 6820 5448 6848
rect 4580 6808 4586 6820
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 7098 6848 7104 6860
rect 5500 6820 6316 6848
rect 5500 6808 5506 6820
rect 6288 6792 6316 6820
rect 6748 6820 7104 6848
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 6748 6789 6776 6820
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 6733 6783 6791 6789
rect 6733 6780 6745 6783
rect 6328 6752 6745 6780
rect 6328 6740 6334 6752
rect 6733 6749 6745 6752
rect 6779 6749 6791 6783
rect 9232 6780 9260 6956
rect 11716 6916 11744 6956
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12124 6956 15700 6984
rect 12124 6944 12130 6956
rect 11716 6888 12434 6916
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 12406 6848 12434 6888
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 13262 6916 13268 6928
rect 12676 6888 13268 6916
rect 12676 6876 12682 6888
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 13998 6876 14004 6928
rect 14056 6916 14062 6928
rect 15672 6916 15700 6956
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 17034 6984 17040 6996
rect 15896 6956 17040 6984
rect 15896 6944 15902 6956
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17862 6984 17868 6996
rect 17184 6956 17868 6984
rect 17184 6944 17190 6956
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 17972 6956 18797 6984
rect 17972 6916 18000 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 18785 6947 18843 6953
rect 19058 6944 19064 6996
rect 19116 6984 19122 6996
rect 19116 6956 20024 6984
rect 19116 6944 19122 6956
rect 14056 6888 15608 6916
rect 15672 6888 18000 6916
rect 14056 6876 14062 6888
rect 15580 6860 15608 6888
rect 18138 6876 18144 6928
rect 18196 6916 18202 6928
rect 19996 6916 20024 6956
rect 20070 6944 20076 6996
rect 20128 6984 20134 6996
rect 22738 6984 22744 6996
rect 20128 6956 22744 6984
rect 20128 6944 20134 6956
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 22278 6916 22284 6928
rect 18196 6888 19380 6916
rect 19996 6888 20852 6916
rect 18196 6876 18202 6888
rect 15580 6848 15792 6860
rect 16868 6848 16988 6860
rect 17126 6848 17132 6860
rect 10744 6820 12020 6848
rect 12406 6820 15516 6848
rect 15580 6832 17132 6848
rect 15764 6820 16896 6832
rect 16960 6820 17132 6832
rect 10744 6808 10750 6820
rect 6733 6743 6791 6749
rect 8312 6752 9260 6780
rect 4062 6712 4068 6724
rect 3174 6684 4068 6712
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 4798 6712 4804 6724
rect 4759 6684 4804 6712
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 6638 6712 6644 6724
rect 6026 6684 6644 6712
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 7006 6712 7012 6724
rect 6967 6684 7012 6712
rect 7006 6672 7012 6684
rect 7064 6672 7070 6724
rect 7466 6672 7472 6724
rect 7524 6672 7530 6724
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 4154 6644 4160 6656
rect 1912 6616 4160 6644
rect 1912 6604 1918 6616
rect 4154 6604 4160 6616
rect 4212 6644 4218 6656
rect 8312 6644 8340 6752
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 9364 6752 9597 6780
rect 9364 6740 9370 6752
rect 9585 6749 9597 6752
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10410 6780 10416 6792
rect 9732 6752 9777 6780
rect 10323 6752 10416 6780
rect 9732 6740 9738 6752
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 10428 6712 10456 6740
rect 10686 6712 10692 6724
rect 9180 6684 10456 6712
rect 10647 6684 10692 6712
rect 9180 6672 9186 6684
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 11992 6712 12020 6820
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12802 6780 12808 6792
rect 12483 6752 12808 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12452 6712 12480 6743
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 14274 6780 14280 6792
rect 13311 6752 14280 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14458 6780 14464 6792
rect 14419 6752 14464 6780
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 15102 6780 15108 6792
rect 14608 6752 14653 6780
rect 14752 6752 15108 6780
rect 14608 6740 14614 6752
rect 11072 6684 11178 6712
rect 11992 6684 12480 6712
rect 11072 6656 11100 6684
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 13541 6715 13599 6721
rect 13541 6712 13553 6715
rect 12676 6684 13553 6712
rect 12676 6672 12682 6684
rect 13541 6681 13553 6684
rect 13587 6681 13599 6715
rect 14292 6712 14320 6740
rect 14752 6712 14780 6752
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 14292 6684 14780 6712
rect 15381 6715 15439 6721
rect 13541 6675 13599 6681
rect 15381 6681 15393 6715
rect 15427 6681 15439 6715
rect 15488 6712 15516 6820
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 17494 6848 17500 6860
rect 17455 6820 17500 6848
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 19242 6848 19248 6860
rect 18104 6820 19248 6848
rect 18104 6808 18110 6820
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19352 6848 19380 6888
rect 20162 6848 20168 6860
rect 19352 6820 20024 6848
rect 20123 6820 20168 6848
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 15838 6780 15844 6792
rect 15712 6752 15844 6780
rect 15712 6740 15718 6752
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 16264 6752 16528 6780
rect 16264 6740 16270 6752
rect 16500 6712 16528 6752
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 18693 6783 18751 6789
rect 18693 6780 18705 6783
rect 18656 6752 18705 6780
rect 18656 6740 18662 6752
rect 18693 6749 18705 6752
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 19429 6783 19487 6789
rect 18932 6774 19380 6780
rect 19429 6774 19441 6783
rect 18932 6752 19441 6774
rect 18932 6740 18938 6752
rect 19352 6749 19441 6752
rect 19475 6749 19487 6783
rect 19352 6746 19487 6749
rect 19429 6743 19487 6746
rect 19610 6740 19616 6792
rect 19668 6774 19674 6792
rect 19996 6782 20024 6820
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 20824 6857 20852 6888
rect 22020 6888 22284 6916
rect 20809 6851 20867 6857
rect 20809 6817 20821 6851
rect 20855 6817 20867 6851
rect 20809 6811 20867 6817
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21232 6820 21465 6848
rect 21232 6808 21238 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 20073 6783 20131 6789
rect 20073 6782 20085 6783
rect 19668 6746 19748 6774
rect 19996 6754 20085 6782
rect 19668 6740 19674 6746
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 15488 6684 16436 6712
rect 16500 6684 16681 6712
rect 15381 6675 15439 6681
rect 4212 6616 8340 6644
rect 8481 6647 8539 6653
rect 4212 6604 4218 6616
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 9214 6644 9220 6656
rect 8527 6616 9220 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 10594 6644 10600 6656
rect 10008 6616 10600 6644
rect 10008 6604 10014 6616
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 11054 6604 11060 6656
rect 11112 6604 11118 6656
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 12526 6644 12532 6656
rect 11664 6616 12532 6644
rect 11664 6604 11670 6616
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 14182 6644 14188 6656
rect 12860 6616 14188 6644
rect 12860 6604 12866 6616
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 15396 6644 15424 6675
rect 16114 6644 16120 6656
rect 14332 6616 16120 6644
rect 14332 6604 14338 6616
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16408 6644 16436 6684
rect 16669 6681 16681 6684
rect 16715 6681 16727 6715
rect 16669 6675 16727 6681
rect 16761 6715 16819 6721
rect 16761 6681 16773 6715
rect 16807 6712 16819 6715
rect 19058 6712 19064 6724
rect 16807 6684 19064 6712
rect 16807 6681 16819 6684
rect 16761 6675 16819 6681
rect 19058 6672 19064 6684
rect 19116 6672 19122 6724
rect 19720 6712 19748 6746
rect 20073 6749 20085 6754
rect 20119 6749 20131 6783
rect 20714 6780 20720 6792
rect 20627 6752 20720 6780
rect 20073 6743 20131 6749
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 20990 6740 20996 6792
rect 21048 6780 21054 6792
rect 22020 6789 22048 6888
rect 22278 6876 22284 6888
rect 22336 6876 22342 6928
rect 23382 6848 23388 6860
rect 23343 6820 23388 6848
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 24670 6848 24676 6860
rect 24631 6820 24676 6848
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 27246 6808 27252 6860
rect 27304 6848 27310 6860
rect 27893 6851 27951 6857
rect 27893 6848 27905 6851
rect 27304 6820 27905 6848
rect 27304 6808 27310 6820
rect 27893 6817 27905 6820
rect 27939 6817 27951 6851
rect 27893 6811 27951 6817
rect 31018 6808 31024 6860
rect 31076 6848 31082 6860
rect 33045 6851 33103 6857
rect 33045 6848 33057 6851
rect 31076 6820 33057 6848
rect 31076 6808 31082 6820
rect 33045 6817 33057 6820
rect 33091 6817 33103 6851
rect 33045 6811 33103 6817
rect 21361 6783 21419 6789
rect 21361 6780 21373 6783
rect 21048 6752 21373 6780
rect 21048 6740 21054 6752
rect 21361 6749 21373 6752
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 22005 6783 22063 6789
rect 22005 6749 22017 6783
rect 22051 6749 22063 6783
rect 22005 6743 22063 6749
rect 22094 6740 22100 6792
rect 22152 6780 22158 6792
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 22152 6752 22661 6780
rect 22152 6740 22158 6752
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 23293 6783 23351 6789
rect 23293 6749 23305 6783
rect 23339 6749 23351 6783
rect 23293 6743 23351 6749
rect 20732 6712 20760 6740
rect 19720 6684 20760 6712
rect 20806 6672 20812 6724
rect 20864 6712 20870 6724
rect 23308 6712 23336 6743
rect 23750 6740 23756 6792
rect 23808 6780 23814 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 23808 6752 24593 6780
rect 23808 6740 23814 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 25866 6780 25872 6792
rect 25827 6752 25872 6780
rect 24581 6743 24639 6749
rect 25866 6740 25872 6752
rect 25924 6740 25930 6792
rect 27801 6783 27859 6789
rect 27801 6749 27813 6783
rect 27847 6780 27859 6783
rect 30374 6780 30380 6792
rect 27847 6752 30380 6780
rect 27847 6749 27859 6752
rect 27801 6743 27859 6749
rect 30374 6740 30380 6752
rect 30432 6740 30438 6792
rect 32953 6783 33011 6789
rect 32953 6749 32965 6783
rect 32999 6780 33011 6783
rect 35710 6780 35716 6792
rect 32999 6752 35716 6780
rect 32999 6749 33011 6752
rect 32953 6743 33011 6749
rect 35710 6740 35716 6752
rect 35768 6740 35774 6792
rect 20864 6684 23336 6712
rect 20864 6672 20870 6684
rect 19426 6644 19432 6656
rect 16408 6616 19432 6644
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 19521 6647 19579 6653
rect 19521 6613 19533 6647
rect 19567 6644 19579 6647
rect 20530 6644 20536 6656
rect 19567 6616 20536 6644
rect 19567 6613 19579 6616
rect 19521 6607 19579 6613
rect 20530 6604 20536 6616
rect 20588 6604 20594 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22738 6644 22744 6656
rect 22152 6616 22197 6644
rect 22699 6616 22744 6644
rect 22152 6604 22158 6616
rect 22738 6604 22744 6616
rect 22796 6604 22802 6656
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 23348 6616 25973 6644
rect 23348 6604 23354 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 4522 6440 4528 6452
rect 2056 6412 4528 6440
rect 2056 6313 2084 6412
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 7466 6440 7472 6452
rect 5951 6412 7472 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 8260 6412 9873 6440
rect 8260 6400 8266 6412
rect 9861 6409 9873 6412
rect 9907 6440 9919 6443
rect 10042 6440 10048 6452
rect 9907 6412 10048 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10336 6412 10640 6440
rect 2314 6372 2320 6384
rect 2275 6344 2320 6372
rect 2314 6332 2320 6344
rect 2372 6332 2378 6384
rect 4065 6375 4123 6381
rect 4065 6341 4077 6375
rect 4111 6372 4123 6375
rect 4154 6372 4160 6384
rect 4111 6344 4160 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 5718 6332 5724 6384
rect 5776 6372 5782 6384
rect 6549 6375 6607 6381
rect 6549 6372 6561 6375
rect 5776 6344 6561 6372
rect 5776 6332 5782 6344
rect 6549 6341 6561 6344
rect 6595 6341 6607 6375
rect 6549 6335 6607 6341
rect 7098 6332 7104 6384
rect 7156 6372 7162 6384
rect 7285 6375 7343 6381
rect 7285 6372 7297 6375
rect 7156 6344 7297 6372
rect 7156 6332 7162 6344
rect 7285 6341 7297 6344
rect 7331 6341 7343 6375
rect 8662 6372 8668 6384
rect 7285 6335 7343 6341
rect 7944 6344 8668 6372
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 3970 6304 3976 6316
rect 3450 6276 3976 6304
rect 2041 6267 2099 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 7944 6304 7972 6344
rect 8662 6332 8668 6344
rect 8720 6332 8726 6384
rect 9674 6332 9680 6384
rect 9732 6372 9738 6384
rect 10336 6372 10364 6412
rect 9732 6344 10364 6372
rect 10612 6372 10640 6412
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 10744 6412 10789 6440
rect 10744 6400 10750 6412
rect 10870 6400 10876 6452
rect 10928 6440 10934 6452
rect 10928 6412 11192 6440
rect 10928 6400 10934 6412
rect 10962 6372 10968 6384
rect 10612 6344 10968 6372
rect 9732 6332 9738 6344
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 11164 6372 11192 6412
rect 11532 6412 11836 6440
rect 11532 6372 11560 6412
rect 11164 6344 11560 6372
rect 11808 6372 11836 6412
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 18874 6440 18880 6452
rect 12216 6412 18880 6440
rect 12216 6400 12222 6412
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 19702 6440 19708 6452
rect 19300 6412 19708 6440
rect 19300 6400 19306 6412
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 21174 6440 21180 6452
rect 19812 6412 21180 6440
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11808 6344 11989 6372
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 13722 6372 13728 6384
rect 13202 6344 13728 6372
rect 11977 6335 12035 6341
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 14182 6372 14188 6384
rect 14143 6344 14188 6372
rect 14182 6332 14188 6344
rect 14240 6332 14246 6384
rect 15105 6375 15163 6381
rect 15105 6341 15117 6375
rect 15151 6372 15163 6375
rect 15378 6372 15384 6384
rect 15151 6344 15384 6372
rect 15151 6341 15163 6344
rect 15105 6335 15163 6341
rect 15378 6332 15384 6344
rect 15436 6332 15442 6384
rect 16574 6332 16580 6384
rect 16632 6372 16638 6384
rect 17037 6375 17095 6381
rect 17037 6372 17049 6375
rect 16632 6344 17049 6372
rect 16632 6332 16638 6344
rect 17037 6341 17049 6344
rect 17083 6341 17095 6375
rect 17037 6335 17095 6341
rect 17126 6332 17132 6384
rect 17184 6372 17190 6384
rect 19812 6372 19840 6412
rect 21174 6400 21180 6412
rect 21232 6400 21238 6452
rect 22278 6440 22284 6452
rect 22239 6412 22284 6440
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 23566 6440 23572 6452
rect 23527 6412 23572 6440
rect 23566 6400 23572 6412
rect 23624 6400 23630 6452
rect 23937 6443 23995 6449
rect 23937 6409 23949 6443
rect 23983 6440 23995 6443
rect 24394 6440 24400 6452
rect 23983 6412 24400 6440
rect 23983 6409 23995 6412
rect 23937 6403 23995 6409
rect 24394 6400 24400 6412
rect 24452 6400 24458 6452
rect 20070 6372 20076 6384
rect 17184 6344 19840 6372
rect 20031 6344 20076 6372
rect 17184 6332 17190 6344
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 20162 6332 20168 6384
rect 20220 6372 20226 6384
rect 20714 6372 20720 6384
rect 20220 6344 20720 6372
rect 20220 6332 20226 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 20898 6332 20904 6384
rect 20956 6372 20962 6384
rect 21913 6375 21971 6381
rect 21913 6372 21925 6375
rect 20956 6344 21925 6372
rect 20956 6332 20962 6344
rect 21913 6341 21925 6344
rect 21959 6341 21971 6375
rect 21913 6335 21971 6341
rect 8110 6304 8116 6316
rect 5859 6276 7972 6304
rect 8071 6276 8116 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 4540 6236 4568 6267
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 9490 6264 9496 6316
rect 9548 6264 9554 6316
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 10560 6276 10609 6304
rect 10560 6264 10566 6276
rect 10597 6273 10609 6276
rect 10643 6273 10655 6307
rect 10597 6267 10655 6273
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11664 6276 11713 6304
rect 11664 6264 11670 6276
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 15657 6307 15715 6313
rect 15657 6273 15669 6307
rect 15703 6304 15715 6307
rect 16482 6304 16488 6316
rect 15703 6276 16488 6304
rect 15703 6273 15715 6276
rect 15657 6267 15715 6273
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 17644 6276 17689 6304
rect 17644 6264 17650 6276
rect 17770 6264 17776 6316
rect 17828 6304 17834 6316
rect 18138 6304 18144 6316
rect 17828 6276 18144 6304
rect 17828 6264 17834 6276
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18417 6307 18475 6313
rect 18417 6273 18429 6307
rect 18463 6304 18475 6307
rect 18598 6304 18604 6316
rect 18463 6276 18604 6304
rect 18463 6273 18475 6276
rect 18417 6267 18475 6273
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 19058 6264 19064 6316
rect 19116 6304 19122 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 19116 6276 19349 6304
rect 19116 6264 19122 6276
rect 19337 6273 19349 6276
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6304 19487 6307
rect 19610 6304 19616 6316
rect 19475 6276 19616 6304
rect 19475 6273 19487 6276
rect 19429 6267 19487 6273
rect 19610 6264 19616 6276
rect 19668 6264 19674 6316
rect 19978 6304 19984 6316
rect 19939 6276 19984 6304
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20254 6304 20260 6316
rect 20180 6276 20260 6304
rect 8389 6239 8447 6245
rect 4540 6208 8248 6236
rect 3694 6128 3700 6180
rect 3752 6168 3758 6180
rect 4709 6171 4767 6177
rect 4709 6168 4721 6171
rect 3752 6140 4721 6168
rect 3752 6128 3758 6140
rect 4709 6137 4721 6140
rect 4755 6137 4767 6171
rect 4709 6131 4767 6137
rect 4982 6128 4988 6180
rect 5040 6168 5046 6180
rect 5442 6168 5448 6180
rect 5040 6140 5448 6168
rect 5040 6128 5046 6140
rect 5442 6128 5448 6140
rect 5500 6168 5506 6180
rect 8110 6168 8116 6180
rect 5500 6140 8116 6168
rect 5500 6128 5506 6140
rect 8110 6128 8116 6140
rect 8168 6128 8174 6180
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 7834 6100 7840 6112
rect 3476 6072 7840 6100
rect 3476 6060 3482 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8220 6100 8248 6208
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 10686 6236 10692 6248
rect 8435 6208 10692 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 10870 6196 10876 6248
rect 10928 6236 10934 6248
rect 10928 6208 13216 6236
rect 10928 6196 10934 6208
rect 10962 6128 10968 6180
rect 11020 6168 11026 6180
rect 13188 6168 13216 6208
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13320 6208 14105 6236
rect 13320 6196 13326 6208
rect 14093 6205 14105 6208
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15160 6208 15853 6236
rect 15160 6196 15166 6208
rect 15841 6205 15853 6208
rect 15887 6205 15899 6239
rect 16942 6236 16948 6248
rect 16903 6208 16948 6236
rect 15841 6199 15899 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 20180 6236 20208 6276
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20496 6276 20637 6304
rect 20496 6264 20502 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 21174 6264 21180 6316
rect 21232 6304 21238 6316
rect 21269 6307 21327 6313
rect 21269 6304 21281 6307
rect 21232 6276 21281 6304
rect 21232 6264 21238 6276
rect 21269 6273 21281 6276
rect 21315 6273 21327 6307
rect 21818 6304 21824 6316
rect 21779 6276 21824 6304
rect 21269 6267 21327 6273
rect 21818 6264 21824 6276
rect 21876 6264 21882 6316
rect 22296 6304 22324 6400
rect 22462 6332 22468 6384
rect 22520 6372 22526 6384
rect 22520 6344 23428 6372
rect 22520 6332 22526 6344
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 22296 6276 22845 6304
rect 22833 6273 22845 6276
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6273 23351 6307
rect 23293 6267 23351 6273
rect 20717 6239 20775 6245
rect 17045 6208 20208 6236
rect 20272 6208 20484 6236
rect 13449 6171 13507 6177
rect 13449 6168 13461 6171
rect 11020 6140 11192 6168
rect 13188 6140 13461 6168
rect 11020 6128 11026 6140
rect 9674 6100 9680 6112
rect 8220 6072 9680 6100
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 11164 6100 11192 6140
rect 13449 6137 13461 6140
rect 13495 6168 13507 6171
rect 17045 6168 17073 6208
rect 20272 6168 20300 6208
rect 13495 6140 17073 6168
rect 17144 6140 20300 6168
rect 20456 6168 20484 6208
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 22554 6236 22560 6248
rect 20763 6208 22560 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 20990 6168 20996 6180
rect 20456 6140 20996 6168
rect 13495 6137 13507 6140
rect 13449 6131 13507 6137
rect 14642 6100 14648 6112
rect 11164 6072 14648 6100
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 17144 6100 17172 6140
rect 20990 6128 20996 6140
rect 21048 6128 21054 6180
rect 21358 6168 21364 6180
rect 21319 6140 21364 6168
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 23308 6168 23336 6267
rect 23400 6236 23428 6344
rect 23584 6304 23612 6400
rect 24121 6307 24179 6313
rect 24121 6304 24133 6307
rect 23584 6276 24133 6304
rect 24121 6273 24133 6276
rect 24167 6273 24179 6307
rect 24121 6267 24179 6273
rect 32309 6307 32367 6313
rect 32309 6273 32321 6307
rect 32355 6304 32367 6307
rect 35802 6304 35808 6316
rect 32355 6276 35808 6304
rect 32355 6273 32367 6276
rect 32309 6267 32367 6273
rect 35802 6264 35808 6276
rect 35860 6264 35866 6316
rect 23400 6208 31754 6236
rect 21836 6140 23336 6168
rect 31726 6168 31754 6208
rect 38010 6168 38016 6180
rect 31726 6140 38016 6168
rect 16908 6072 17172 6100
rect 16908 6060 16914 6072
rect 17494 6060 17500 6112
rect 17552 6100 17558 6112
rect 18509 6103 18567 6109
rect 18509 6100 18521 6103
rect 17552 6072 18521 6100
rect 17552 6060 17558 6072
rect 18509 6069 18521 6072
rect 18555 6069 18567 6103
rect 18509 6063 18567 6069
rect 19242 6060 19248 6112
rect 19300 6100 19306 6112
rect 20162 6100 20168 6112
rect 19300 6072 20168 6100
rect 19300 6060 19306 6072
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 20438 6060 20444 6112
rect 20496 6100 20502 6112
rect 21836 6100 21864 6140
rect 38010 6128 38016 6140
rect 38068 6128 38074 6180
rect 20496 6072 21864 6100
rect 22649 6103 22707 6109
rect 20496 6060 20502 6072
rect 22649 6069 22661 6103
rect 22695 6100 22707 6103
rect 22922 6100 22928 6112
rect 22695 6072 22928 6100
rect 22695 6069 22707 6072
rect 22649 6063 22707 6069
rect 22922 6060 22928 6072
rect 22980 6060 22986 6112
rect 23106 6100 23112 6112
rect 23067 6072 23112 6100
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 24946 6060 24952 6112
rect 25004 6100 25010 6112
rect 32401 6103 32459 6109
rect 32401 6100 32413 6103
rect 25004 6072 32413 6100
rect 25004 6060 25010 6072
rect 32401 6069 32413 6072
rect 32447 6069 32459 6103
rect 32401 6063 32459 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1844 5899 1902 5905
rect 1844 5865 1856 5899
rect 1890 5896 1902 5899
rect 3050 5896 3056 5908
rect 1890 5868 3056 5896
rect 1890 5865 1902 5868
rect 1844 5859 1902 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 3418 5896 3424 5908
rect 3375 5868 3424 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 6730 5896 6736 5908
rect 4028 5868 6736 5896
rect 4028 5856 4034 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7064 5868 8064 5896
rect 7064 5856 7070 5868
rect 5350 5788 5356 5840
rect 5408 5788 5414 5840
rect 5718 5828 5724 5840
rect 5679 5800 5724 5828
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 8036 5837 8064 5868
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 9030 5896 9036 5908
rect 8536 5868 9036 5896
rect 8536 5856 8542 5868
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 9398 5896 9404 5908
rect 9263 5868 9404 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 10045 5899 10103 5905
rect 9508 5868 9996 5896
rect 8021 5831 8079 5837
rect 8021 5797 8033 5831
rect 8067 5828 8079 5831
rect 9508 5828 9536 5868
rect 8067 5800 9536 5828
rect 9968 5828 9996 5868
rect 10045 5865 10057 5899
rect 10091 5896 10103 5899
rect 10318 5896 10324 5908
rect 10091 5868 10324 5896
rect 10091 5865 10103 5868
rect 10045 5859 10103 5865
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 16850 5896 16856 5908
rect 10428 5868 16856 5896
rect 10428 5828 10456 5868
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 16945 5899 17003 5905
rect 16945 5865 16957 5899
rect 16991 5896 17003 5899
rect 17034 5896 17040 5908
rect 16991 5868 17040 5896
rect 16991 5865 17003 5868
rect 16945 5859 17003 5865
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17862 5856 17868 5908
rect 17920 5896 17926 5908
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 17920 5868 18153 5896
rect 17920 5856 17926 5868
rect 18141 5865 18153 5868
rect 18187 5865 18199 5899
rect 18141 5859 18199 5865
rect 18690 5856 18696 5908
rect 18748 5896 18754 5908
rect 18785 5899 18843 5905
rect 18785 5896 18797 5899
rect 18748 5868 18797 5896
rect 18748 5856 18754 5868
rect 18785 5865 18797 5868
rect 18831 5865 18843 5899
rect 18785 5859 18843 5865
rect 18874 5856 18880 5908
rect 18932 5896 18938 5908
rect 19978 5896 19984 5908
rect 18932 5868 19984 5896
rect 18932 5856 18938 5868
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20073 5899 20131 5905
rect 20073 5865 20085 5899
rect 20119 5896 20131 5899
rect 20346 5896 20352 5908
rect 20119 5868 20352 5896
rect 20119 5865 20131 5868
rect 20073 5859 20131 5865
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 21453 5899 21511 5905
rect 21453 5896 21465 5899
rect 20772 5868 21465 5896
rect 20772 5856 20778 5868
rect 21453 5865 21465 5868
rect 21499 5865 21511 5899
rect 21453 5859 21511 5865
rect 21726 5856 21732 5908
rect 21784 5896 21790 5908
rect 23842 5896 23848 5908
rect 21784 5868 23848 5896
rect 21784 5856 21790 5868
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 37550 5856 37556 5908
rect 37608 5896 37614 5908
rect 37645 5899 37703 5905
rect 37645 5896 37657 5899
rect 37608 5868 37657 5896
rect 37608 5856 37614 5868
rect 37645 5865 37657 5868
rect 37691 5865 37703 5899
rect 37645 5859 37703 5865
rect 12342 5828 12348 5840
rect 9968 5800 10456 5828
rect 10612 5800 11652 5828
rect 12303 5800 12348 5828
rect 8067 5797 8079 5800
rect 8021 5791 8079 5797
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5760 1642 5772
rect 4249 5763 4307 5769
rect 1636 5732 4016 5760
rect 1636 5720 1642 5732
rect 3988 5704 4016 5732
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4982 5760 4988 5772
rect 4295 5732 4988 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4982 5720 4988 5732
rect 5040 5720 5046 5772
rect 5368 5760 5396 5788
rect 6270 5760 6276 5772
rect 5368 5732 6276 5760
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6546 5760 6552 5772
rect 6459 5732 6552 5760
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 10612 5760 10640 5800
rect 6604 5732 10640 5760
rect 6604 5720 6610 5732
rect 11238 5720 11244 5772
rect 11296 5720 11302 5772
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8662 5692 8668 5704
rect 7892 5664 8668 5692
rect 7892 5652 7898 5664
rect 8662 5652 8668 5664
rect 8720 5652 8726 5704
rect 9122 5692 9128 5704
rect 9083 5664 9128 5692
rect 9122 5652 9128 5664
rect 9180 5692 9186 5704
rect 9950 5692 9956 5704
rect 9180 5664 9956 5692
rect 9180 5652 9186 5664
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10100 5664 10732 5692
rect 10100 5652 10106 5664
rect 6822 5624 6828 5636
rect 3082 5596 4660 5624
rect 5474 5596 6828 5624
rect 4632 5556 4660 5596
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 10318 5624 10324 5636
rect 7774 5596 10324 5624
rect 10318 5584 10324 5596
rect 10376 5584 10382 5636
rect 10704 5624 10732 5664
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10836 5664 10977 5692
rect 10836 5652 10842 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5692 11115 5695
rect 11256 5692 11284 5720
rect 11624 5701 11652 5800
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 13998 5828 14004 5840
rect 12584 5800 14004 5828
rect 12584 5788 12590 5800
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 14366 5828 14372 5840
rect 14327 5800 14372 5828
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 14642 5788 14648 5840
rect 14700 5828 14706 5840
rect 23106 5828 23112 5840
rect 14700 5800 23112 5828
rect 14700 5788 14706 5800
rect 23106 5788 23112 5800
rect 23164 5788 23170 5840
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 13081 5763 13139 5769
rect 13081 5760 13093 5763
rect 12676 5732 13093 5760
rect 12676 5720 12682 5732
rect 13081 5729 13093 5732
rect 13127 5729 13139 5763
rect 13081 5723 13139 5729
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14240 5732 17816 5760
rect 14240 5720 14246 5732
rect 11103 5664 11284 5692
rect 11609 5695 11667 5701
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 11609 5661 11621 5695
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 11848 5664 12265 5692
rect 11848 5652 11854 5664
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12860 5664 12909 5692
rect 12860 5652 12866 5664
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 14274 5692 14280 5704
rect 12897 5655 12955 5661
rect 13004 5664 14280 5692
rect 10704 5596 11192 5624
rect 10870 5556 10876 5568
rect 4632 5528 10876 5556
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 11164 5556 11192 5596
rect 11238 5584 11244 5636
rect 11296 5624 11302 5636
rect 12342 5624 12348 5636
rect 11296 5596 12348 5624
rect 11296 5584 11302 5596
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 13004 5624 13032 5664
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 16850 5692 16856 5704
rect 16172 5664 16856 5692
rect 16172 5652 16178 5664
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17788 5692 17816 5732
rect 17862 5720 17868 5772
rect 17920 5760 17926 5772
rect 19794 5760 19800 5772
rect 17920 5732 19800 5760
rect 17920 5720 17926 5732
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 19886 5720 19892 5772
rect 19944 5760 19950 5772
rect 21174 5760 21180 5772
rect 19944 5732 21180 5760
rect 19944 5720 19950 5732
rect 21174 5720 21180 5732
rect 21232 5720 21238 5772
rect 21910 5720 21916 5772
rect 21968 5760 21974 5772
rect 37660 5760 37688 5859
rect 21968 5732 23336 5760
rect 37660 5732 38056 5760
rect 21968 5720 21974 5732
rect 18049 5695 18107 5701
rect 17788 5664 18000 5692
rect 12820 5596 13032 5624
rect 11606 5556 11612 5568
rect 11164 5528 11612 5556
rect 11606 5516 11612 5528
rect 11664 5516 11670 5568
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 11882 5556 11888 5568
rect 11747 5528 11888 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 12820 5556 12848 5596
rect 13998 5584 14004 5636
rect 14056 5624 14062 5636
rect 15010 5624 15016 5636
rect 14056 5596 14504 5624
rect 14971 5596 15016 5624
rect 14056 5584 14062 5596
rect 12676 5528 12848 5556
rect 14476 5556 14504 5596
rect 15010 5584 15016 5596
rect 15068 5584 15074 5636
rect 15102 5584 15108 5636
rect 15160 5624 15166 5636
rect 15160 5596 15205 5624
rect 15160 5584 15166 5596
rect 15838 5584 15844 5636
rect 15896 5624 15902 5636
rect 16025 5627 16083 5633
rect 16025 5624 16037 5627
rect 15896 5596 16037 5624
rect 15896 5584 15902 5596
rect 16025 5593 16037 5596
rect 16071 5593 16083 5627
rect 17862 5624 17868 5636
rect 16025 5587 16083 5593
rect 16132 5596 17868 5624
rect 16132 5556 16160 5596
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 17972 5624 18000 5664
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18230 5692 18236 5704
rect 18095 5664 18236 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18690 5692 18696 5704
rect 18651 5664 18696 5692
rect 18690 5652 18696 5664
rect 18748 5652 18754 5704
rect 18782 5652 18788 5704
rect 18840 5692 18846 5704
rect 19981 5695 20039 5701
rect 19981 5692 19993 5695
rect 18840 5664 19993 5692
rect 18840 5652 18846 5664
rect 19981 5661 19993 5664
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 20070 5652 20076 5704
rect 20128 5692 20134 5704
rect 20709 5695 20767 5701
rect 20709 5692 20721 5695
rect 20128 5664 20721 5692
rect 20128 5652 20134 5664
rect 20709 5661 20721 5664
rect 20755 5661 20767 5695
rect 20709 5655 20767 5661
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 20864 5664 20909 5692
rect 20864 5652 20870 5664
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 21048 5664 21373 5692
rect 21048 5652 21054 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 22186 5692 22192 5704
rect 22147 5664 22192 5692
rect 21361 5655 21419 5661
rect 22186 5652 22192 5664
rect 22244 5652 22250 5704
rect 22646 5692 22652 5704
rect 22607 5664 22652 5692
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 23308 5701 23336 5732
rect 23293 5695 23351 5701
rect 23293 5661 23305 5695
rect 23339 5661 23351 5695
rect 23293 5655 23351 5661
rect 37369 5695 37427 5701
rect 37369 5661 37381 5695
rect 37415 5692 37427 5695
rect 37734 5692 37740 5704
rect 37415 5664 37740 5692
rect 37415 5661 37427 5664
rect 37369 5655 37427 5661
rect 37734 5652 37740 5664
rect 37792 5652 37798 5704
rect 38028 5701 38056 5732
rect 38013 5695 38071 5701
rect 38013 5661 38025 5695
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 22741 5627 22799 5633
rect 22741 5624 22753 5627
rect 17972 5596 20208 5624
rect 14476 5528 16160 5556
rect 12676 5516 12682 5528
rect 16850 5516 16856 5568
rect 16908 5556 16914 5568
rect 20070 5556 20076 5568
rect 16908 5528 20076 5556
rect 16908 5516 16914 5528
rect 20070 5516 20076 5528
rect 20128 5516 20134 5568
rect 20180 5556 20208 5596
rect 20732 5596 22753 5624
rect 20732 5556 20760 5596
rect 22741 5593 22753 5596
rect 22787 5593 22799 5627
rect 22741 5587 22799 5593
rect 22002 5556 22008 5568
rect 20180 5528 20760 5556
rect 21963 5528 22008 5556
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 23382 5556 23388 5568
rect 23343 5528 23388 5556
rect 23382 5516 23388 5528
rect 23440 5516 23446 5568
rect 37185 5559 37243 5565
rect 37185 5525 37197 5559
rect 37231 5556 37243 5559
rect 37550 5556 37556 5568
rect 37231 5528 37556 5556
rect 37231 5525 37243 5528
rect 37185 5519 37243 5525
rect 37550 5516 37556 5528
rect 37608 5516 37614 5568
rect 38194 5556 38200 5568
rect 38155 5528 38200 5556
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 5902 5352 5908 5364
rect 4908 5324 5908 5352
rect 2222 5244 2228 5296
rect 2280 5284 2286 5296
rect 2317 5287 2375 5293
rect 2317 5284 2329 5287
rect 2280 5256 2329 5284
rect 2280 5244 2286 5256
rect 2317 5253 2329 5256
rect 2363 5253 2375 5287
rect 4908 5284 4936 5324
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6546 5352 6552 5364
rect 6043 5324 6552 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 6914 5352 6920 5364
rect 6840 5324 6920 5352
rect 6086 5284 6092 5296
rect 3542 5256 4936 5284
rect 5750 5256 6092 5284
rect 2317 5247 2375 5253
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 6270 5244 6276 5296
rect 6328 5284 6334 5296
rect 6454 5284 6460 5296
rect 6328 5256 6460 5284
rect 6328 5244 6334 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6840 5293 6868 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 8846 5352 8852 5364
rect 7156 5324 8294 5352
rect 8807 5324 8852 5352
rect 7156 5312 7162 5324
rect 6825 5287 6883 5293
rect 6825 5253 6837 5287
rect 6871 5253 6883 5287
rect 8266 5284 8294 5324
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9398 5352 9404 5364
rect 9232 5324 9404 5352
rect 9232 5284 9260 5324
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 9582 5352 9588 5364
rect 9539 5324 9588 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 11054 5352 11060 5364
rect 10100 5324 10548 5352
rect 11015 5324 11060 5352
rect 10100 5312 10106 5324
rect 8266 5256 9260 5284
rect 9324 5256 9720 5284
rect 6825 5247 6883 5253
rect 1578 5176 1584 5228
rect 1636 5216 1642 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1636 5188 2053 5216
rect 1636 5176 1642 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 8478 5216 8484 5228
rect 7958 5188 8484 5216
rect 2041 5179 2099 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9214 5216 9220 5228
rect 8803 5188 9220 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 4062 5148 4068 5160
rect 2924 5120 4068 5148
rect 2924 5108 2930 5120
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4249 5151 4307 5157
rect 4249 5148 4261 5151
rect 4212 5120 4261 5148
rect 4212 5108 4218 5120
rect 4249 5117 4261 5120
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4982 5148 4988 5160
rect 4571 5120 4988 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 3789 5015 3847 5021
rect 3789 4981 3801 5015
rect 3835 5012 3847 5015
rect 3878 5012 3884 5024
rect 3835 4984 3884 5012
rect 3835 4981 3847 4984
rect 3789 4975 3847 4981
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 4264 5012 4292 5111
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 6535 5108 6541 5160
rect 6593 5157 6599 5160
rect 6593 5151 6607 5157
rect 6595 5148 6607 5151
rect 6595 5120 6638 5148
rect 6595 5117 6607 5120
rect 6593 5111 6607 5117
rect 6593 5108 6599 5111
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 9324 5148 9352 5256
rect 9393 5217 9451 5223
rect 9393 5183 9405 5217
rect 9439 5216 9451 5217
rect 9582 5216 9588 5228
rect 9439 5188 9588 5216
rect 9439 5183 9451 5188
rect 9393 5177 9451 5183
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 6972 5120 9352 5148
rect 9692 5148 9720 5256
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10520 5284 10548 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11790 5352 11796 5364
rect 11164 5324 11796 5352
rect 11164 5284 11192 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 11940 5324 12480 5352
rect 11940 5312 11946 5324
rect 12345 5287 12403 5293
rect 12345 5284 12357 5287
rect 10008 5256 10456 5284
rect 10520 5256 11192 5284
rect 11256 5256 12357 5284
rect 10008 5244 10014 5256
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10100 5188 10333 5216
rect 10100 5176 10106 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10428 5216 10456 5256
rect 10686 5216 10692 5228
rect 10428 5188 10692 5216
rect 10321 5179 10379 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10836 5188 10977 5216
rect 10836 5176 10842 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11256 5148 11284 5256
rect 12345 5253 12357 5256
rect 12391 5253 12403 5287
rect 12452 5284 12480 5324
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12584 5324 13001 5352
rect 12584 5312 12590 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 13096 5324 13768 5352
rect 13096 5284 13124 5324
rect 12452 5256 13124 5284
rect 12345 5247 12403 5253
rect 13170 5244 13176 5296
rect 13228 5284 13234 5296
rect 13633 5287 13691 5293
rect 13633 5284 13645 5287
rect 13228 5256 13645 5284
rect 13228 5244 13234 5256
rect 13633 5253 13645 5256
rect 13679 5253 13691 5287
rect 13633 5247 13691 5253
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 9692 5120 11284 5148
rect 11532 5188 12265 5216
rect 6972 5108 6978 5120
rect 6362 5080 6368 5092
rect 5644 5052 6368 5080
rect 4614 5012 4620 5024
rect 4264 4984 4620 5012
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5644 5012 5672 5052
rect 6362 5040 6368 5052
rect 6420 5040 6426 5092
rect 11238 5080 11244 5092
rect 8220 5052 11244 5080
rect 5040 4984 5672 5012
rect 5040 4972 5046 4984
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 8220 5012 8248 5052
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 5776 4984 8248 5012
rect 8297 5015 8355 5021
rect 5776 4972 5782 4984
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 8386 5012 8392 5024
rect 8343 4984 8392 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 9732 4984 10425 5012
rect 9732 4972 9738 4984
rect 10413 4981 10425 4984
rect 10459 4981 10471 5015
rect 10413 4975 10471 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11532 5012 11560 5188
rect 12253 5185 12265 5188
rect 12299 5216 12311 5219
rect 12897 5219 12955 5225
rect 12299 5188 12388 5216
rect 12897 5214 12909 5219
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12360 5148 12388 5188
rect 12820 5186 12909 5214
rect 12618 5148 12624 5160
rect 12360 5120 12624 5148
rect 12618 5108 12624 5120
rect 12676 5148 12682 5160
rect 12820 5148 12848 5186
rect 12897 5185 12909 5186
rect 12943 5185 12955 5219
rect 13541 5219 13599 5225
rect 13541 5216 13553 5219
rect 12897 5179 12955 5185
rect 13188 5188 13553 5216
rect 13188 5160 13216 5188
rect 13541 5185 13553 5188
rect 13587 5185 13599 5219
rect 13740 5216 13768 5324
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 14148 5324 14289 5352
rect 14148 5312 14154 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14424 5324 14933 5352
rect 14424 5312 14430 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15252 5324 15516 5352
rect 15252 5312 15258 5324
rect 14458 5244 14464 5296
rect 14516 5284 14522 5296
rect 15488 5284 15516 5324
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16209 5355 16267 5361
rect 16209 5352 16221 5355
rect 15804 5324 16221 5352
rect 15804 5312 15810 5324
rect 16209 5321 16221 5324
rect 16255 5321 16267 5355
rect 16209 5315 16267 5321
rect 16482 5312 16488 5364
rect 16540 5352 16546 5364
rect 17402 5352 17408 5364
rect 16540 5324 17408 5352
rect 16540 5312 16546 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 19429 5355 19487 5361
rect 18196 5324 19334 5352
rect 18196 5312 18202 5324
rect 18785 5287 18843 5293
rect 14516 5256 15194 5284
rect 15488 5256 18736 5284
rect 14516 5244 14522 5256
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13740 5188 14197 5216
rect 13541 5179 13599 5185
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14332 5188 14841 5216
rect 14332 5176 14338 5188
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 15166 5216 15194 5256
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15166 5188 15485 5216
rect 14829 5179 14887 5185
rect 15473 5185 15485 5188
rect 15519 5216 15531 5219
rect 15746 5216 15752 5228
rect 15519 5188 15752 5216
rect 15519 5185 15531 5188
rect 15473 5179 15531 5185
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 16114 5216 16120 5228
rect 16075 5188 16120 5216
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 16298 5176 16304 5228
rect 16356 5216 16362 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 16356 5188 17417 5216
rect 16356 5176 16362 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17828 5188 18061 5216
rect 17828 5176 17834 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18708 5225 18736 5256
rect 18785 5253 18797 5287
rect 18831 5284 18843 5287
rect 19150 5284 19156 5296
rect 18831 5256 19156 5284
rect 18831 5253 18843 5256
rect 18785 5247 18843 5253
rect 19150 5244 19156 5256
rect 19208 5244 19214 5296
rect 19306 5284 19334 5324
rect 19429 5321 19441 5355
rect 19475 5352 19487 5355
rect 24118 5352 24124 5364
rect 19475 5324 24124 5352
rect 19475 5321 19487 5324
rect 19429 5315 19487 5321
rect 24118 5312 24124 5324
rect 24176 5312 24182 5364
rect 21913 5287 21971 5293
rect 21913 5284 21925 5287
rect 19306 5256 21925 5284
rect 21913 5253 21925 5256
rect 21959 5253 21971 5287
rect 21913 5247 21971 5253
rect 18693 5219 18751 5225
rect 18196 5188 18241 5216
rect 18196 5176 18202 5188
rect 18693 5185 18705 5219
rect 18739 5185 18751 5219
rect 19337 5219 19395 5225
rect 19337 5214 19349 5219
rect 18693 5179 18751 5185
rect 19260 5186 19349 5214
rect 12676 5120 12848 5148
rect 12676 5108 12682 5120
rect 13170 5108 13176 5160
rect 13228 5108 13234 5160
rect 13280 5120 15700 5148
rect 11606 5040 11612 5092
rect 11664 5080 11670 5092
rect 11664 5052 12388 5080
rect 11664 5040 11670 5052
rect 10744 4984 11560 5012
rect 10744 4972 10750 4984
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 12158 5012 12164 5024
rect 11756 4984 12164 5012
rect 11756 4972 11762 4984
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12360 5012 12388 5052
rect 13280 5012 13308 5120
rect 15565 5083 15623 5089
rect 15565 5080 15577 5083
rect 13832 5052 15577 5080
rect 12360 4984 13308 5012
rect 13446 4972 13452 5024
rect 13504 5012 13510 5024
rect 13832 5012 13860 5052
rect 15565 5049 15577 5052
rect 15611 5049 15623 5083
rect 15672 5080 15700 5120
rect 17494 5108 17500 5160
rect 17552 5148 17558 5160
rect 18598 5148 18604 5160
rect 17552 5120 17597 5148
rect 17696 5120 18604 5148
rect 17552 5108 17558 5120
rect 17696 5080 17724 5120
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 19260 5148 19288 5186
rect 19337 5185 19349 5186
rect 19383 5185 19395 5219
rect 19337 5179 19395 5185
rect 20073 5219 20131 5225
rect 20073 5185 20085 5219
rect 20119 5216 20131 5219
rect 20254 5216 20260 5228
rect 20119 5188 20260 5216
rect 20119 5185 20131 5188
rect 20073 5179 20131 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5185 20775 5219
rect 21818 5216 21824 5228
rect 21779 5188 21824 5216
rect 20717 5179 20775 5185
rect 18708 5120 19288 5148
rect 15672 5052 17724 5080
rect 15565 5043 15623 5049
rect 17862 5040 17868 5092
rect 17920 5080 17926 5092
rect 18230 5080 18236 5092
rect 17920 5052 18236 5080
rect 17920 5040 17926 5052
rect 18230 5040 18236 5052
rect 18288 5040 18294 5092
rect 13504 4984 13860 5012
rect 13504 4972 13510 4984
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 18708 5012 18736 5120
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 20732 5148 20760 5179
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 22278 5176 22284 5228
rect 22336 5216 22342 5228
rect 22833 5219 22891 5225
rect 22833 5216 22845 5219
rect 22336 5188 22845 5216
rect 22336 5176 22342 5188
rect 22833 5185 22845 5188
rect 22879 5185 22891 5219
rect 22833 5179 22891 5185
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 23293 5219 23351 5225
rect 23293 5216 23305 5219
rect 22980 5188 23305 5216
rect 22980 5176 22986 5188
rect 23293 5185 23305 5188
rect 23339 5185 23351 5219
rect 23293 5179 23351 5185
rect 32398 5176 32404 5228
rect 32456 5216 32462 5228
rect 38013 5219 38071 5225
rect 38013 5216 38025 5219
rect 32456 5188 38025 5216
rect 32456 5176 32462 5188
rect 38013 5185 38025 5188
rect 38059 5185 38071 5219
rect 38013 5179 38071 5185
rect 19484 5120 20760 5148
rect 19484 5108 19490 5120
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 23385 5151 23443 5157
rect 23385 5148 23397 5151
rect 20864 5120 23397 5148
rect 20864 5108 20870 5120
rect 23385 5117 23397 5120
rect 23431 5117 23443 5151
rect 23385 5111 23443 5117
rect 18782 5040 18788 5092
rect 18840 5080 18846 5092
rect 19242 5080 19248 5092
rect 18840 5052 19248 5080
rect 18840 5040 18846 5052
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 20165 5083 20223 5089
rect 20165 5080 20177 5083
rect 19444 5052 20177 5080
rect 13964 4984 18736 5012
rect 13964 4972 13970 4984
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 19444 5012 19472 5052
rect 20165 5049 20177 5052
rect 20211 5049 20223 5083
rect 20165 5043 20223 5049
rect 20530 5040 20536 5092
rect 20588 5080 20594 5092
rect 22649 5083 22707 5089
rect 22649 5080 22661 5083
rect 20588 5052 22661 5080
rect 20588 5040 20594 5052
rect 22649 5049 22661 5052
rect 22695 5049 22707 5083
rect 22649 5043 22707 5049
rect 19024 4984 19472 5012
rect 19024 4972 19030 4984
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19978 5012 19984 5024
rect 19576 4984 19984 5012
rect 19576 4972 19582 4984
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20438 4972 20444 5024
rect 20496 5012 20502 5024
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20496 4984 20821 5012
rect 20496 4972 20502 4984
rect 20809 4981 20821 4984
rect 20855 4981 20867 5015
rect 22278 5012 22284 5024
rect 22239 4984 22284 5012
rect 20809 4975 20867 4981
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 38194 5012 38200 5024
rect 38155 4984 38200 5012
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 2556 4780 7604 4808
rect 2556 4768 2562 4780
rect 3326 4700 3332 4752
rect 3384 4740 3390 4752
rect 3421 4743 3479 4749
rect 3421 4740 3433 4743
rect 3384 4712 3433 4740
rect 3384 4700 3390 4712
rect 3421 4709 3433 4712
rect 3467 4709 3479 4743
rect 3421 4703 3479 4709
rect 3786 4700 3792 4752
rect 3844 4740 3850 4752
rect 4893 4743 4951 4749
rect 4893 4740 4905 4743
rect 3844 4712 4905 4740
rect 3844 4700 3850 4712
rect 4893 4709 4905 4712
rect 4939 4709 4951 4743
rect 7282 4740 7288 4752
rect 7243 4712 7288 4740
rect 4893 4703 4951 4709
rect 7282 4700 7288 4712
rect 7340 4700 7346 4752
rect 7576 4740 7604 4780
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7708 4780 7849 4808
rect 7708 4768 7714 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8481 4811 8539 4817
rect 8260 4780 8432 4808
rect 8260 4768 8266 4780
rect 8294 4740 8300 4752
rect 7576 4712 8300 4740
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8404 4740 8432 4780
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 8754 4808 8760 4820
rect 8527 4780 8760 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 8938 4768 8944 4820
rect 8996 4808 9002 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 8996 4780 9229 4808
rect 8996 4768 9002 4780
rect 9217 4777 9229 4780
rect 9263 4777 9275 4811
rect 9217 4771 9275 4777
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 10413 4811 10471 4817
rect 9456 4780 10364 4808
rect 9456 4768 9462 4780
rect 10336 4740 10364 4780
rect 10413 4777 10425 4811
rect 10459 4808 10471 4811
rect 10594 4808 10600 4820
rect 10459 4780 10600 4808
rect 10459 4777 10471 4780
rect 10413 4771 10471 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 10888 4780 11376 4808
rect 10888 4740 10916 4780
rect 8404 4712 10272 4740
rect 10336 4712 10916 4740
rect 1578 4632 1584 4684
rect 1636 4672 1642 4684
rect 1673 4675 1731 4681
rect 1673 4672 1685 4675
rect 1636 4644 1685 4672
rect 1636 4632 1642 4644
rect 1673 4641 1685 4644
rect 1719 4641 1731 4675
rect 1673 4635 1731 4641
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 2038 4672 2044 4684
rect 1995 4644 2044 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 10244 4672 10272 4712
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 11057 4743 11115 4749
rect 11057 4740 11069 4743
rect 11020 4712 11069 4740
rect 11020 4700 11026 4712
rect 11057 4709 11069 4712
rect 11103 4709 11115 4743
rect 11057 4703 11115 4709
rect 3016 4644 8432 4672
rect 10244 4644 10548 4672
rect 3016 4632 3022 4644
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 4430 4604 4436 4616
rect 3835 4576 4436 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4604 4770 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4764 4576 5273 4604
rect 4764 4564 4770 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5408 4576 5549 4604
rect 5408 4564 5414 4576
rect 5537 4573 5549 4576
rect 5583 4573 5595 4607
rect 5537 4567 5595 4573
rect 7190 4564 7196 4616
rect 7248 4604 7254 4616
rect 7650 4604 7656 4616
rect 7248 4576 7656 4604
rect 7248 4564 7254 4576
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 8202 4604 8208 4616
rect 7791 4576 8208 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8404 4613 8432 4644
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8938 4564 8944 4616
rect 8996 4604 9002 4616
rect 9125 4607 9183 4613
rect 9125 4604 9137 4607
rect 8996 4576 9137 4604
rect 8996 4564 9002 4576
rect 9125 4573 9137 4576
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10321 4607 10379 4613
rect 10321 4604 10333 4607
rect 10008 4576 10333 4604
rect 10008 4564 10014 4576
rect 10321 4573 10333 4576
rect 10367 4573 10379 4607
rect 10520 4604 10548 4644
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 11348 4672 11376 4780
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 11572 4780 11713 4808
rect 11572 4768 11578 4780
rect 11701 4777 11713 4780
rect 11747 4777 11759 4811
rect 11701 4771 11759 4777
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 12434 4808 12440 4820
rect 11848 4780 12440 4808
rect 11848 4768 11854 4780
rect 12434 4768 12440 4780
rect 12492 4808 12498 4820
rect 12802 4808 12808 4820
rect 12492 4780 12808 4808
rect 12492 4768 12498 4780
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12986 4808 12992 4820
rect 12947 4780 12992 4808
rect 12986 4768 12992 4780
rect 13044 4768 13050 4820
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 16482 4808 16488 4820
rect 14752 4780 16488 4808
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 11480 4712 13645 4740
rect 11480 4700 11486 4712
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 14458 4740 14464 4752
rect 13633 4703 13691 4709
rect 14108 4712 14464 4740
rect 10744 4644 11100 4672
rect 11348 4644 13124 4672
rect 10744 4632 10750 4644
rect 10870 4604 10876 4616
rect 10520 4576 10876 4604
rect 10321 4567 10379 4573
rect 10870 4564 10876 4576
rect 10928 4604 10934 4616
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 10928 4576 10977 4604
rect 10928 4564 10934 4576
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 11072 4604 11100 4644
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11072 4576 11621 4604
rect 10965 4567 11023 4573
rect 11609 4573 11621 4576
rect 11655 4604 11667 4607
rect 11790 4604 11796 4616
rect 11655 4576 11796 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 12250 4604 12256 4616
rect 12211 4576 12256 4604
rect 12250 4564 12256 4576
rect 12308 4604 12314 4616
rect 12308 4576 12480 4604
rect 12308 4564 12314 4576
rect 5718 4536 5724 4548
rect 3174 4508 5724 4536
rect 5718 4496 5724 4508
rect 5776 4496 5782 4548
rect 5813 4539 5871 4545
rect 5813 4505 5825 4539
rect 5859 4505 5871 4539
rect 9674 4536 9680 4548
rect 7038 4508 9680 4536
rect 5813 4499 5871 4505
rect 3970 4468 3976 4480
rect 3931 4440 3976 4468
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 4430 4468 4436 4480
rect 4343 4440 4436 4468
rect 4430 4428 4436 4440
rect 4488 4468 4494 4480
rect 4798 4468 4804 4480
rect 4488 4440 4804 4468
rect 4488 4428 4494 4440
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5828 4468 5856 4499
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 9824 4508 11744 4536
rect 9824 4496 9830 4508
rect 8386 4468 8392 4480
rect 5828 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 11606 4468 11612 4480
rect 8996 4440 11612 4468
rect 8996 4428 9002 4440
rect 11606 4428 11612 4440
rect 11664 4428 11670 4480
rect 11716 4468 11744 4508
rect 12066 4496 12072 4548
rect 12124 4536 12130 4548
rect 12345 4539 12403 4545
rect 12345 4536 12357 4539
rect 12124 4508 12357 4536
rect 12124 4496 12130 4508
rect 12345 4505 12357 4508
rect 12391 4505 12403 4539
rect 12452 4536 12480 4576
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 12897 4607 12955 4613
rect 12897 4604 12909 4607
rect 12584 4576 12909 4604
rect 12584 4564 12590 4576
rect 12897 4573 12909 4576
rect 12943 4604 12955 4607
rect 12986 4604 12992 4616
rect 12943 4576 12992 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 12710 4536 12716 4548
rect 12452 4508 12716 4536
rect 12345 4499 12403 4505
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 13096 4536 13124 4644
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13446 4672 13452 4684
rect 13228 4644 13452 4672
rect 13228 4632 13234 4644
rect 13446 4632 13452 4644
rect 13504 4672 13510 4684
rect 14108 4672 14136 4712
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 13504 4644 14136 4672
rect 13504 4632 13510 4644
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 14642 4672 14648 4684
rect 14240 4644 14648 4672
rect 14240 4632 14246 4644
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13906 4604 13912 4616
rect 13587 4576 13912 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14056 4576 14565 4604
rect 14056 4564 14062 4576
rect 14553 4573 14565 4576
rect 14599 4604 14611 4607
rect 14752 4604 14780 4780
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 16666 4768 16672 4820
rect 16724 4808 16730 4820
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 16724 4780 17877 4808
rect 16724 4768 16730 4780
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 20809 4811 20867 4817
rect 20809 4808 20821 4811
rect 17865 4771 17923 4777
rect 17972 4780 20821 4808
rect 15010 4700 15016 4752
rect 15068 4740 15074 4752
rect 16577 4743 16635 4749
rect 15068 4712 16344 4740
rect 15068 4700 15074 4712
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 14599 4576 14780 4604
rect 14599 4573 14611 4576
rect 14553 4567 14611 4573
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15197 4607 15255 4613
rect 15197 4604 15209 4607
rect 15068 4576 15209 4604
rect 15068 4564 15074 4576
rect 15197 4573 15209 4576
rect 15243 4573 15255 4607
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15197 4567 15255 4573
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 13170 4536 13176 4548
rect 13096 4508 13176 4536
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 15933 4539 15991 4545
rect 15933 4536 15945 4539
rect 13780 4508 15945 4536
rect 13780 4496 13786 4508
rect 15933 4505 15945 4508
rect 15979 4505 15991 4539
rect 16316 4536 16344 4712
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 16758 4740 16764 4752
rect 16623 4712 16764 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 17034 4700 17040 4752
rect 17092 4740 17098 4752
rect 17221 4743 17279 4749
rect 17221 4740 17233 4743
rect 17092 4712 17233 4740
rect 17092 4700 17098 4712
rect 17221 4709 17233 4712
rect 17267 4709 17279 4743
rect 17221 4703 17279 4709
rect 17402 4700 17408 4752
rect 17460 4740 17466 4752
rect 17770 4740 17776 4752
rect 17460 4712 17776 4740
rect 17460 4700 17466 4712
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 17972 4672 18000 4780
rect 20809 4777 20821 4780
rect 20855 4777 20867 4811
rect 20809 4771 20867 4777
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22152 4780 22197 4808
rect 22152 4768 22158 4780
rect 18509 4743 18567 4749
rect 18509 4709 18521 4743
rect 18555 4740 18567 4743
rect 22370 4740 22376 4752
rect 18555 4712 22376 4740
rect 18555 4709 18567 4712
rect 18509 4703 18567 4709
rect 22370 4700 22376 4712
rect 22428 4700 22434 4752
rect 21361 4675 21419 4681
rect 21361 4672 21373 4675
rect 16724 4644 18000 4672
rect 18064 4644 21373 4672
rect 16724 4632 16730 4644
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16448 4576 16497 4604
rect 16448 4564 16454 4576
rect 16485 4573 16497 4576
rect 16531 4604 16543 4607
rect 17129 4607 17187 4613
rect 17129 4604 17141 4607
rect 16531 4576 17141 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 17129 4573 17141 4576
rect 17175 4573 17187 4607
rect 17770 4604 17776 4616
rect 17731 4576 17776 4604
rect 17129 4567 17187 4573
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 18064 4536 18092 4644
rect 21361 4641 21373 4644
rect 21407 4641 21419 4675
rect 23474 4672 23480 4684
rect 21361 4635 21419 4641
rect 22664 4644 23480 4672
rect 18322 4564 18328 4616
rect 18380 4604 18386 4616
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 18380 4576 18429 4604
rect 18380 4564 18386 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 20073 4607 20131 4613
rect 20073 4604 20085 4607
rect 19668 4576 20085 4604
rect 19668 4564 19674 4576
rect 20073 4573 20085 4576
rect 20119 4604 20131 4607
rect 20717 4607 20775 4613
rect 20119 4576 20300 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 19518 4536 19524 4548
rect 16316 4508 18092 4536
rect 19479 4508 19524 4536
rect 15933 4499 15991 4505
rect 19518 4496 19524 4508
rect 19576 4496 19582 4548
rect 20162 4536 20168 4548
rect 20123 4508 20168 4536
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 20272 4536 20300 4576
rect 20717 4573 20729 4607
rect 20763 4604 20775 4607
rect 20806 4604 20812 4616
rect 20763 4576 20812 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 21174 4564 21180 4616
rect 21232 4604 21238 4616
rect 21818 4604 21824 4616
rect 21232 4576 21824 4604
rect 21232 4564 21238 4576
rect 21818 4564 21824 4576
rect 21876 4604 21882 4616
rect 22664 4613 22692 4644
rect 23474 4632 23480 4644
rect 23532 4632 23538 4684
rect 22005 4607 22063 4613
rect 22005 4604 22017 4607
rect 21876 4576 22017 4604
rect 21876 4564 21882 4576
rect 22005 4573 22017 4576
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 22649 4607 22707 4613
rect 22649 4573 22661 4607
rect 22695 4573 22707 4607
rect 22649 4567 22707 4573
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4573 23351 4607
rect 31294 4604 31300 4616
rect 31255 4576 31300 4604
rect 23293 4567 23351 4573
rect 21082 4536 21088 4548
rect 20272 4508 21088 4536
rect 21082 4496 21088 4508
rect 21140 4496 21146 4548
rect 21358 4496 21364 4548
rect 21416 4536 21422 4548
rect 23308 4536 23336 4567
rect 31294 4564 31300 4576
rect 31352 4564 31358 4616
rect 38013 4607 38071 4613
rect 38013 4604 38025 4607
rect 31726 4576 38025 4604
rect 21416 4508 23336 4536
rect 21416 4496 21422 4508
rect 15194 4468 15200 4480
rect 11716 4440 15200 4468
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15746 4428 15752 4480
rect 15804 4468 15810 4480
rect 17494 4468 17500 4480
rect 15804 4440 17500 4468
rect 15804 4428 15810 4440
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17586 4428 17592 4480
rect 17644 4468 17650 4480
rect 19426 4468 19432 4480
rect 17644 4440 19432 4468
rect 17644 4428 17650 4440
rect 19426 4428 19432 4440
rect 19484 4428 19490 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 20622 4468 20628 4480
rect 20036 4440 20628 4468
rect 20036 4428 20042 4440
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 22741 4471 22799 4477
rect 22741 4468 22753 4471
rect 20772 4440 22753 4468
rect 20772 4428 20778 4440
rect 22741 4437 22753 4440
rect 22787 4437 22799 4471
rect 22741 4431 22799 4437
rect 23385 4471 23443 4477
rect 23385 4437 23397 4471
rect 23431 4468 23443 4471
rect 24118 4468 24124 4480
rect 23431 4440 24124 4468
rect 23431 4437 23443 4440
rect 23385 4431 23443 4437
rect 24118 4428 24124 4440
rect 24176 4428 24182 4480
rect 31113 4471 31171 4477
rect 31113 4437 31125 4471
rect 31159 4468 31171 4471
rect 31726 4468 31754 4576
rect 38013 4573 38025 4576
rect 38059 4573 38071 4607
rect 38013 4567 38071 4573
rect 38194 4468 38200 4480
rect 31159 4440 31754 4468
rect 38155 4440 38200 4468
rect 31159 4437 31171 4440
rect 31113 4431 31171 4437
rect 38194 4428 38200 4440
rect 38252 4428 38258 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 2409 4267 2467 4273
rect 2409 4233 2421 4267
rect 2455 4264 2467 4267
rect 2774 4264 2780 4276
rect 2455 4236 2780 4264
rect 2455 4233 2467 4236
rect 2409 4227 2467 4233
rect 2774 4224 2780 4236
rect 2832 4224 2838 4276
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 3878 4264 3884 4276
rect 3200 4236 3884 4264
rect 3200 4224 3206 4236
rect 3878 4224 3884 4236
rect 3936 4264 3942 4276
rect 9125 4267 9183 4273
rect 3936 4236 8708 4264
rect 3936 4224 3942 4236
rect 1670 4196 1676 4208
rect 1631 4168 1676 4196
rect 1670 4156 1676 4168
rect 1728 4156 1734 4208
rect 3053 4199 3111 4205
rect 3053 4165 3065 4199
rect 3099 4196 3111 4199
rect 3234 4196 3240 4208
rect 3099 4168 3240 4196
rect 3099 4165 3111 4168
rect 3053 4159 3111 4165
rect 3234 4156 3240 4168
rect 3292 4156 3298 4208
rect 3694 4156 3700 4208
rect 3752 4196 3758 4208
rect 3973 4199 4031 4205
rect 3973 4196 3985 4199
rect 3752 4168 3985 4196
rect 3752 4156 3758 4168
rect 3973 4165 3985 4168
rect 4019 4165 4031 4199
rect 8202 4196 8208 4208
rect 5198 4168 8208 4196
rect 3973 4159 4031 4165
rect 8202 4156 8208 4168
rect 8260 4156 8266 4208
rect 8680 4196 8708 4236
rect 9125 4233 9137 4267
rect 9171 4264 9183 4267
rect 9306 4264 9312 4276
rect 9171 4236 9312 4264
rect 9171 4233 9183 4236
rect 9125 4227 9183 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 9640 4236 12112 4264
rect 9640 4224 9646 4236
rect 8938 4196 8944 4208
rect 8680 4168 8944 4196
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 9950 4156 9956 4208
rect 10008 4196 10014 4208
rect 11422 4196 11428 4208
rect 10008 4168 11428 4196
rect 10008 4156 10014 4168
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1857 4131 1915 4137
rect 1857 4128 1869 4131
rect 900 4100 1869 4128
rect 900 4088 906 4100
rect 1857 4097 1869 4100
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 7745 4131 7803 4137
rect 7745 4097 7757 4131
rect 7791 4128 7803 4131
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 7791 4100 8401 4128
rect 7791 4097 7803 4100
rect 7745 4091 7803 4097
rect 8389 4097 8401 4100
rect 8435 4128 8447 4131
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8435 4100 9045 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 9033 4097 9045 4100
rect 9079 4128 9091 4131
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9079 4100 9689 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9677 4097 9689 4100
rect 9723 4128 9735 4131
rect 10321 4131 10379 4137
rect 10321 4128 10333 4131
rect 9723 4100 10333 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 10321 4097 10333 4100
rect 10367 4128 10379 4131
rect 10502 4128 10508 4140
rect 10367 4100 10508 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 2332 3992 2360 4091
rect 3694 4060 3700 4072
rect 3655 4032 3700 4060
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 6564 4060 6592 4091
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 10980 4137 11008 4168
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 12084 4196 12112 4236
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 14366 4264 14372 4276
rect 12216 4236 14372 4264
rect 12216 4224 12222 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 14642 4224 14648 4276
rect 14700 4264 14706 4276
rect 17034 4264 17040 4276
rect 14700 4236 17040 4264
rect 14700 4224 14706 4236
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 17276 4236 19334 4264
rect 17276 4224 17282 4236
rect 12526 4196 12532 4208
rect 12084 4168 12532 4196
rect 12526 4156 12532 4168
rect 12584 4156 12590 4208
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 17770 4196 17776 4208
rect 12768 4168 17776 4196
rect 12768 4156 12774 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 19306 4196 19334 4236
rect 19426 4224 19432 4276
rect 19484 4264 19490 4276
rect 31294 4264 31300 4276
rect 19484 4236 31300 4264
rect 19484 4224 19490 4236
rect 31294 4224 31300 4236
rect 31352 4224 31358 4276
rect 20714 4196 20720 4208
rect 18288 4168 18552 4196
rect 19306 4168 20720 4196
rect 18288 4156 18294 4168
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11974 4128 11980 4140
rect 11103 4100 11980 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12434 4128 12440 4140
rect 12299 4100 12440 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12860 4100 12909 4128
rect 12860 4088 12866 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4128 13047 4131
rect 13354 4128 13360 4140
rect 13035 4100 13360 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13722 4128 13728 4140
rect 13587 4100 13728 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13722 4088 13728 4100
rect 13780 4128 13786 4140
rect 13906 4128 13912 4140
rect 13780 4100 13912 4128
rect 13780 4088 13786 4100
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14185 4131 14243 4137
rect 14185 4128 14197 4131
rect 14148 4100 14197 4128
rect 14148 4088 14154 4100
rect 14185 4097 14197 4100
rect 14231 4097 14243 4131
rect 14185 4091 14243 4097
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14332 4100 14377 4128
rect 14332 4088 14338 4100
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14829 4131 14887 4137
rect 14829 4128 14841 4131
rect 14516 4100 14841 4128
rect 14516 4088 14522 4100
rect 14829 4097 14841 4100
rect 14875 4097 14887 4131
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 14829 4091 14887 4097
rect 15212 4100 15485 4128
rect 15102 4060 15108 4072
rect 3804 4032 5212 4060
rect 6564 4032 15108 4060
rect 2958 3992 2964 4004
rect 2332 3964 2964 3992
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3992 3295 3995
rect 3804 3992 3832 4032
rect 5184 4004 5212 4032
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 15212 4004 15240 4100
rect 15473 4097 15485 4100
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 15562 4088 15568 4140
rect 15620 4128 15626 4140
rect 15620 4100 15665 4128
rect 15620 4088 15626 4100
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15896 4100 16129 4128
rect 15896 4088 15902 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16666 4088 16672 4140
rect 16724 4128 16730 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16724 4100 16865 4128
rect 16724 4088 16730 4100
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 17494 4128 17500 4140
rect 17455 4100 17500 4128
rect 16853 4091 16911 4097
rect 17494 4088 17500 4100
rect 17552 4128 17558 4140
rect 17862 4128 17868 4140
rect 17552 4100 17868 4128
rect 17552 4088 17558 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 18414 4128 18420 4140
rect 18187 4100 18420 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 18524 4128 18552 4168
rect 20714 4156 20720 4168
rect 20772 4156 20778 4208
rect 23106 4156 23112 4208
rect 23164 4196 23170 4208
rect 23385 4199 23443 4205
rect 23385 4196 23397 4199
rect 23164 4168 23397 4196
rect 23164 4156 23170 4168
rect 23385 4165 23397 4168
rect 23431 4165 23443 4199
rect 23385 4159 23443 4165
rect 18785 4131 18843 4137
rect 18785 4128 18797 4131
rect 18524 4100 18797 4128
rect 18785 4097 18797 4100
rect 18831 4097 18843 4131
rect 19426 4128 19432 4140
rect 19387 4100 19432 4128
rect 18785 4091 18843 4097
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 20257 4131 20315 4137
rect 19576 4100 19621 4128
rect 19576 4088 19582 4100
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 20898 4128 20904 4140
rect 20859 4100 20904 4128
rect 20257 4091 20315 4097
rect 20272 4060 20300 4091
rect 20898 4088 20904 4100
rect 20956 4088 20962 4140
rect 21450 4088 21456 4140
rect 21508 4128 21514 4140
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21508 4126 21864 4128
rect 21928 4126 22017 4128
rect 21508 4100 22017 4126
rect 21508 4088 21514 4100
rect 21836 4098 21956 4100
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22462 4088 22468 4140
rect 22520 4128 22526 4140
rect 22649 4131 22707 4137
rect 22649 4128 22661 4131
rect 22520 4100 22661 4128
rect 22520 4088 22526 4100
rect 22649 4097 22661 4100
rect 22695 4097 22707 4131
rect 23290 4128 23296 4140
rect 23251 4100 23296 4128
rect 22649 4091 22707 4097
rect 23290 4088 23296 4100
rect 23348 4088 23354 4140
rect 24118 4128 24124 4140
rect 24079 4100 24124 4128
rect 24118 4088 24124 4100
rect 24176 4088 24182 4140
rect 38010 4128 38016 4140
rect 37971 4100 38016 4128
rect 38010 4088 38016 4100
rect 38068 4088 38074 4140
rect 22097 4063 22155 4069
rect 22097 4060 22109 4063
rect 15488 4032 20116 4060
rect 20272 4032 22109 4060
rect 3283 3964 3832 3992
rect 3283 3961 3295 3964
rect 3237 3955 3295 3961
rect 5166 3952 5172 4004
rect 5224 3952 5230 4004
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 6733 3995 6791 4001
rect 6733 3992 6745 3995
rect 6512 3964 6745 3992
rect 6512 3952 6518 3964
rect 6733 3961 6745 3964
rect 6779 3961 6791 3995
rect 6733 3955 6791 3961
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 8846 3992 8852 4004
rect 8527 3964 8852 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 10134 3992 10140 4004
rect 8956 3964 10140 3992
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 5350 3924 5356 3936
rect 3752 3896 5356 3924
rect 3752 3884 3758 3896
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5442 3884 5448 3936
rect 5500 3924 5506 3936
rect 7837 3927 7895 3933
rect 5500 3896 5545 3924
rect 5500 3884 5506 3896
rect 7837 3893 7849 3927
rect 7883 3924 7895 3927
rect 8956 3924 8984 3964
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 12066 3992 12072 4004
rect 10459 3964 12072 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12342 3992 12348 4004
rect 12303 3964 12348 3992
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 12986 3952 12992 4004
rect 13044 3992 13050 4004
rect 14458 3992 14464 4004
rect 13044 3964 14464 3992
rect 13044 3952 13050 3964
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 14550 3952 14556 4004
rect 14608 3992 14614 4004
rect 15194 3992 15200 4004
rect 14608 3964 15200 3992
rect 14608 3952 14614 3964
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 7883 3896 8984 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9398 3924 9404 3936
rect 9272 3896 9404 3924
rect 9272 3884 9278 3896
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9769 3927 9827 3933
rect 9769 3893 9781 3927
rect 9815 3924 9827 3927
rect 10226 3924 10232 3936
rect 9815 3896 10232 3924
rect 9815 3893 9827 3896
rect 9769 3887 9827 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 12158 3924 12164 3936
rect 10376 3896 12164 3924
rect 10376 3884 10382 3896
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13078 3924 13084 3936
rect 12492 3896 13084 3924
rect 12492 3884 12498 3896
rect 13078 3884 13084 3896
rect 13136 3884 13142 3936
rect 13630 3924 13636 3936
rect 13591 3896 13636 3924
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 14568 3924 14596 3952
rect 13780 3896 14596 3924
rect 13780 3884 13786 3896
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 14792 3896 14933 3924
rect 14792 3884 14798 3896
rect 14921 3893 14933 3896
rect 14967 3893 14979 3927
rect 14921 3887 14979 3893
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15488 3924 15516 4032
rect 15562 3952 15568 4004
rect 15620 3992 15626 4004
rect 16209 3995 16267 4001
rect 16209 3992 16221 3995
rect 15620 3964 16221 3992
rect 15620 3952 15626 3964
rect 16209 3961 16221 3964
rect 16255 3961 16267 3995
rect 16209 3955 16267 3961
rect 17310 3952 17316 4004
rect 17368 3992 17374 4004
rect 17589 3995 17647 4001
rect 17589 3992 17601 3995
rect 17368 3964 17601 3992
rect 17368 3952 17374 3964
rect 17589 3961 17601 3964
rect 17635 3961 17647 3995
rect 17589 3955 17647 3961
rect 17678 3952 17684 4004
rect 17736 3992 17742 4004
rect 18877 3995 18935 4001
rect 18877 3992 18889 3995
rect 17736 3964 18889 3992
rect 17736 3952 17742 3964
rect 18877 3961 18889 3964
rect 18923 3961 18935 3995
rect 19978 3992 19984 4004
rect 18877 3955 18935 3961
rect 18984 3964 19984 3992
rect 15160 3896 15516 3924
rect 15160 3884 15166 3896
rect 15930 3884 15936 3936
rect 15988 3924 15994 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 15988 3896 16957 3924
rect 15988 3884 15994 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18138 3924 18144 3936
rect 17828 3896 18144 3924
rect 17828 3884 17834 3896
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 18233 3927 18291 3933
rect 18233 3893 18245 3927
rect 18279 3924 18291 3927
rect 18322 3924 18328 3936
rect 18279 3896 18328 3924
rect 18279 3893 18291 3896
rect 18233 3887 18291 3893
rect 18322 3884 18328 3896
rect 18380 3884 18386 3936
rect 18414 3884 18420 3936
rect 18472 3924 18478 3936
rect 18984 3924 19012 3964
rect 19978 3952 19984 3964
rect 20036 3952 20042 4004
rect 20088 4001 20116 4032
rect 22097 4029 22109 4032
rect 22143 4029 22155 4063
rect 22097 4023 22155 4029
rect 20073 3995 20131 4001
rect 20073 3961 20085 3995
rect 20119 3961 20131 3995
rect 23014 3992 23020 4004
rect 20073 3955 20131 3961
rect 20180 3964 23020 3992
rect 18472 3896 19012 3924
rect 18472 3884 18478 3896
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 20180 3924 20208 3964
rect 23014 3952 23020 3964
rect 23072 3952 23078 4004
rect 20714 3924 20720 3936
rect 19208 3896 20208 3924
rect 20675 3896 20720 3924
rect 19208 3884 19214 3896
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 20990 3884 20996 3936
rect 21048 3924 21054 3936
rect 22741 3927 22799 3933
rect 22741 3924 22753 3927
rect 21048 3896 22753 3924
rect 21048 3884 21054 3896
rect 22741 3893 22753 3896
rect 22787 3893 22799 3927
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 22741 3887 22799 3893
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 37182 3884 37188 3936
rect 37240 3924 37246 3936
rect 38197 3927 38255 3933
rect 38197 3924 38209 3927
rect 37240 3896 38209 3924
rect 37240 3884 37246 3896
rect 38197 3893 38209 3896
rect 38243 3893 38255 3927
rect 38197 3887 38255 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 6733 3723 6791 3729
rect 6733 3720 6745 3723
rect 4028 3692 6745 3720
rect 4028 3680 4034 3692
rect 6733 3689 6745 3692
rect 6779 3689 6791 3723
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 6733 3683 6791 3689
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 9548 3692 10425 3720
rect 9548 3680 9554 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 11701 3723 11759 3729
rect 11701 3720 11713 3723
rect 10652 3692 11713 3720
rect 10652 3680 10658 3692
rect 11701 3689 11713 3692
rect 11747 3689 11759 3723
rect 11701 3683 11759 3689
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 12216 3692 12357 3720
rect 12216 3680 12222 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12618 3720 12624 3732
rect 12345 3683 12403 3689
rect 12452 3692 12624 3720
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 9769 3655 9827 3661
rect 9769 3652 9781 3655
rect 9732 3624 9781 3652
rect 9732 3612 9738 3624
rect 9769 3621 9781 3624
rect 9815 3621 9827 3655
rect 9769 3615 9827 3621
rect 11057 3655 11115 3661
rect 11057 3621 11069 3655
rect 11103 3652 11115 3655
rect 11330 3652 11336 3664
rect 11103 3624 11336 3652
rect 11103 3621 11115 3624
rect 11057 3615 11115 3621
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 11790 3612 11796 3664
rect 11848 3652 11854 3664
rect 12452 3652 12480 3692
rect 12618 3680 12624 3692
rect 12676 3720 12682 3732
rect 12986 3720 12992 3732
rect 12676 3692 12992 3720
rect 12676 3680 12682 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13228 3692 13645 3720
rect 13228 3680 13234 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 16574 3720 16580 3732
rect 16163 3692 16580 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 18046 3720 18052 3732
rect 18007 3692 18052 3720
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 18785 3723 18843 3729
rect 18785 3720 18797 3723
rect 18564 3692 18797 3720
rect 18564 3680 18570 3692
rect 18785 3689 18797 3692
rect 18831 3689 18843 3723
rect 18785 3683 18843 3689
rect 19150 3680 19156 3732
rect 19208 3720 19214 3732
rect 19886 3720 19892 3732
rect 19208 3692 19892 3720
rect 19208 3680 19214 3692
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 19996 3692 20484 3720
rect 11848 3624 12480 3652
rect 11848 3612 11854 3624
rect 14182 3612 14188 3664
rect 14240 3652 14246 3664
rect 18230 3652 18236 3664
rect 14240 3624 18236 3652
rect 14240 3612 14246 3624
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 19996 3652 20024 3692
rect 18616 3624 20024 3652
rect 20073 3655 20131 3661
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 1673 3587 1731 3593
rect 1673 3584 1685 3587
rect 1636 3556 1685 3584
rect 1636 3544 1642 3556
rect 1673 3553 1685 3556
rect 1719 3553 1731 3587
rect 1673 3547 1731 3553
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 3510 3584 3516 3596
rect 1995 3556 3516 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4614 3584 4620 3596
rect 4387 3556 4620 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 7190 3584 7196 3596
rect 4764 3556 7196 3584
rect 4764 3544 4770 3556
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 10778 3584 10784 3596
rect 9456 3556 10784 3584
rect 9456 3544 9462 3556
rect 10778 3544 10784 3556
rect 10836 3584 10842 3596
rect 10836 3556 12204 3584
rect 10836 3544 10842 3556
rect 4154 3516 4160 3528
rect 3082 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 5994 3516 6000 3528
rect 5750 3488 6000 3516
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6546 3516 6552 3528
rect 6507 3488 6552 3516
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 8294 3516 8300 3528
rect 7331 3488 8300 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 9122 3516 9128 3528
rect 8435 3488 9128 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 10226 3516 10232 3528
rect 9723 3488 10232 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 4617 3451 4675 3457
rect 3252 3420 3556 3448
rect 658 3340 664 3392
rect 716 3380 722 3392
rect 3252 3380 3280 3420
rect 716 3352 3280 3380
rect 716 3340 722 3352
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 3384 3352 3433 3380
rect 3384 3340 3390 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 3528 3380 3556 3420
rect 4617 3417 4629 3451
rect 4663 3448 4675 3451
rect 4706 3448 4712 3460
rect 4663 3420 4712 3448
rect 4663 3417 4675 3420
rect 4617 3411 4675 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 5920 3420 7512 3448
rect 5920 3380 5948 3420
rect 3528 3352 5948 3380
rect 6089 3383 6147 3389
rect 3421 3343 3479 3349
rect 6089 3349 6101 3383
rect 6135 3380 6147 3383
rect 7374 3380 7380 3392
rect 6135 3352 7380 3380
rect 6135 3349 6147 3352
rect 6089 3343 6147 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7484 3389 7512 3420
rect 9766 3408 9772 3460
rect 9824 3448 9830 3460
rect 10042 3448 10048 3460
rect 9824 3420 10048 3448
rect 9824 3408 9830 3420
rect 10042 3408 10048 3420
rect 10100 3448 10106 3460
rect 10336 3448 10364 3479
rect 10502 3476 10508 3528
rect 10560 3516 10566 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10560 3488 10977 3516
rect 10560 3476 10566 3488
rect 10965 3485 10977 3488
rect 11011 3516 11023 3519
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11011 3488 11621 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 11609 3485 11621 3488
rect 11655 3516 11667 3519
rect 11882 3516 11888 3528
rect 11655 3488 11888 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12176 3516 12204 3556
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 16850 3584 16856 3596
rect 12676 3556 16856 3584
rect 12676 3544 12682 3556
rect 16850 3544 16856 3556
rect 16908 3544 16914 3596
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17000 3556 17325 3584
rect 17000 3544 17006 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 18616 3584 18644 3624
rect 20073 3621 20085 3655
rect 20119 3621 20131 3655
rect 20073 3615 20131 3621
rect 20088 3584 20116 3615
rect 17828 3556 18644 3584
rect 18708 3556 20116 3584
rect 20456 3584 20484 3692
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 20809 3723 20867 3729
rect 20809 3720 20821 3723
rect 20680 3692 20821 3720
rect 20680 3680 20686 3692
rect 20809 3689 20821 3692
rect 20855 3689 20867 3723
rect 24578 3720 24584 3732
rect 24539 3692 24584 3720
rect 20809 3683 20867 3689
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 35802 3680 35808 3732
rect 35860 3720 35866 3732
rect 36725 3723 36783 3729
rect 36725 3720 36737 3723
rect 35860 3692 36737 3720
rect 35860 3680 35866 3692
rect 36725 3689 36737 3692
rect 36771 3689 36783 3723
rect 36725 3683 36783 3689
rect 21910 3612 21916 3664
rect 21968 3652 21974 3664
rect 21968 3624 31754 3652
rect 21968 3612 21974 3624
rect 22186 3584 22192 3596
rect 20456 3556 22192 3584
rect 17828 3544 17834 3556
rect 12245 3519 12303 3525
rect 12245 3516 12257 3519
rect 12176 3488 12257 3516
rect 12245 3485 12257 3488
rect 12291 3516 12303 3519
rect 12897 3519 12955 3525
rect 12291 3488 12848 3516
rect 12291 3485 12303 3488
rect 12245 3479 12303 3485
rect 10594 3448 10600 3460
rect 10100 3420 10600 3448
rect 10100 3408 10106 3420
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 12434 3448 12440 3460
rect 10928 3420 12440 3448
rect 10928 3408 10934 3420
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 12820 3448 12848 3488
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 12986 3516 12992 3528
rect 12943 3488 12992 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13136 3488 13553 3516
rect 13136 3476 13142 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14516 3488 14749 3516
rect 14516 3476 14522 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 14884 3488 14929 3516
rect 14884 3476 14890 3488
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15252 3488 15393 3516
rect 15252 3476 15258 3488
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15528 3488 16037 3516
rect 15528 3476 15534 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16025 3479 16083 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 17954 3516 17960 3528
rect 17915 3488 17960 3516
rect 16669 3479 16727 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18046 3476 18052 3528
rect 18104 3516 18110 3528
rect 18414 3516 18420 3528
rect 18104 3488 18420 3516
rect 18104 3476 18110 3488
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 18708 3525 18736 3556
rect 22186 3544 22192 3556
rect 22244 3544 22250 3596
rect 31726 3584 31754 3624
rect 35710 3612 35716 3664
rect 35768 3652 35774 3664
rect 37369 3655 37427 3661
rect 37369 3652 37381 3655
rect 35768 3624 37381 3652
rect 35768 3612 35774 3624
rect 37369 3621 37381 3624
rect 37415 3621 37427 3655
rect 37369 3615 37427 3621
rect 38289 3587 38347 3593
rect 38289 3584 38301 3587
rect 31726 3556 38301 3584
rect 38289 3553 38301 3556
rect 38335 3553 38347 3587
rect 38289 3547 38347 3553
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19300 3488 19441 3516
rect 19300 3476 19306 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20257 3479 20315 3485
rect 12820 3420 15608 3448
rect 7469 3383 7527 3389
rect 7469 3349 7481 3383
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 12618 3380 12624 3392
rect 7800 3352 12624 3380
rect 7800 3340 7806 3352
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12986 3380 12992 3392
rect 12947 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 15470 3380 15476 3392
rect 15431 3352 15476 3380
rect 15470 3340 15476 3352
rect 15528 3340 15534 3392
rect 15580 3380 15608 3420
rect 15654 3408 15660 3460
rect 15712 3448 15718 3460
rect 16761 3451 16819 3457
rect 16761 3448 16773 3451
rect 15712 3420 16773 3448
rect 15712 3408 15718 3420
rect 16761 3417 16773 3420
rect 16807 3417 16819 3451
rect 16761 3411 16819 3417
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 20272 3448 20300 3479
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20680 3488 20729 3516
rect 20680 3476 20686 3488
rect 20717 3485 20729 3488
rect 20763 3516 20775 3519
rect 21174 3516 21180 3528
rect 20763 3488 21180 3516
rect 20763 3485 20775 3488
rect 20717 3479 20775 3485
rect 21174 3476 21180 3488
rect 21232 3476 21238 3528
rect 21358 3516 21364 3528
rect 21319 3488 21364 3516
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 22002 3516 22008 3528
rect 21963 3488 22008 3516
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22833 3519 22891 3525
rect 22833 3516 22845 3519
rect 22336 3488 22845 3516
rect 22336 3476 22342 3488
rect 22833 3485 22845 3488
rect 22879 3485 22891 3519
rect 24026 3516 24032 3528
rect 23987 3488 24032 3516
rect 22833 3479 22891 3485
rect 24026 3476 24032 3488
rect 24084 3476 24090 3528
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 36909 3519 36967 3525
rect 36909 3485 36921 3519
rect 36955 3516 36967 3519
rect 37274 3516 37280 3528
rect 36955 3488 37280 3516
rect 36955 3485 36967 3488
rect 36909 3479 36967 3485
rect 16908 3420 20300 3448
rect 16908 3408 16914 3420
rect 21082 3408 21088 3460
rect 21140 3448 21146 3460
rect 24780 3448 24808 3479
rect 37274 3476 37280 3488
rect 37332 3476 37338 3528
rect 37553 3519 37611 3525
rect 37553 3485 37565 3519
rect 37599 3516 37611 3519
rect 39298 3516 39304 3528
rect 37599 3488 39304 3516
rect 37599 3485 37611 3488
rect 37553 3479 37611 3485
rect 39298 3476 39304 3488
rect 39356 3476 39362 3528
rect 21140 3420 24808 3448
rect 38105 3451 38163 3457
rect 21140 3408 21146 3420
rect 38105 3417 38117 3451
rect 38151 3448 38163 3451
rect 38286 3448 38292 3460
rect 38151 3420 38292 3448
rect 38151 3417 38163 3420
rect 38105 3411 38163 3417
rect 38286 3408 38292 3420
rect 38344 3408 38350 3460
rect 16574 3380 16580 3392
rect 15580 3352 16580 3380
rect 16574 3340 16580 3352
rect 16632 3340 16638 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 19242 3380 19248 3392
rect 17368 3352 19248 3380
rect 17368 3340 17374 3352
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 19521 3383 19579 3389
rect 19521 3349 19533 3383
rect 19567 3380 19579 3383
rect 19978 3380 19984 3392
rect 19567 3352 19984 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 21450 3380 21456 3392
rect 21411 3352 21456 3380
rect 21450 3340 21456 3352
rect 21508 3340 21514 3392
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21600 3352 21833 3380
rect 21600 3340 21606 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 22278 3380 22284 3392
rect 22239 3352 22284 3380
rect 21821 3343 21879 3349
rect 22278 3340 22284 3352
rect 22336 3340 22342 3392
rect 22646 3380 22652 3392
rect 22607 3352 22652 3380
rect 22646 3340 22652 3352
rect 22704 3340 22710 3392
rect 23845 3383 23903 3389
rect 23845 3349 23857 3383
rect 23891 3380 23903 3383
rect 23934 3380 23940 3392
rect 23891 3352 23940 3380
rect 23891 3349 23903 3352
rect 23845 3343 23903 3349
rect 23934 3340 23940 3352
rect 23992 3340 23998 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 3142 3176 3148 3188
rect 1872 3148 3148 3176
rect 1872 3117 1900 3148
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3329 3179 3387 3185
rect 3329 3145 3341 3179
rect 3375 3176 3387 3179
rect 3510 3176 3516 3188
rect 3375 3148 3516 3176
rect 3375 3145 3387 3148
rect 3329 3139 3387 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 6733 3179 6791 3185
rect 6733 3176 6745 3179
rect 3620 3148 6745 3176
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3077 1915 3111
rect 1857 3071 1915 3077
rect 1578 3040 1584 3052
rect 1539 3012 1584 3040
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 2958 3000 2964 3052
rect 3016 3000 3022 3052
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 3620 2972 3648 3148
rect 6733 3145 6745 3148
rect 6779 3145 6791 3179
rect 9858 3176 9864 3188
rect 9819 3148 9864 3176
rect 6733 3139 6791 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11146 3176 11152 3188
rect 10152 3148 11152 3176
rect 8202 3108 8208 3120
rect 5290 3080 8208 3108
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 9217 3111 9275 3117
rect 9217 3077 9229 3111
rect 9263 3108 9275 3111
rect 10152 3108 10180 3148
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12710 3176 12716 3188
rect 11256 3148 12716 3176
rect 10686 3108 10692 3120
rect 9263 3080 10180 3108
rect 10647 3080 10692 3108
rect 9263 3077 9275 3080
rect 9217 3071 9275 3077
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3752 3012 3801 3040
rect 3752 3000 3758 3012
rect 3789 3009 3801 3012
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 6546 3040 6552 3052
rect 5408 3012 6224 3040
rect 6507 3012 6552 3040
rect 5408 3000 5414 3012
rect 4062 2972 4068 2984
rect 2648 2944 3648 2972
rect 4023 2944 4068 2972
rect 2648 2932 2654 2944
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 5902 2972 5908 2984
rect 4212 2944 5908 2972
rect 4212 2932 4218 2944
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 6196 2972 6224 3012
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7282 3040 7288 3052
rect 7243 3012 7288 3040
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9398 3040 9404 3052
rect 9171 3012 9404 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 8036 2972 8064 3003
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9732 3012 9781 3040
rect 9732 3000 9738 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10376 3012 10517 3040
rect 10376 3000 10382 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 11146 2972 11152 2984
rect 6196 2944 7604 2972
rect 8036 2944 11152 2972
rect 7469 2907 7527 2913
rect 7469 2904 7481 2907
rect 3252 2876 3464 2904
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 3252 2836 3280 2876
rect 1360 2808 3280 2836
rect 3436 2836 3464 2876
rect 5092 2876 7481 2904
rect 5092 2836 5120 2876
rect 7469 2873 7481 2876
rect 7515 2873 7527 2907
rect 7576 2904 7604 2944
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11256 2904 11284 3148
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 12894 3176 12900 3188
rect 12855 3148 12900 3176
rect 12894 3136 12900 3148
rect 12952 3136 12958 3188
rect 13538 3176 13544 3188
rect 13499 3148 13544 3176
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 14734 3176 14740 3188
rect 13688 3148 14740 3176
rect 13688 3136 13694 3148
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 15473 3179 15531 3185
rect 15473 3176 15485 3179
rect 15436 3148 15485 3176
rect 15436 3136 15442 3148
rect 15473 3145 15485 3148
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 18141 3179 18199 3185
rect 18141 3145 18153 3179
rect 18187 3145 18199 3179
rect 18141 3139 18199 3145
rect 18156 3108 18184 3139
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19576 3148 19625 3176
rect 19576 3136 19582 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 19613 3139 19671 3145
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 21542 3176 21548 3188
rect 20220 3148 21548 3176
rect 20220 3136 20226 3148
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 22005 3179 22063 3185
rect 22005 3145 22017 3179
rect 22051 3176 22063 3179
rect 22830 3176 22836 3188
rect 22051 3148 22836 3176
rect 22051 3145 22063 3148
rect 22005 3139 22063 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 23290 3136 23296 3188
rect 23348 3176 23354 3188
rect 25777 3179 25835 3185
rect 25777 3176 25789 3179
rect 23348 3148 25789 3176
rect 23348 3136 23354 3148
rect 25777 3145 25789 3148
rect 25823 3145 25835 3179
rect 25777 3139 25835 3145
rect 25866 3136 25872 3188
rect 25924 3176 25930 3188
rect 27801 3179 27859 3185
rect 27801 3176 27813 3179
rect 25924 3148 27813 3176
rect 25924 3136 25930 3148
rect 27801 3145 27813 3148
rect 27847 3145 27859 3179
rect 27801 3139 27859 3145
rect 30374 3136 30380 3188
rect 30432 3176 30438 3188
rect 32953 3179 33011 3185
rect 32953 3176 32965 3179
rect 30432 3148 32965 3176
rect 30432 3136 30438 3148
rect 32953 3145 32965 3148
rect 32999 3145 33011 3179
rect 32953 3139 33011 3145
rect 34422 3136 34428 3188
rect 34480 3176 34486 3188
rect 36725 3179 36783 3185
rect 36725 3176 36737 3179
rect 34480 3148 36737 3176
rect 34480 3136 34486 3148
rect 36725 3145 36737 3148
rect 36771 3145 36783 3179
rect 36725 3139 36783 3145
rect 11716 3080 18184 3108
rect 11716 3049 11744 3080
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 18288 3080 21128 3108
rect 18288 3068 18294 3080
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 12342 3040 12348 3052
rect 11701 3003 11759 3009
rect 11808 3012 12348 3040
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 11808 2972 11836 3012
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12492 3012 12817 3040
rect 12492 3000 12498 3012
rect 12805 3009 12817 3012
rect 12851 3040 12863 3043
rect 13354 3040 13360 3052
rect 12851 3012 13360 3040
rect 12851 3009 12863 3012
rect 12805 3003 12863 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13630 3040 13636 3052
rect 13495 3012 13636 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 13780 3012 14105 3040
rect 13780 3000 13786 3012
rect 14093 3009 14105 3012
rect 14139 3040 14151 3043
rect 14550 3040 14556 3052
rect 14139 3012 14556 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 14734 3040 14740 3052
rect 14695 3012 14740 3040
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15838 3040 15844 3052
rect 15427 3012 15844 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 16114 3040 16120 3052
rect 16075 3012 16120 3040
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16298 3040 16304 3052
rect 16259 3012 16304 3040
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 18046 3040 18052 3052
rect 16899 3012 18052 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18322 3040 18328 3052
rect 18283 3012 18328 3040
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 18966 3040 18972 3052
rect 18927 3012 18972 3040
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19150 3000 19156 3052
rect 19208 3040 19214 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19208 3012 19441 3040
rect 19208 3000 19214 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19429 3003 19487 3009
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20036 3012 20361 3040
rect 20036 3000 20042 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20990 3040 20996 3052
rect 20951 3012 20996 3040
rect 20349 3003 20407 3009
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 11480 2944 11836 2972
rect 11480 2932 11486 2944
rect 12618 2932 12624 2984
rect 12676 2972 12682 2984
rect 21100 2972 21128 3080
rect 21450 3068 21456 3120
rect 21508 3108 21514 3120
rect 24949 3111 25007 3117
rect 21508 3080 23520 3108
rect 21508 3068 21514 3080
rect 21910 3000 21916 3052
rect 21968 3040 21974 3052
rect 23492 3049 23520 3080
rect 24949 3077 24961 3111
rect 24995 3108 25007 3111
rect 28810 3108 28816 3120
rect 24995 3080 28816 3108
rect 24995 3077 25007 3080
rect 24949 3071 25007 3077
rect 28810 3068 28816 3080
rect 28868 3068 28874 3120
rect 22189 3043 22247 3049
rect 22189 3040 22201 3043
rect 21968 3012 22201 3040
rect 21968 3000 21974 3012
rect 22189 3009 22201 3012
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23934 3040 23940 3052
rect 23895 3012 23940 3040
rect 23477 3003 23535 3009
rect 22848 2972 22876 3003
rect 23934 3000 23940 3012
rect 23992 3000 23998 3052
rect 25406 3040 25412 3052
rect 25367 3012 25412 3040
rect 25406 3000 25412 3012
rect 25464 3040 25470 3052
rect 25961 3043 26019 3049
rect 25961 3040 25973 3043
rect 25464 3012 25973 3040
rect 25464 3000 25470 3012
rect 25961 3009 25973 3012
rect 26007 3009 26019 3043
rect 26602 3040 26608 3052
rect 26563 3012 26608 3040
rect 25961 3003 26019 3009
rect 26602 3000 26608 3012
rect 26660 3000 26666 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 27985 3043 28043 3049
rect 27985 3040 27997 3043
rect 27764 3012 27997 3040
rect 27764 3000 27770 3012
rect 27985 3009 27997 3012
rect 28031 3009 28043 3043
rect 27985 3003 28043 3009
rect 32858 3000 32864 3052
rect 32916 3040 32922 3052
rect 33137 3043 33195 3049
rect 33137 3040 33149 3043
rect 32916 3012 33149 3040
rect 32916 3000 32922 3012
rect 33137 3009 33149 3012
rect 33183 3009 33195 3043
rect 36906 3040 36912 3052
rect 36867 3012 36912 3040
rect 33137 3003 33195 3009
rect 36906 3000 36912 3012
rect 36964 3000 36970 3052
rect 37550 3000 37556 3052
rect 37608 3040 37614 3052
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37608 3012 38025 3040
rect 37608 3000 37614 3012
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 12676 2944 20852 2972
rect 21100 2944 22876 2972
rect 12676 2932 12682 2944
rect 11698 2904 11704 2916
rect 7576 2876 11284 2904
rect 11348 2876 11704 2904
rect 7469 2867 7527 2873
rect 5534 2836 5540 2848
rect 3436 2808 5120 2836
rect 5495 2808 5540 2836
rect 1360 2796 1366 2808
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 8202 2836 8208 2848
rect 8163 2808 8208 2836
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 11348 2836 11376 2876
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 12710 2864 12716 2916
rect 12768 2904 12774 2916
rect 14829 2907 14887 2913
rect 14829 2904 14841 2907
rect 12768 2876 14841 2904
rect 12768 2864 12774 2876
rect 14829 2873 14841 2876
rect 14875 2873 14887 2907
rect 14829 2867 14887 2873
rect 16850 2864 16856 2916
rect 16908 2904 16914 2916
rect 20824 2913 20852 2944
rect 18785 2907 18843 2913
rect 18785 2904 18797 2907
rect 16908 2876 18797 2904
rect 16908 2864 16914 2876
rect 18785 2873 18797 2876
rect 18831 2873 18843 2907
rect 20165 2907 20223 2913
rect 20165 2904 20177 2907
rect 18785 2867 18843 2873
rect 18892 2876 20177 2904
rect 8444 2808 11376 2836
rect 8444 2796 8450 2808
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 11885 2839 11943 2845
rect 11885 2836 11897 2839
rect 11664 2808 11897 2836
rect 11664 2796 11670 2808
rect 11885 2805 11897 2808
rect 11931 2805 11943 2839
rect 11885 2799 11943 2805
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 13630 2836 13636 2848
rect 12032 2808 13636 2836
rect 12032 2796 12038 2808
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 14185 2839 14243 2845
rect 14185 2836 14197 2839
rect 13872 2808 14197 2836
rect 13872 2796 13878 2808
rect 14185 2805 14197 2808
rect 14231 2805 14243 2839
rect 14185 2799 14243 2805
rect 16758 2796 16764 2848
rect 16816 2836 16822 2848
rect 17037 2839 17095 2845
rect 17037 2836 17049 2839
rect 16816 2808 17049 2836
rect 16816 2796 16822 2808
rect 17037 2805 17049 2808
rect 17083 2805 17095 2839
rect 17037 2799 17095 2805
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 18892 2836 18920 2876
rect 20165 2873 20177 2876
rect 20211 2873 20223 2907
rect 20165 2867 20223 2873
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2873 20867 2907
rect 20809 2867 20867 2873
rect 20898 2864 20904 2916
rect 20956 2904 20962 2916
rect 22186 2904 22192 2916
rect 20956 2876 22192 2904
rect 20956 2864 20962 2876
rect 22186 2864 22192 2876
rect 22244 2904 22250 2916
rect 23198 2904 23204 2916
rect 22244 2876 23204 2904
rect 22244 2864 22250 2876
rect 23198 2864 23204 2876
rect 23256 2864 23262 2916
rect 26421 2907 26479 2913
rect 26421 2873 26433 2907
rect 26467 2904 26479 2907
rect 28902 2904 28908 2916
rect 26467 2876 28908 2904
rect 26467 2873 26479 2876
rect 26421 2867 26479 2873
rect 28902 2864 28908 2876
rect 28960 2864 28966 2916
rect 17552 2808 18920 2836
rect 17552 2796 17558 2808
rect 19058 2796 19064 2848
rect 19116 2836 19122 2848
rect 22649 2839 22707 2845
rect 22649 2836 22661 2839
rect 19116 2808 22661 2836
rect 19116 2796 19122 2808
rect 22649 2805 22661 2808
rect 22695 2805 22707 2839
rect 23290 2836 23296 2848
rect 23251 2808 23296 2836
rect 22649 2799 22707 2805
rect 23290 2796 23296 2808
rect 23348 2796 23354 2848
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23900 2808 24133 2836
rect 23900 2796 23906 2808
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 25038 2836 25044 2848
rect 24999 2808 25044 2836
rect 24121 2799 24179 2805
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 38010 2796 38016 2848
rect 38068 2836 38074 2848
rect 38197 2839 38255 2845
rect 38197 2836 38209 2839
rect 38068 2808 38209 2836
rect 38068 2796 38074 2808
rect 38197 2805 38209 2808
rect 38243 2805 38255 2839
rect 38197 2799 38255 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 3200 2604 3341 2632
rect 3200 2592 3206 2604
rect 3329 2601 3341 2604
rect 3375 2632 3387 2635
rect 4062 2632 4068 2644
rect 3375 2604 4068 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 5718 2632 5724 2644
rect 4448 2604 5724 2632
rect 4448 2564 4476 2604
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 12710 2632 12716 2644
rect 6886 2604 11928 2632
rect 4614 2564 4620 2576
rect 3896 2536 4476 2564
rect 4575 2536 4620 2564
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 3896 2496 3924 2536
rect 4614 2524 4620 2536
rect 4672 2524 4678 2576
rect 5258 2564 5264 2576
rect 5219 2536 5264 2564
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 4632 2496 4660 2524
rect 1903 2468 3924 2496
rect 3988 2468 4660 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 3988 2437 4016 2468
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 5721 2431 5779 2437
rect 3973 2391 4031 2397
rect 4632 2400 5212 2428
rect 4632 2360 4660 2400
rect 5074 2360 5080 2372
rect 3082 2332 4660 2360
rect 5035 2332 5080 2360
rect 5074 2320 5080 2332
rect 5132 2320 5138 2372
rect 5184 2360 5212 2400
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 6886 2428 6914 2604
rect 10870 2564 10876 2576
rect 7208 2536 10876 2564
rect 7208 2437 7236 2536
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 10962 2496 10968 2508
rect 7944 2468 10968 2496
rect 7944 2437 7972 2468
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 11790 2456 11796 2508
rect 11848 2456 11854 2508
rect 5767 2400 6914 2428
rect 7193 2431 7251 2437
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 9122 2428 9128 2440
rect 9083 2400 9128 2428
rect 7929 2391 7987 2397
rect 9122 2388 9128 2400
rect 9180 2388 9186 2440
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9272 2400 9317 2428
rect 9272 2388 9278 2400
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 10042 2428 10048 2440
rect 10003 2400 10048 2428
rect 9769 2391 9827 2397
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2428 11759 2431
rect 11808 2428 11836 2456
rect 11747 2400 11836 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 5184 2332 11805 2360
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11900 2360 11928 2604
rect 12360 2604 12716 2632
rect 12360 2437 12388 2604
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 14458 2632 14464 2644
rect 14108 2604 14464 2632
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 13722 2564 13728 2576
rect 12492 2536 13728 2564
rect 12492 2524 12498 2536
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 14108 2496 14136 2604
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 16853 2635 16911 2641
rect 16853 2601 16865 2635
rect 16899 2632 16911 2635
rect 19150 2632 19156 2644
rect 16899 2604 19156 2632
rect 16899 2601 16911 2604
rect 16853 2595 16911 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 19242 2592 19248 2644
rect 19300 2632 19306 2644
rect 19426 2632 19432 2644
rect 19300 2592 19334 2632
rect 19387 2604 19432 2632
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 25869 2635 25927 2641
rect 25869 2601 25881 2635
rect 25915 2632 25927 2635
rect 26142 2632 26148 2644
rect 25915 2604 26148 2632
rect 25915 2601 25927 2604
rect 25869 2595 25927 2601
rect 26142 2592 26148 2604
rect 26200 2592 26206 2644
rect 28276 2604 31248 2632
rect 18874 2564 18880 2576
rect 12584 2468 14136 2496
rect 14292 2536 18880 2564
rect 12584 2456 12590 2468
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12618 2428 12624 2440
rect 12492 2400 12624 2428
rect 12492 2388 12498 2400
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 14292 2437 14320 2536
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 19306 2564 19334 2592
rect 21082 2564 21088 2576
rect 19306 2536 21088 2564
rect 21082 2524 21088 2536
rect 21140 2524 21146 2576
rect 22281 2567 22339 2573
rect 22281 2533 22293 2567
rect 22327 2564 22339 2567
rect 24854 2564 24860 2576
rect 22327 2536 24860 2564
rect 22327 2533 22339 2536
rect 22281 2527 22339 2533
rect 24854 2524 24860 2536
rect 24912 2524 24918 2576
rect 25130 2524 25136 2576
rect 25188 2564 25194 2576
rect 27433 2567 27491 2573
rect 27433 2564 27445 2567
rect 25188 2536 27445 2564
rect 25188 2524 25194 2536
rect 27433 2533 27445 2536
rect 27479 2533 27491 2567
rect 27433 2527 27491 2533
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 19334 2496 19340 2508
rect 17819 2468 19340 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 20346 2496 20352 2508
rect 20307 2468 20352 2496
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22244 2468 24716 2496
rect 22244 2456 22250 2468
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 12860 2400 13553 2428
rect 12860 2388 12866 2400
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 14921 2391 14979 2397
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 16850 2360 16856 2372
rect 11900 2332 16856 2360
rect 11793 2323 11851 2329
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 17052 2360 17080 2391
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 18748 2400 19625 2428
rect 18748 2388 18754 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 20036 2400 20085 2428
rect 20036 2388 20042 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 21542 2388 21548 2440
rect 21600 2428 21606 2440
rect 23290 2428 23296 2440
rect 21600 2400 22232 2428
rect 23251 2400 23296 2428
rect 21600 2388 21606 2400
rect 20438 2360 20444 2372
rect 17052 2332 20444 2360
rect 20438 2320 20444 2332
rect 20496 2320 20502 2372
rect 21266 2320 21272 2372
rect 21324 2360 21330 2372
rect 22097 2363 22155 2369
rect 22097 2360 22109 2363
rect 21324 2332 22109 2360
rect 21324 2320 21330 2332
rect 22097 2329 22109 2332
rect 22143 2329 22155 2363
rect 22204 2360 22232 2400
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24688 2428 24716 2468
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 28276 2496 28304 2604
rect 30745 2567 30803 2573
rect 30745 2564 30757 2567
rect 24820 2468 28304 2496
rect 28368 2536 30757 2564
rect 24820 2456 24826 2468
rect 24857 2431 24915 2437
rect 24857 2428 24869 2431
rect 24688 2400 24869 2428
rect 24581 2391 24639 2397
rect 24857 2397 24869 2400
rect 24903 2397 24915 2431
rect 24857 2391 24915 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25832 2400 26065 2428
rect 25832 2388 25838 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 28368 2428 28396 2536
rect 30745 2533 30757 2536
rect 30791 2564 30803 2567
rect 31220 2564 31248 2604
rect 34790 2592 34796 2644
rect 34848 2632 34854 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 34848 2604 35081 2632
rect 34848 2592 34854 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 35897 2567 35955 2573
rect 35897 2564 35909 2567
rect 30791 2536 31156 2564
rect 31220 2536 35909 2564
rect 30791 2533 30803 2536
rect 30745 2527 30803 2533
rect 30190 2456 30196 2508
rect 30248 2496 30254 2508
rect 30248 2468 30328 2496
rect 30248 2456 30254 2468
rect 26053 2391 26111 2397
rect 26206 2400 28396 2428
rect 26206 2360 26234 2400
rect 28442 2388 28448 2440
rect 28500 2428 28506 2440
rect 29914 2428 29920 2440
rect 28500 2400 28545 2428
rect 29875 2400 29920 2428
rect 28500 2388 28506 2400
rect 29914 2388 29920 2400
rect 29972 2388 29978 2440
rect 30300 2437 30328 2468
rect 31128 2437 31156 2536
rect 35897 2533 35909 2536
rect 35943 2533 35955 2567
rect 35897 2527 35955 2533
rect 37642 2496 37648 2508
rect 36648 2468 37648 2496
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2397 30343 2431
rect 30285 2391 30343 2397
rect 31113 2431 31171 2437
rect 31113 2397 31125 2431
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 33594 2428 33600 2440
rect 33555 2400 33600 2428
rect 32309 2391 32367 2397
rect 22204 2332 26234 2360
rect 22097 2323 22155 2329
rect 26418 2320 26424 2372
rect 26476 2360 26482 2372
rect 27249 2363 27307 2369
rect 27249 2360 27261 2363
rect 26476 2332 27261 2360
rect 26476 2320 26482 2332
rect 27249 2329 27261 2332
rect 27295 2329 27307 2363
rect 27249 2323 27307 2329
rect 28902 2320 28908 2372
rect 28960 2360 28966 2372
rect 32324 2360 32352 2391
rect 33594 2388 33600 2400
rect 33652 2388 33658 2440
rect 36648 2437 36676 2468
rect 37642 2456 37648 2468
rect 37700 2456 37706 2508
rect 36633 2431 36691 2437
rect 36633 2397 36645 2431
rect 36679 2397 36691 2431
rect 36633 2391 36691 2397
rect 37366 2388 37372 2440
rect 37424 2428 37430 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 37424 2400 37473 2428
rect 37424 2388 37430 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37734 2428 37740 2440
rect 37695 2400 37740 2428
rect 37461 2391 37519 2397
rect 37734 2388 37740 2400
rect 37792 2388 37798 2440
rect 28960 2332 32352 2360
rect 28960 2320 28966 2332
rect 34790 2320 34796 2372
rect 34848 2360 34854 2372
rect 34977 2363 35035 2369
rect 34977 2360 34989 2363
rect 34848 2332 34989 2360
rect 34848 2320 34854 2332
rect 34977 2329 34989 2332
rect 35023 2329 35035 2363
rect 34977 2323 35035 2329
rect 35434 2320 35440 2372
rect 35492 2360 35498 2372
rect 35713 2363 35771 2369
rect 35713 2360 35725 2363
rect 35492 2332 35725 2360
rect 35492 2320 35498 2332
rect 35713 2329 35725 2332
rect 35759 2329 35771 2363
rect 35713 2323 35771 2329
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3936 2264 4169 2292
rect 3936 2252 3942 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5868 2264 5917 2292
rect 5868 2252 5874 2264
rect 5905 2261 5917 2264
rect 5951 2261 5963 2295
rect 6546 2292 6552 2304
rect 6507 2264 6552 2292
rect 5905 2255 5963 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 8110 2292 8116 2304
rect 8071 2264 8116 2292
rect 7377 2255 7435 2261
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 12158 2292 12164 2304
rect 11204 2264 12164 2292
rect 11204 2252 11210 2264
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12308 2264 12541 2292
rect 12308 2252 12314 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 13630 2292 13636 2304
rect 13591 2264 13636 2292
rect 12529 2255 12587 2261
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 14366 2292 14372 2304
rect 14327 2264 14372 2292
rect 14366 2252 14372 2264
rect 14424 2252 14430 2304
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 20806 2292 20812 2304
rect 14516 2264 20812 2292
rect 14516 2252 14522 2264
rect 20806 2252 20812 2264
rect 20864 2252 20870 2304
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23477 2295 23535 2301
rect 23477 2292 23489 2295
rect 23256 2264 23489 2292
rect 23256 2252 23262 2264
rect 23477 2261 23489 2264
rect 23523 2261 23535 2295
rect 23477 2255 23535 2261
rect 28350 2252 28356 2304
rect 28408 2292 28414 2304
rect 28629 2295 28687 2301
rect 28629 2292 28641 2295
rect 28408 2264 28641 2292
rect 28408 2252 28414 2264
rect 28629 2261 28641 2264
rect 28675 2261 28687 2295
rect 28629 2255 28687 2261
rect 29730 2252 29736 2304
rect 29788 2292 29794 2304
rect 29788 2264 29833 2292
rect 29788 2252 29794 2264
rect 30374 2252 30380 2304
rect 30432 2292 30438 2304
rect 30432 2264 30477 2292
rect 30432 2252 30438 2264
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 31297 2295 31355 2301
rect 31297 2292 31309 2295
rect 30984 2264 31309 2292
rect 30984 2252 30990 2264
rect 31297 2261 31309 2264
rect 31343 2261 31355 2295
rect 31297 2255 31355 2261
rect 32214 2252 32220 2304
rect 32272 2292 32278 2304
rect 32493 2295 32551 2301
rect 32493 2292 32505 2295
rect 32272 2264 32505 2292
rect 32272 2252 32278 2264
rect 32493 2261 32505 2264
rect 32539 2261 32551 2295
rect 32493 2255 32551 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 33560 2264 33793 2292
rect 33560 2252 33566 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 36722 2252 36728 2304
rect 36780 2292 36786 2304
rect 36817 2295 36875 2301
rect 36817 2292 36829 2295
rect 36780 2264 36829 2292
rect 36780 2252 36786 2264
rect 36817 2261 36829 2264
rect 36863 2261 36875 2295
rect 36817 2255 36875 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 6270 2048 6276 2100
rect 6328 2088 6334 2100
rect 9950 2088 9956 2100
rect 6328 2060 9956 2088
rect 6328 2048 6334 2060
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 10042 2048 10048 2100
rect 10100 2088 10106 2100
rect 10100 2060 12664 2088
rect 10100 2048 10106 2060
rect 3418 1980 3424 2032
rect 3476 2020 3482 2032
rect 12526 2020 12532 2032
rect 3476 1992 12532 2020
rect 3476 1980 3482 1992
rect 12526 1980 12532 1992
rect 12584 1980 12590 2032
rect 12636 2020 12664 2060
rect 12710 2048 12716 2100
rect 12768 2088 12774 2100
rect 20162 2088 20168 2100
rect 12768 2060 20168 2088
rect 12768 2048 12774 2060
rect 20162 2048 20168 2060
rect 20220 2048 20226 2100
rect 28442 2048 28448 2100
rect 28500 2088 28506 2100
rect 30742 2088 30748 2100
rect 28500 2060 30748 2088
rect 28500 2048 28506 2060
rect 30742 2048 30748 2060
rect 30800 2048 30806 2100
rect 17770 2020 17776 2032
rect 12636 1992 17776 2020
rect 17770 1980 17776 1992
rect 17828 1980 17834 2032
rect 19058 1980 19064 2032
rect 19116 2020 19122 2032
rect 20070 2020 20076 2032
rect 19116 1992 20076 2020
rect 19116 1980 19122 1992
rect 20070 1980 20076 1992
rect 20128 1980 20134 2032
rect 28810 1980 28816 2032
rect 28868 2020 28874 2032
rect 37734 2020 37740 2032
rect 28868 1992 37740 2020
rect 28868 1980 28874 1992
rect 37734 1980 37740 1992
rect 37792 1980 37798 2032
rect 3326 1912 3332 1964
rect 3384 1952 3390 1964
rect 5350 1952 5356 1964
rect 3384 1924 5356 1952
rect 3384 1912 3390 1924
rect 5350 1912 5356 1924
rect 5408 1952 5414 1964
rect 17218 1952 17224 1964
rect 5408 1924 17224 1952
rect 5408 1912 5414 1924
rect 17218 1912 17224 1924
rect 17276 1912 17282 1964
rect 9122 1844 9128 1896
rect 9180 1884 9186 1896
rect 22646 1884 22652 1896
rect 9180 1856 22652 1884
rect 9180 1844 9186 1856
rect 22646 1844 22652 1856
rect 22704 1844 22710 1896
rect 5994 1776 6000 1828
rect 6052 1816 6058 1828
rect 22738 1816 22744 1828
rect 6052 1788 22744 1816
rect 6052 1776 6058 1788
rect 22738 1776 22744 1788
rect 22796 1776 22802 1828
rect 6638 1708 6644 1760
rect 6696 1748 6702 1760
rect 22094 1748 22100 1760
rect 6696 1720 22100 1748
rect 6696 1708 6702 1720
rect 22094 1708 22100 1720
rect 22152 1708 22158 1760
rect 6546 1640 6552 1692
rect 6604 1680 6610 1692
rect 6604 1652 6914 1680
rect 6604 1640 6610 1652
rect 6886 1612 6914 1652
rect 9950 1640 9956 1692
rect 10008 1680 10014 1692
rect 17126 1680 17132 1692
rect 10008 1652 17132 1680
rect 10008 1640 10014 1652
rect 17126 1640 17132 1652
rect 17184 1640 17190 1692
rect 13262 1612 13268 1624
rect 6886 1584 13268 1612
rect 13262 1572 13268 1584
rect 13320 1572 13326 1624
rect 17218 1572 17224 1624
rect 17276 1612 17282 1624
rect 23750 1612 23756 1624
rect 17276 1584 23756 1612
rect 17276 1572 17282 1584
rect 23750 1572 23756 1584
rect 23808 1572 23814 1624
rect 7558 1504 7564 1556
rect 7616 1544 7622 1556
rect 13630 1544 13636 1556
rect 7616 1516 13636 1544
rect 7616 1504 7622 1516
rect 13630 1504 13636 1516
rect 13688 1504 13694 1556
rect 15562 1544 15568 1556
rect 14016 1516 15568 1544
rect 8018 1436 8024 1488
rect 8076 1476 8082 1488
rect 14016 1476 14044 1516
rect 15562 1504 15568 1516
rect 15620 1504 15626 1556
rect 8076 1448 14044 1476
rect 8076 1436 8082 1448
rect 15194 1436 15200 1488
rect 15252 1476 15258 1488
rect 26602 1476 26608 1488
rect 15252 1448 26608 1476
rect 15252 1436 15258 1448
rect 26602 1436 26608 1448
rect 26660 1436 26666 1488
rect 5902 1368 5908 1420
rect 5960 1408 5966 1420
rect 14366 1408 14372 1420
rect 5960 1380 14372 1408
rect 5960 1368 5966 1380
rect 14366 1368 14372 1380
rect 14424 1368 14430 1420
rect 28994 1368 29000 1420
rect 29052 1408 29058 1420
rect 29914 1408 29920 1420
rect 29052 1380 29920 1408
rect 29052 1368 29058 1380
rect 29914 1368 29920 1380
rect 29972 1368 29978 1420
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 8202 1340 8208 1352
rect 72 1312 8208 1340
rect 72 1300 78 1312
rect 8202 1300 8208 1312
rect 8260 1300 8266 1352
rect 9030 1300 9036 1352
rect 9088 1340 9094 1352
rect 20714 1340 20720 1352
rect 9088 1312 20720 1340
rect 9088 1300 9094 1312
rect 20714 1300 20720 1312
rect 20772 1300 20778 1352
rect 5534 1232 5540 1284
rect 5592 1272 5598 1284
rect 17954 1272 17960 1284
rect 5592 1244 17960 1272
rect 5592 1232 5598 1244
rect 17954 1232 17960 1244
rect 18012 1232 18018 1284
rect 12894 1164 12900 1216
rect 12952 1204 12958 1216
rect 17310 1204 17316 1216
rect 12952 1176 17316 1204
rect 12952 1164 12958 1176
rect 17310 1164 17316 1176
rect 17368 1164 17374 1216
rect 3510 756 3516 808
rect 3568 796 3574 808
rect 8110 796 8116 808
rect 3568 768 8116 796
rect 3568 756 3574 768
rect 8110 756 8116 768
rect 8168 756 8174 808
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16764 37408 16816 37460
rect 22744 37408 22796 37460
rect 32220 37408 32272 37460
rect 20168 37340 20220 37392
rect 2872 37272 2924 37324
rect 10324 37315 10376 37324
rect 1952 37204 2004 37256
rect 2964 37204 3016 37256
rect 10324 37281 10333 37315
rect 10333 37281 10367 37315
rect 10367 37281 10376 37315
rect 10324 37272 10376 37281
rect 14832 37272 14884 37324
rect 20628 37315 20680 37324
rect 20628 37281 20637 37315
rect 20637 37281 20671 37315
rect 20671 37281 20680 37315
rect 20628 37272 20680 37281
rect 22560 37272 22612 37324
rect 30932 37315 30984 37324
rect 30932 37281 30941 37315
rect 30941 37281 30975 37315
rect 30975 37281 30984 37315
rect 30932 37272 30984 37281
rect 34152 37272 34204 37324
rect 5724 37204 5776 37256
rect 5816 37204 5868 37256
rect 7104 37204 7156 37256
rect 9128 37247 9180 37256
rect 9128 37213 9137 37247
rect 9137 37213 9171 37247
rect 9171 37213 9180 37247
rect 9128 37204 9180 37213
rect 10600 37247 10652 37256
rect 10600 37213 10609 37247
rect 10609 37213 10643 37247
rect 10643 37213 10652 37247
rect 10600 37204 10652 37213
rect 12992 37247 13044 37256
rect 2780 37068 2832 37120
rect 6828 37136 6880 37188
rect 4620 37068 4672 37120
rect 10784 37136 10836 37188
rect 12992 37213 13001 37247
rect 13001 37213 13035 37247
rect 13035 37213 13044 37247
rect 12992 37204 13044 37213
rect 13544 37204 13596 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 18052 37204 18104 37256
rect 20076 37204 20128 37256
rect 20904 37247 20956 37256
rect 20904 37213 20913 37247
rect 20913 37213 20947 37247
rect 20947 37213 20956 37247
rect 20904 37204 20956 37213
rect 24584 37247 24636 37256
rect 16120 37136 16172 37188
rect 16580 37136 16632 37188
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 25320 37247 25372 37256
rect 25320 37213 25329 37247
rect 25329 37213 25363 37247
rect 25363 37213 25372 37247
rect 25320 37204 25372 37213
rect 26240 37204 26292 37256
rect 27528 37204 27580 37256
rect 29736 37247 29788 37256
rect 26976 37136 27028 37188
rect 27068 37136 27120 37188
rect 8392 37068 8444 37120
rect 11612 37068 11664 37120
rect 12900 37068 12952 37120
rect 15016 37068 15068 37120
rect 17960 37068 18012 37120
rect 19984 37068 20036 37120
rect 24492 37068 24544 37120
rect 25136 37068 25188 37120
rect 26424 37068 26476 37120
rect 27712 37136 27764 37188
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 31208 37247 31260 37256
rect 31208 37213 31217 37247
rect 31217 37213 31251 37247
rect 31251 37213 31260 37247
rect 31208 37204 31260 37213
rect 33048 37247 33100 37256
rect 33048 37213 33057 37247
rect 33057 37213 33091 37247
rect 33091 37213 33100 37247
rect 33048 37204 33100 37213
rect 33784 37247 33836 37256
rect 33784 37213 33793 37247
rect 33793 37213 33827 37247
rect 33827 37213 33836 37247
rect 33784 37204 33836 37213
rect 36084 37204 36136 37256
rect 36728 37204 36780 37256
rect 28632 37111 28684 37120
rect 28632 37077 28641 37111
rect 28641 37077 28675 37111
rect 28675 37077 28684 37111
rect 28632 37068 28684 37077
rect 28724 37068 28776 37120
rect 36544 37136 36596 37188
rect 29644 37068 29696 37120
rect 31760 37068 31812 37120
rect 33508 37068 33560 37120
rect 35900 37068 35952 37120
rect 37648 37111 37700 37120
rect 37648 37077 37657 37111
rect 37657 37077 37691 37111
rect 37691 37077 37700 37111
rect 37648 37068 37700 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1308 36864 1360 36916
rect 8760 36864 8812 36916
rect 11060 36864 11112 36916
rect 15200 36864 15252 36916
rect 3148 36839 3200 36848
rect 3148 36805 3157 36839
rect 3157 36805 3191 36839
rect 3191 36805 3200 36839
rect 3148 36796 3200 36805
rect 3884 36796 3936 36848
rect 15476 36796 15528 36848
rect 17408 36796 17460 36848
rect 19340 36864 19392 36916
rect 22100 36864 22152 36916
rect 23480 36907 23532 36916
rect 23480 36873 23489 36907
rect 23489 36873 23523 36907
rect 23523 36873 23532 36907
rect 23480 36864 23532 36873
rect 24768 36864 24820 36916
rect 28632 36864 28684 36916
rect 36820 36907 36872 36916
rect 36820 36873 36829 36907
rect 36829 36873 36863 36907
rect 36863 36873 36872 36907
rect 36820 36864 36872 36873
rect 2320 36728 2372 36780
rect 3056 36728 3108 36780
rect 6460 36728 6512 36780
rect 9036 36728 9088 36780
rect 11704 36771 11756 36780
rect 11704 36737 11713 36771
rect 11713 36737 11747 36771
rect 11747 36737 11756 36771
rect 11704 36728 11756 36737
rect 9220 36660 9272 36712
rect 9404 36703 9456 36712
rect 9404 36669 9413 36703
rect 9413 36669 9447 36703
rect 9447 36669 9456 36703
rect 9404 36660 9456 36669
rect 10968 36660 11020 36712
rect 19432 36771 19484 36780
rect 19432 36737 19441 36771
rect 19441 36737 19475 36771
rect 19475 36737 19484 36771
rect 19432 36728 19484 36737
rect 20904 36796 20956 36848
rect 21272 36728 21324 36780
rect 22376 36728 22428 36780
rect 23388 36728 23440 36780
rect 5356 36592 5408 36644
rect 10324 36592 10376 36644
rect 15844 36635 15896 36644
rect 15844 36601 15853 36635
rect 15853 36601 15887 36635
rect 15887 36601 15896 36635
rect 15844 36592 15896 36601
rect 3148 36524 3200 36576
rect 5540 36524 5592 36576
rect 10692 36524 10744 36576
rect 18696 36524 18748 36576
rect 21272 36592 21324 36644
rect 26976 36728 27028 36780
rect 29000 36728 29052 36780
rect 38016 36796 38068 36848
rect 35900 36771 35952 36780
rect 35900 36737 35909 36771
rect 35909 36737 35943 36771
rect 35943 36737 35952 36771
rect 35900 36728 35952 36737
rect 28724 36660 28776 36712
rect 33048 36660 33100 36712
rect 38660 36592 38712 36644
rect 28448 36524 28500 36576
rect 28540 36524 28592 36576
rect 37832 36524 37884 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1768 36363 1820 36372
rect 1768 36329 1777 36363
rect 1777 36329 1811 36363
rect 1811 36329 1820 36363
rect 1768 36320 1820 36329
rect 2320 36320 2372 36372
rect 5724 36320 5776 36372
rect 15844 36320 15896 36372
rect 21916 36320 21968 36372
rect 22376 36363 22428 36372
rect 22376 36329 22385 36363
rect 22385 36329 22419 36363
rect 22419 36329 22428 36363
rect 22376 36320 22428 36329
rect 24492 36320 24544 36372
rect 31208 36320 31260 36372
rect 37464 36363 37516 36372
rect 37464 36329 37473 36363
rect 37473 36329 37507 36363
rect 37507 36329 37516 36363
rect 37464 36320 37516 36329
rect 20 36184 72 36236
rect 3148 36184 3200 36236
rect 10968 36184 11020 36236
rect 28724 36184 28776 36236
rect 5540 36159 5592 36168
rect 5540 36125 5549 36159
rect 5549 36125 5583 36159
rect 5583 36125 5592 36159
rect 5540 36116 5592 36125
rect 12256 36116 12308 36168
rect 24492 36116 24544 36168
rect 2872 36048 2924 36100
rect 21548 36048 21600 36100
rect 33784 36116 33836 36168
rect 36176 36116 36228 36168
rect 29920 36048 29972 36100
rect 4068 35980 4120 36032
rect 36176 36023 36228 36032
rect 36176 35989 36185 36023
rect 36185 35989 36219 36023
rect 36219 35989 36228 36023
rect 36176 35980 36228 35989
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 12992 35776 13044 35828
rect 11888 35683 11940 35692
rect 11888 35649 11897 35683
rect 11897 35649 11931 35683
rect 11931 35649 11940 35683
rect 11888 35640 11940 35649
rect 39304 35708 39356 35760
rect 1584 35615 1636 35624
rect 1584 35581 1593 35615
rect 1593 35581 1627 35615
rect 1627 35581 1636 35615
rect 1584 35572 1636 35581
rect 2136 35572 2188 35624
rect 35532 35572 35584 35624
rect 34520 35436 34572 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 38292 35232 38344 35284
rect 11704 35164 11756 35216
rect 28080 35164 28132 35216
rect 10692 35071 10744 35080
rect 10692 35037 10701 35071
rect 10701 35037 10735 35071
rect 10735 35037 10744 35071
rect 10692 35028 10744 35037
rect 37280 35028 37332 35080
rect 13360 34892 13412 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 5816 34688 5868 34740
rect 29736 34688 29788 34740
rect 35900 34688 35952 34740
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 4068 34552 4120 34604
rect 11152 34620 11204 34672
rect 10784 34595 10836 34604
rect 10784 34561 10793 34595
rect 10793 34561 10827 34595
rect 10827 34561 10836 34595
rect 10784 34552 10836 34561
rect 27804 34595 27856 34604
rect 27804 34561 27813 34595
rect 27813 34561 27847 34595
rect 27847 34561 27856 34595
rect 27804 34552 27856 34561
rect 29000 34552 29052 34604
rect 37188 34484 37240 34536
rect 37740 34527 37792 34536
rect 37740 34493 37749 34527
rect 37749 34493 37783 34527
rect 37783 34493 37792 34527
rect 37740 34484 37792 34493
rect 10508 34348 10560 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 11888 34144 11940 34196
rect 27528 34187 27580 34196
rect 27528 34153 27537 34187
rect 27537 34153 27571 34187
rect 27571 34153 27580 34187
rect 27528 34144 27580 34153
rect 12532 33940 12584 33992
rect 22100 33940 22152 33992
rect 24768 33940 24820 33992
rect 26884 33940 26936 33992
rect 23572 33872 23624 33924
rect 23664 33804 23716 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 24584 33600 24636 33652
rect 112 33464 164 33516
rect 23664 33507 23716 33516
rect 20 33396 72 33448
rect 23664 33473 23673 33507
rect 23673 33473 23707 33507
rect 23707 33473 23716 33507
rect 23664 33464 23716 33473
rect 34520 33464 34572 33516
rect 38108 33507 38160 33516
rect 38108 33473 38117 33507
rect 38117 33473 38151 33507
rect 38151 33473 38160 33507
rect 38108 33464 38160 33473
rect 3424 33328 3476 33380
rect 20444 33328 20496 33380
rect 3976 33260 4028 33312
rect 21180 33260 21232 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 2872 33056 2924 33108
rect 1124 32988 1176 33040
rect 1492 32920 1544 32972
rect 2688 32852 2740 32904
rect 6828 32852 6880 32904
rect 36176 32852 36228 32904
rect 1768 32759 1820 32768
rect 1768 32725 1777 32759
rect 1777 32725 1811 32759
rect 1811 32725 1820 32759
rect 1768 32716 1820 32725
rect 2228 32759 2280 32768
rect 2228 32725 2237 32759
rect 2237 32725 2271 32759
rect 2271 32725 2280 32759
rect 2228 32716 2280 32725
rect 7196 32716 7248 32768
rect 25320 32716 25372 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 2228 32512 2280 32564
rect 22560 32512 22612 32564
rect 5356 32444 5408 32496
rect 27160 32444 27212 32496
rect 3056 32419 3108 32428
rect 3056 32385 3065 32419
rect 3065 32385 3099 32419
rect 3099 32385 3108 32419
rect 3056 32376 3108 32385
rect 3700 32419 3752 32428
rect 3700 32385 3709 32419
rect 3709 32385 3743 32419
rect 3743 32385 3752 32419
rect 3700 32376 3752 32385
rect 28540 32419 28592 32428
rect 28540 32385 28549 32419
rect 28549 32385 28583 32419
rect 28583 32385 28592 32419
rect 28540 32376 28592 32385
rect 33784 32376 33836 32428
rect 4988 32308 5040 32360
rect 37464 32351 37516 32360
rect 37464 32317 37473 32351
rect 37473 32317 37507 32351
rect 37507 32317 37516 32351
rect 37464 32308 37516 32317
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 1952 32172 2004 32224
rect 2688 32172 2740 32224
rect 6644 32172 6696 32224
rect 28540 32172 28592 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2964 32011 3016 32020
rect 2964 31977 2973 32011
rect 2973 31977 3007 32011
rect 3007 31977 3016 32011
rect 2964 31968 3016 31977
rect 35532 32011 35584 32020
rect 35532 31977 35541 32011
rect 35541 31977 35575 32011
rect 35575 31977 35584 32011
rect 35532 31968 35584 31977
rect 3792 31900 3844 31952
rect 848 31764 900 31816
rect 5632 31900 5684 31952
rect 5448 31832 5500 31884
rect 17960 31807 18012 31816
rect 17960 31773 17969 31807
rect 17969 31773 18003 31807
rect 18003 31773 18012 31807
rect 17960 31764 18012 31773
rect 19340 31764 19392 31816
rect 33876 31764 33928 31816
rect 37188 31764 37240 31816
rect 37556 31764 37608 31816
rect 5080 31696 5132 31748
rect 7288 31696 7340 31748
rect 11704 31628 11756 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4988 31467 5040 31476
rect 4988 31433 4997 31467
rect 4997 31433 5031 31467
rect 5031 31433 5040 31467
rect 4988 31424 5040 31433
rect 19432 31424 19484 31476
rect 756 31356 808 31408
rect 1400 31288 1452 31340
rect 3516 31288 3568 31340
rect 6552 31288 6604 31340
rect 12072 31288 12124 31340
rect 18696 31331 18748 31340
rect 18696 31297 18705 31331
rect 18705 31297 18739 31331
rect 18739 31297 18748 31331
rect 18696 31288 18748 31297
rect 20628 31331 20680 31340
rect 1860 31152 1912 31204
rect 9128 31220 9180 31272
rect 12440 31263 12492 31272
rect 12440 31229 12449 31263
rect 12449 31229 12483 31263
rect 12483 31229 12492 31263
rect 12440 31220 12492 31229
rect 17592 31220 17644 31272
rect 20628 31297 20637 31331
rect 20637 31297 20671 31331
rect 20671 31297 20680 31331
rect 20628 31288 20680 31297
rect 20352 31152 20404 31204
rect 1032 31084 1084 31136
rect 4712 31084 4764 31136
rect 10232 31084 10284 31136
rect 19984 31084 20036 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6552 30923 6604 30932
rect 6552 30889 6561 30923
rect 6561 30889 6595 30923
rect 6595 30889 6604 30923
rect 6552 30880 6604 30889
rect 12256 30880 12308 30932
rect 12716 30812 12768 30864
rect 1216 30744 1268 30796
rect 6736 30744 6788 30796
rect 11704 30787 11756 30796
rect 664 30676 716 30728
rect 3424 30719 3476 30728
rect 3424 30685 3433 30719
rect 3433 30685 3467 30719
rect 3467 30685 3476 30719
rect 3424 30676 3476 30685
rect 5080 30719 5132 30728
rect 5080 30685 5089 30719
rect 5089 30685 5123 30719
rect 5123 30685 5132 30719
rect 5080 30676 5132 30685
rect 5816 30719 5868 30728
rect 5816 30685 5825 30719
rect 5825 30685 5859 30719
rect 5859 30685 5868 30719
rect 5816 30676 5868 30685
rect 6460 30719 6512 30728
rect 6460 30685 6469 30719
rect 6469 30685 6503 30719
rect 6503 30685 6512 30719
rect 6460 30676 6512 30685
rect 6644 30676 6696 30728
rect 9036 30676 9088 30728
rect 2136 30608 2188 30660
rect 5540 30608 5592 30660
rect 11704 30753 11713 30787
rect 11713 30753 11747 30787
rect 11747 30753 11756 30787
rect 11704 30744 11756 30753
rect 21364 30744 21416 30796
rect 10416 30676 10468 30728
rect 10968 30719 11020 30728
rect 10968 30685 10977 30719
rect 10977 30685 11011 30719
rect 11011 30685 11020 30719
rect 10968 30676 11020 30685
rect 12900 30676 12952 30728
rect 15016 30719 15068 30728
rect 15016 30685 15025 30719
rect 15025 30685 15059 30719
rect 15059 30685 15068 30719
rect 15016 30676 15068 30685
rect 12532 30608 12584 30660
rect 12808 30608 12860 30660
rect 15384 30608 15436 30660
rect 2044 30583 2096 30592
rect 2044 30549 2053 30583
rect 2053 30549 2087 30583
rect 2087 30549 2096 30583
rect 2044 30540 2096 30549
rect 2964 30540 3016 30592
rect 4436 30583 4488 30592
rect 4436 30549 4445 30583
rect 4445 30549 4479 30583
rect 4479 30549 4488 30583
rect 4436 30540 4488 30549
rect 5172 30583 5224 30592
rect 5172 30549 5181 30583
rect 5181 30549 5215 30583
rect 5215 30549 5224 30583
rect 5172 30540 5224 30549
rect 6920 30540 6972 30592
rect 7104 30583 7156 30592
rect 7104 30549 7113 30583
rect 7113 30549 7147 30583
rect 7147 30549 7156 30583
rect 7104 30540 7156 30549
rect 8392 30583 8444 30592
rect 8392 30549 8401 30583
rect 8401 30549 8435 30583
rect 8435 30549 8444 30583
rect 8392 30540 8444 30549
rect 9496 30540 9548 30592
rect 11244 30540 11296 30592
rect 18788 30540 18840 30592
rect 19984 30651 20036 30660
rect 19984 30617 19993 30651
rect 19993 30617 20027 30651
rect 20027 30617 20036 30651
rect 19984 30608 20036 30617
rect 22836 30651 22888 30660
rect 22836 30617 22845 30651
rect 22845 30617 22879 30651
rect 22879 30617 22888 30651
rect 38108 30651 38160 30660
rect 22836 30608 22888 30617
rect 38108 30617 38117 30651
rect 38117 30617 38151 30651
rect 38151 30617 38160 30651
rect 38108 30608 38160 30617
rect 25320 30540 25372 30592
rect 38200 30583 38252 30592
rect 38200 30549 38209 30583
rect 38209 30549 38243 30583
rect 38243 30549 38252 30583
rect 38200 30540 38252 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 5172 30268 5224 30320
rect 10692 30336 10744 30388
rect 10784 30336 10836 30388
rect 3976 30243 4028 30252
rect 3976 30209 3985 30243
rect 3985 30209 4019 30243
rect 4019 30209 4028 30243
rect 3976 30200 4028 30209
rect 5540 30200 5592 30252
rect 8392 30268 8444 30320
rect 8944 30311 8996 30320
rect 8944 30277 8953 30311
rect 8953 30277 8987 30311
rect 8987 30277 8996 30311
rect 8944 30268 8996 30277
rect 9220 30268 9272 30320
rect 9956 30268 10008 30320
rect 1768 30107 1820 30116
rect 1768 30073 1777 30107
rect 1777 30073 1811 30107
rect 1811 30073 1820 30107
rect 1768 30064 1820 30073
rect 4620 30132 4672 30184
rect 5724 30175 5776 30184
rect 5724 30141 5733 30175
rect 5733 30141 5767 30175
rect 5767 30141 5776 30175
rect 5724 30132 5776 30141
rect 10140 30200 10192 30252
rect 10600 30200 10652 30252
rect 12624 30336 12676 30388
rect 16120 30379 16172 30388
rect 16120 30345 16129 30379
rect 16129 30345 16163 30379
rect 16163 30345 16172 30379
rect 16120 30336 16172 30345
rect 13360 30311 13412 30320
rect 13360 30277 13369 30311
rect 13369 30277 13403 30311
rect 13403 30277 13412 30311
rect 13360 30268 13412 30277
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12256 30200 12308 30252
rect 8852 30132 8904 30184
rect 9220 30175 9272 30184
rect 9220 30141 9229 30175
rect 9229 30141 9263 30175
rect 9263 30141 9272 30175
rect 9220 30132 9272 30141
rect 9312 30132 9364 30184
rect 14372 30175 14424 30184
rect 14372 30141 14381 30175
rect 14381 30141 14415 30175
rect 14415 30141 14424 30175
rect 18512 30268 18564 30320
rect 20168 30268 20220 30320
rect 21364 30311 21416 30320
rect 21364 30277 21373 30311
rect 21373 30277 21407 30311
rect 21407 30277 21416 30311
rect 21364 30268 21416 30277
rect 22560 30311 22612 30320
rect 22560 30277 22569 30311
rect 22569 30277 22603 30311
rect 22603 30277 22612 30311
rect 22560 30268 22612 30277
rect 16304 30243 16356 30252
rect 16304 30209 16313 30243
rect 16313 30209 16347 30243
rect 16347 30209 16356 30243
rect 16304 30200 16356 30209
rect 21272 30243 21324 30252
rect 21272 30209 21281 30243
rect 21281 30209 21315 30243
rect 21315 30209 21324 30243
rect 21272 30200 21324 30209
rect 27436 30200 27488 30252
rect 14372 30132 14424 30141
rect 16488 30132 16540 30184
rect 1676 29996 1728 30048
rect 3332 29996 3384 30048
rect 4160 29996 4212 30048
rect 8760 30064 8812 30116
rect 7012 30039 7064 30048
rect 7012 30005 7021 30039
rect 7021 30005 7055 30039
rect 7055 30005 7064 30039
rect 7012 29996 7064 30005
rect 7748 30039 7800 30048
rect 7748 30005 7757 30039
rect 7757 30005 7791 30039
rect 7791 30005 7800 30039
rect 7748 29996 7800 30005
rect 8116 29996 8168 30048
rect 11704 30039 11756 30048
rect 11704 30005 11713 30039
rect 11713 30005 11747 30039
rect 11747 30005 11756 30039
rect 11704 29996 11756 30005
rect 12532 29996 12584 30048
rect 12624 29996 12676 30048
rect 14740 29996 14792 30048
rect 14924 30039 14976 30048
rect 14924 30005 14933 30039
rect 14933 30005 14967 30039
rect 14967 30005 14976 30039
rect 14924 29996 14976 30005
rect 15476 29996 15528 30048
rect 22100 30132 22152 30184
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 7564 29792 7616 29844
rect 8208 29792 8260 29844
rect 11704 29724 11756 29776
rect 11796 29724 11848 29776
rect 13912 29724 13964 29776
rect 6184 29656 6236 29708
rect 9772 29656 9824 29708
rect 10508 29699 10560 29708
rect 10508 29665 10517 29699
rect 10517 29665 10551 29699
rect 10551 29665 10560 29699
rect 11060 29699 11112 29708
rect 10508 29656 10560 29665
rect 11060 29665 11069 29699
rect 11069 29665 11103 29699
rect 11103 29665 11112 29699
rect 11060 29656 11112 29665
rect 12440 29699 12492 29708
rect 12440 29665 12449 29699
rect 12449 29665 12483 29699
rect 12483 29665 12492 29699
rect 12900 29699 12952 29708
rect 12440 29656 12492 29665
rect 12900 29665 12909 29699
rect 12909 29665 12943 29699
rect 12943 29665 12952 29699
rect 12900 29656 12952 29665
rect 14372 29792 14424 29844
rect 15384 29792 15436 29844
rect 15568 29792 15620 29844
rect 18696 29792 18748 29844
rect 15292 29724 15344 29776
rect 20720 29724 20772 29776
rect 18328 29656 18380 29708
rect 18880 29656 18932 29708
rect 2596 29631 2648 29640
rect 2596 29597 2605 29631
rect 2605 29597 2639 29631
rect 2639 29597 2648 29631
rect 2596 29588 2648 29597
rect 4068 29588 4120 29640
rect 4804 29588 4856 29640
rect 6092 29588 6144 29640
rect 3608 29520 3660 29572
rect 4988 29520 5040 29572
rect 8668 29588 8720 29640
rect 8760 29588 8812 29640
rect 10140 29588 10192 29640
rect 14556 29631 14608 29640
rect 14556 29597 14565 29631
rect 14565 29597 14599 29631
rect 14599 29597 14608 29631
rect 14556 29588 14608 29597
rect 14740 29588 14792 29640
rect 16488 29588 16540 29640
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 20904 29588 20956 29640
rect 22836 29792 22888 29844
rect 27804 29792 27856 29844
rect 24492 29588 24544 29640
rect 26056 29631 26108 29640
rect 26056 29597 26065 29631
rect 26065 29597 26099 29631
rect 26099 29597 26108 29631
rect 26056 29588 26108 29597
rect 26976 29588 27028 29640
rect 38292 29631 38344 29640
rect 38292 29597 38301 29631
rect 38301 29597 38335 29631
rect 38335 29597 38344 29631
rect 38292 29588 38344 29597
rect 9864 29520 9916 29572
rect 10600 29563 10652 29572
rect 10600 29529 10618 29563
rect 10618 29529 10652 29563
rect 10600 29520 10652 29529
rect 10784 29520 10836 29572
rect 12624 29520 12676 29572
rect 14280 29520 14332 29572
rect 19524 29563 19576 29572
rect 19524 29529 19533 29563
rect 19533 29529 19567 29563
rect 19567 29529 19576 29563
rect 19524 29520 19576 29529
rect 1768 29495 1820 29504
rect 1768 29461 1777 29495
rect 1777 29461 1811 29495
rect 1811 29461 1820 29495
rect 1768 29452 1820 29461
rect 3792 29452 3844 29504
rect 5356 29452 5408 29504
rect 6368 29452 6420 29504
rect 7472 29452 7524 29504
rect 7840 29495 7892 29504
rect 7840 29461 7849 29495
rect 7849 29461 7883 29495
rect 7883 29461 7892 29495
rect 7840 29452 7892 29461
rect 7932 29452 7984 29504
rect 9128 29452 9180 29504
rect 9772 29495 9824 29504
rect 9772 29461 9781 29495
rect 9781 29461 9815 29495
rect 9815 29461 9824 29495
rect 9772 29452 9824 29461
rect 14464 29452 14516 29504
rect 15752 29495 15804 29504
rect 15752 29461 15761 29495
rect 15761 29461 15795 29495
rect 15795 29461 15804 29495
rect 15752 29452 15804 29461
rect 23940 29452 23992 29504
rect 24032 29452 24084 29504
rect 26516 29452 26568 29504
rect 37004 29452 37056 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 572 29248 624 29300
rect 2136 29180 2188 29232
rect 2412 29112 2464 29164
rect 2872 29112 2924 29164
rect 3884 29112 3936 29164
rect 2780 29044 2832 29096
rect 5080 29112 5132 29164
rect 7196 29180 7248 29232
rect 7656 29180 7708 29232
rect 8944 29248 8996 29300
rect 11796 29248 11848 29300
rect 9312 29180 9364 29232
rect 10232 29223 10284 29232
rect 10232 29189 10241 29223
rect 10241 29189 10275 29223
rect 10275 29189 10284 29223
rect 10232 29180 10284 29189
rect 6920 29112 6972 29164
rect 8208 29112 8260 29164
rect 8300 29155 8352 29164
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 9404 29155 9456 29164
rect 8300 29112 8352 29121
rect 9404 29121 9413 29155
rect 9413 29121 9447 29155
rect 9447 29121 9456 29155
rect 9404 29112 9456 29121
rect 4804 29044 4856 29096
rect 6828 29044 6880 29096
rect 10784 29087 10836 29096
rect 10784 29053 10793 29087
rect 10793 29053 10827 29087
rect 10827 29053 10836 29087
rect 10784 29044 10836 29053
rect 1308 28976 1360 29028
rect 3148 28976 3200 29028
rect 3976 28976 4028 29028
rect 6920 28976 6972 29028
rect 7196 29019 7248 29028
rect 7196 28985 7205 29019
rect 7205 28985 7239 29019
rect 7239 28985 7248 29019
rect 7196 28976 7248 28985
rect 7564 28976 7616 29028
rect 14280 29248 14332 29300
rect 19524 29248 19576 29300
rect 14648 29180 14700 29232
rect 15568 29180 15620 29232
rect 18972 29223 19024 29232
rect 18972 29189 18981 29223
rect 18981 29189 19015 29223
rect 19015 29189 19024 29223
rect 18972 29180 19024 29189
rect 19432 29180 19484 29232
rect 20444 29223 20496 29232
rect 20444 29189 20453 29223
rect 20453 29189 20487 29223
rect 20487 29189 20496 29223
rect 20444 29180 20496 29189
rect 20628 29180 20680 29232
rect 23572 29223 23624 29232
rect 23572 29189 23581 29223
rect 23581 29189 23615 29223
rect 23615 29189 23624 29223
rect 23572 29180 23624 29189
rect 23664 29223 23716 29232
rect 23664 29189 23673 29223
rect 23673 29189 23707 29223
rect 23707 29189 23716 29223
rect 23664 29180 23716 29189
rect 23940 29180 23992 29232
rect 25228 29223 25280 29232
rect 25228 29189 25237 29223
rect 25237 29189 25271 29223
rect 25271 29189 25280 29223
rect 25228 29180 25280 29189
rect 12716 29087 12768 29096
rect 12716 29053 12725 29087
rect 12725 29053 12759 29087
rect 12759 29053 12768 29087
rect 12716 29044 12768 29053
rect 14372 29112 14424 29164
rect 15292 29155 15344 29164
rect 15292 29121 15301 29155
rect 15301 29121 15335 29155
rect 15335 29121 15344 29155
rect 15292 29112 15344 29121
rect 15660 29112 15712 29164
rect 15936 29112 15988 29164
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 13636 29087 13688 29096
rect 13636 29053 13645 29087
rect 13645 29053 13679 29087
rect 13679 29053 13688 29087
rect 13636 29044 13688 29053
rect 13912 29044 13964 29096
rect 18880 29087 18932 29096
rect 13084 28976 13136 29028
rect 18880 29053 18889 29087
rect 18889 29053 18923 29087
rect 18923 29053 18932 29087
rect 18880 29044 18932 29053
rect 19340 29087 19392 29096
rect 19340 29053 19349 29087
rect 19349 29053 19383 29087
rect 19383 29053 19392 29087
rect 19340 29044 19392 29053
rect 21088 29087 21140 29096
rect 21088 29053 21097 29087
rect 21097 29053 21131 29087
rect 21131 29053 21140 29087
rect 21088 29044 21140 29053
rect 23940 29087 23992 29096
rect 23940 29053 23949 29087
rect 23949 29053 23983 29087
rect 23983 29053 23992 29087
rect 23940 29044 23992 29053
rect 1584 28908 1636 28960
rect 9772 28908 9824 28960
rect 13820 28908 13872 28960
rect 18328 28976 18380 29028
rect 18604 28908 18656 28960
rect 19984 28976 20036 29028
rect 26056 29044 26108 29096
rect 37188 29044 37240 29096
rect 27436 28976 27488 29028
rect 20812 28908 20864 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 5172 28704 5224 28756
rect 2596 28636 2648 28688
rect 6092 28636 6144 28688
rect 1952 28543 2004 28552
rect 1952 28509 1961 28543
rect 1961 28509 1995 28543
rect 1995 28509 2004 28543
rect 1952 28500 2004 28509
rect 4068 28500 4120 28552
rect 4896 28500 4948 28552
rect 9404 28636 9456 28688
rect 10876 28568 10928 28620
rect 16856 28704 16908 28756
rect 15200 28636 15252 28688
rect 18972 28704 19024 28756
rect 20076 28704 20128 28756
rect 23388 28704 23440 28756
rect 26884 28747 26936 28756
rect 26884 28713 26893 28747
rect 26893 28713 26927 28747
rect 26927 28713 26936 28747
rect 26884 28704 26936 28713
rect 19064 28636 19116 28688
rect 20260 28636 20312 28688
rect 21916 28636 21968 28688
rect 32404 28636 32456 28688
rect 24308 28568 24360 28620
rect 25320 28611 25372 28620
rect 25320 28577 25329 28611
rect 25329 28577 25363 28611
rect 25363 28577 25372 28611
rect 25320 28568 25372 28577
rect 25504 28568 25556 28620
rect 7564 28500 7616 28552
rect 6552 28432 6604 28484
rect 7012 28475 7064 28484
rect 7012 28441 7021 28475
rect 7021 28441 7055 28475
rect 7055 28441 7064 28475
rect 7012 28432 7064 28441
rect 8300 28432 8352 28484
rect 9404 28500 9456 28552
rect 9864 28500 9916 28552
rect 10324 28500 10376 28552
rect 2228 28364 2280 28416
rect 2688 28407 2740 28416
rect 2688 28373 2697 28407
rect 2697 28373 2731 28407
rect 2731 28373 2740 28407
rect 2688 28364 2740 28373
rect 3884 28364 3936 28416
rect 4068 28407 4120 28416
rect 4068 28373 4077 28407
rect 4077 28373 4111 28407
rect 4111 28373 4120 28407
rect 4068 28364 4120 28373
rect 4620 28364 4672 28416
rect 5264 28364 5316 28416
rect 6092 28364 6144 28416
rect 8760 28364 8812 28416
rect 9588 28432 9640 28484
rect 11520 28500 11572 28552
rect 16212 28543 16264 28552
rect 16212 28509 16221 28543
rect 16221 28509 16255 28543
rect 16255 28509 16264 28543
rect 16212 28500 16264 28509
rect 16580 28500 16632 28552
rect 16764 28500 16816 28552
rect 17408 28500 17460 28552
rect 17592 28500 17644 28552
rect 12348 28475 12400 28484
rect 12348 28441 12357 28475
rect 12357 28441 12391 28475
rect 12391 28441 12400 28475
rect 12348 28432 12400 28441
rect 13360 28475 13412 28484
rect 9772 28364 9824 28416
rect 10048 28407 10100 28416
rect 10048 28373 10057 28407
rect 10057 28373 10091 28407
rect 10091 28373 10100 28407
rect 10048 28364 10100 28373
rect 10416 28364 10468 28416
rect 13360 28441 13369 28475
rect 13369 28441 13403 28475
rect 13403 28441 13412 28475
rect 13360 28432 13412 28441
rect 13728 28432 13780 28484
rect 14924 28432 14976 28484
rect 15384 28475 15436 28484
rect 15384 28441 15393 28475
rect 15393 28441 15427 28475
rect 15427 28441 15436 28475
rect 15384 28432 15436 28441
rect 19064 28500 19116 28552
rect 20352 28543 20404 28552
rect 20352 28509 20361 28543
rect 20361 28509 20395 28543
rect 20395 28509 20404 28543
rect 20352 28500 20404 28509
rect 20812 28543 20864 28552
rect 20812 28509 20821 28543
rect 20821 28509 20855 28543
rect 20855 28509 20864 28543
rect 20812 28500 20864 28509
rect 21916 28543 21968 28552
rect 21916 28509 21925 28543
rect 21925 28509 21959 28543
rect 21959 28509 21968 28543
rect 21916 28500 21968 28509
rect 23848 28500 23900 28552
rect 27436 28543 27488 28552
rect 27436 28509 27445 28543
rect 27445 28509 27479 28543
rect 27479 28509 27488 28543
rect 27436 28500 27488 28509
rect 37004 28500 37056 28552
rect 12532 28364 12584 28416
rect 19156 28432 19208 28484
rect 24952 28432 25004 28484
rect 25412 28475 25464 28484
rect 25412 28441 25421 28475
rect 25421 28441 25455 28475
rect 25455 28441 25464 28475
rect 25412 28432 25464 28441
rect 26148 28432 26200 28484
rect 15752 28364 15804 28416
rect 19064 28364 19116 28416
rect 19340 28364 19392 28416
rect 20260 28364 20312 28416
rect 21548 28364 21600 28416
rect 25964 28364 26016 28416
rect 32036 28407 32088 28416
rect 32036 28373 32045 28407
rect 32045 28373 32079 28407
rect 32079 28373 32088 28407
rect 32036 28364 32088 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 3884 28092 3936 28144
rect 5816 28092 5868 28144
rect 6460 28092 6512 28144
rect 1584 28067 1636 28076
rect 1584 28033 1593 28067
rect 1593 28033 1627 28067
rect 1627 28033 1636 28067
rect 1584 28024 1636 28033
rect 2872 28024 2924 28076
rect 3424 28024 3476 28076
rect 4804 28024 4856 28076
rect 1768 27931 1820 27940
rect 1768 27897 1777 27931
rect 1777 27897 1811 27931
rect 1811 27897 1820 27931
rect 1768 27888 1820 27897
rect 3884 27888 3936 27940
rect 5724 27956 5776 28008
rect 6920 28160 6972 28212
rect 7380 28092 7432 28144
rect 9036 28160 9088 28212
rect 10968 28160 11020 28212
rect 17132 28160 17184 28212
rect 19248 28160 19300 28212
rect 23756 28160 23808 28212
rect 25412 28160 25464 28212
rect 8484 28067 8536 28076
rect 8484 28033 8493 28067
rect 8493 28033 8527 28067
rect 8527 28033 8536 28067
rect 8484 28024 8536 28033
rect 5540 27888 5592 27940
rect 5908 27820 5960 27872
rect 7104 27956 7156 28008
rect 9680 28092 9732 28144
rect 9772 28092 9824 28144
rect 11152 28092 11204 28144
rect 13820 28092 13872 28144
rect 18604 28135 18656 28144
rect 18604 28101 18613 28135
rect 18613 28101 18647 28135
rect 18647 28101 18656 28135
rect 18604 28092 18656 28101
rect 18972 28092 19024 28144
rect 20076 28092 20128 28144
rect 20260 28092 20312 28144
rect 22100 28135 22152 28144
rect 22100 28101 22109 28135
rect 22109 28101 22143 28135
rect 22143 28101 22152 28135
rect 22100 28092 22152 28101
rect 25964 28160 26016 28212
rect 8944 28024 8996 28076
rect 9956 28067 10008 28076
rect 9956 28033 9965 28067
rect 9965 28033 9999 28067
rect 9999 28033 10008 28067
rect 9956 28024 10008 28033
rect 10140 28024 10192 28076
rect 12440 28024 12492 28076
rect 11428 27956 11480 28008
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 14188 28024 14240 28076
rect 15568 28024 15620 28076
rect 16396 28024 16448 28076
rect 17040 28024 17092 28076
rect 17500 28067 17552 28076
rect 17500 28033 17509 28067
rect 17509 28033 17543 28067
rect 17543 28033 17552 28067
rect 17500 28024 17552 28033
rect 13636 27956 13688 28008
rect 7748 27888 7800 27940
rect 8484 27888 8536 27940
rect 7104 27820 7156 27872
rect 8392 27820 8444 27872
rect 8668 27820 8720 27872
rect 14004 27888 14056 27940
rect 10692 27863 10744 27872
rect 10692 27829 10701 27863
rect 10701 27829 10735 27863
rect 10735 27829 10744 27863
rect 10692 27820 10744 27829
rect 10968 27820 11020 27872
rect 13084 27820 13136 27872
rect 13176 27820 13228 27872
rect 16672 27956 16724 28008
rect 17408 27956 17460 28008
rect 16120 27888 16172 27940
rect 19432 27956 19484 28008
rect 20536 27956 20588 28008
rect 22468 27956 22520 28008
rect 24216 28067 24268 28076
rect 24216 28033 24225 28067
rect 24225 28033 24259 28067
rect 24259 28033 24268 28067
rect 24216 28024 24268 28033
rect 25136 28024 25188 28076
rect 27804 28024 27856 28076
rect 24768 27956 24820 28008
rect 24952 27956 25004 28008
rect 27436 27956 27488 28008
rect 30748 27888 30800 27940
rect 16304 27820 16356 27872
rect 16948 27863 17000 27872
rect 16948 27829 16957 27863
rect 16957 27829 16991 27863
rect 16991 27829 17000 27863
rect 16948 27820 17000 27829
rect 17500 27820 17552 27872
rect 37648 27820 37700 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4804 27616 4856 27668
rect 9772 27616 9824 27668
rect 9864 27616 9916 27668
rect 10048 27548 10100 27600
rect 10324 27548 10376 27600
rect 10968 27548 11020 27600
rect 3240 27455 3292 27464
rect 3240 27421 3249 27455
rect 3249 27421 3283 27455
rect 3283 27421 3292 27455
rect 3240 27412 3292 27421
rect 6000 27480 6052 27532
rect 6828 27480 6880 27532
rect 8208 27480 8260 27532
rect 9404 27480 9456 27532
rect 9588 27523 9640 27532
rect 9588 27489 9597 27523
rect 9597 27489 9631 27523
rect 9631 27489 9640 27523
rect 9588 27480 9640 27489
rect 11060 27480 11112 27532
rect 12716 27480 12768 27532
rect 4804 27412 4856 27464
rect 4988 27412 5040 27464
rect 2872 27344 2924 27396
rect 5632 27387 5684 27396
rect 5632 27353 5641 27387
rect 5641 27353 5675 27387
rect 5675 27353 5684 27387
rect 5632 27344 5684 27353
rect 1768 27319 1820 27328
rect 1768 27285 1777 27319
rect 1777 27285 1811 27319
rect 1811 27285 1820 27319
rect 1768 27276 1820 27285
rect 2412 27276 2464 27328
rect 3332 27319 3384 27328
rect 3332 27285 3341 27319
rect 3341 27285 3375 27319
rect 3375 27285 3384 27319
rect 3332 27276 3384 27285
rect 4804 27276 4856 27328
rect 5172 27276 5224 27328
rect 5448 27276 5500 27328
rect 5816 27344 5868 27396
rect 6920 27412 6972 27464
rect 8760 27412 8812 27464
rect 11888 27412 11940 27464
rect 15108 27616 15160 27668
rect 13084 27548 13136 27600
rect 16212 27548 16264 27600
rect 16396 27616 16448 27668
rect 25136 27616 25188 27668
rect 16580 27548 16632 27600
rect 20720 27591 20772 27600
rect 20720 27557 20729 27591
rect 20729 27557 20763 27591
rect 20763 27557 20772 27591
rect 20720 27548 20772 27557
rect 21456 27548 21508 27600
rect 21916 27548 21968 27600
rect 14004 27480 14056 27532
rect 7012 27344 7064 27396
rect 9220 27387 9272 27396
rect 8392 27276 8444 27328
rect 9220 27353 9229 27387
rect 9229 27353 9263 27387
rect 9263 27353 9272 27387
rect 9220 27344 9272 27353
rect 9680 27344 9732 27396
rect 10968 27344 11020 27396
rect 12532 27344 12584 27396
rect 12992 27344 13044 27396
rect 11060 27276 11112 27328
rect 14280 27344 14332 27396
rect 14648 27344 14700 27396
rect 14096 27276 14148 27328
rect 15200 27344 15252 27396
rect 15292 27344 15344 27396
rect 16120 27387 16172 27396
rect 16120 27353 16129 27387
rect 16129 27353 16163 27387
rect 16163 27353 16172 27387
rect 16120 27344 16172 27353
rect 16212 27387 16264 27396
rect 16212 27353 16221 27387
rect 16221 27353 16255 27387
rect 16255 27353 16264 27387
rect 20812 27480 20864 27532
rect 21548 27480 21600 27532
rect 24768 27548 24820 27600
rect 24860 27480 24912 27532
rect 25504 27480 25556 27532
rect 26516 27480 26568 27532
rect 17040 27412 17092 27464
rect 17868 27412 17920 27464
rect 18512 27412 18564 27464
rect 19156 27412 19208 27464
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 16212 27344 16264 27353
rect 17408 27344 17460 27396
rect 18052 27344 18104 27396
rect 17684 27319 17736 27328
rect 17684 27285 17693 27319
rect 17693 27285 17727 27319
rect 17727 27285 17736 27319
rect 17684 27276 17736 27285
rect 19984 27276 20036 27328
rect 21456 27387 21508 27396
rect 21456 27353 21465 27387
rect 21465 27353 21499 27387
rect 21499 27353 21508 27387
rect 21456 27344 21508 27353
rect 21364 27276 21416 27328
rect 22376 27344 22428 27396
rect 25872 27344 25924 27396
rect 26056 27276 26108 27328
rect 37372 27480 37424 27532
rect 27896 27412 27948 27464
rect 37464 27455 37516 27464
rect 37464 27421 37473 27455
rect 37473 27421 37507 27455
rect 37507 27421 37516 27455
rect 37464 27412 37516 27421
rect 27252 27387 27304 27396
rect 27252 27353 27261 27387
rect 27261 27353 27295 27387
rect 27295 27353 27304 27387
rect 27252 27344 27304 27353
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4896 27072 4948 27124
rect 940 27004 992 27056
rect 2136 26936 2188 26988
rect 2596 26979 2648 26988
rect 2596 26945 2605 26979
rect 2605 26945 2639 26979
rect 2639 26945 2648 26979
rect 2596 26936 2648 26945
rect 3240 26979 3292 26988
rect 3240 26945 3249 26979
rect 3249 26945 3283 26979
rect 3283 26945 3292 26979
rect 3240 26936 3292 26945
rect 1584 26868 1636 26920
rect 4068 26936 4120 26988
rect 5724 26936 5776 26988
rect 5448 26868 5500 26920
rect 6736 26936 6788 26988
rect 7196 27004 7248 27056
rect 9220 27072 9272 27124
rect 11244 27072 11296 27124
rect 12716 27072 12768 27124
rect 14280 27072 14332 27124
rect 14648 27072 14700 27124
rect 21272 27072 21324 27124
rect 21456 27072 21508 27124
rect 25872 27115 25924 27124
rect 25872 27081 25881 27115
rect 25881 27081 25915 27115
rect 25915 27081 25924 27115
rect 25872 27072 25924 27081
rect 27252 27072 27304 27124
rect 30748 27115 30800 27124
rect 7380 26936 7432 26988
rect 8208 26911 8260 26920
rect 6644 26856 6696 26908
rect 8208 26877 8217 26911
rect 8217 26877 8251 26911
rect 8251 26877 8260 26911
rect 8208 26868 8260 26877
rect 4988 26800 5040 26852
rect 6184 26800 6236 26852
rect 9496 27047 9548 27056
rect 9496 27013 9505 27047
rect 9505 27013 9539 27047
rect 9539 27013 9548 27047
rect 9496 27004 9548 27013
rect 10876 27004 10928 27056
rect 12440 27004 12492 27056
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 13176 27004 13228 27056
rect 13360 26936 13412 26988
rect 13544 26979 13596 26988
rect 13544 26945 13553 26979
rect 13553 26945 13587 26979
rect 13587 26945 13596 26979
rect 13544 26936 13596 26945
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 18512 27004 18564 27056
rect 19064 27047 19116 27056
rect 19064 27013 19073 27047
rect 19073 27013 19107 27047
rect 19107 27013 19116 27047
rect 19064 27004 19116 27013
rect 19340 27004 19392 27056
rect 19432 27004 19484 27056
rect 22468 27004 22520 27056
rect 22744 27047 22796 27056
rect 22744 27013 22753 27047
rect 22753 27013 22787 27047
rect 22787 27013 22796 27047
rect 22744 27004 22796 27013
rect 23296 27004 23348 27056
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 16028 26936 16080 26988
rect 17316 26936 17368 26988
rect 17592 26936 17644 26988
rect 18696 26936 18748 26988
rect 12440 26868 12492 26920
rect 12900 26868 12952 26920
rect 13268 26868 13320 26920
rect 20168 26936 20220 26988
rect 20352 26936 20404 26988
rect 20720 26868 20772 26920
rect 2044 26775 2096 26784
rect 2044 26741 2053 26775
rect 2053 26741 2087 26775
rect 2087 26741 2096 26775
rect 2044 26732 2096 26741
rect 2596 26732 2648 26784
rect 5080 26732 5132 26784
rect 6644 26732 6696 26784
rect 7012 26732 7064 26784
rect 7196 26732 7248 26784
rect 7380 26775 7432 26784
rect 7380 26741 7389 26775
rect 7389 26741 7423 26775
rect 7423 26741 7432 26775
rect 7380 26732 7432 26741
rect 9864 26800 9916 26852
rect 12256 26800 12308 26852
rect 15568 26800 15620 26852
rect 10692 26732 10744 26784
rect 11060 26775 11112 26784
rect 11060 26741 11069 26775
rect 11069 26741 11103 26775
rect 11103 26741 11112 26775
rect 11060 26732 11112 26741
rect 13452 26732 13504 26784
rect 14924 26775 14976 26784
rect 14924 26741 14933 26775
rect 14933 26741 14967 26775
rect 14967 26741 14976 26775
rect 14924 26732 14976 26741
rect 15200 26732 15252 26784
rect 16948 26775 17000 26784
rect 16948 26741 16957 26775
rect 16957 26741 16991 26775
rect 16991 26741 17000 26775
rect 16948 26732 17000 26741
rect 17592 26775 17644 26784
rect 17592 26741 17601 26775
rect 17601 26741 17635 26775
rect 17635 26741 17644 26775
rect 17592 26732 17644 26741
rect 18236 26775 18288 26784
rect 18236 26741 18245 26775
rect 18245 26741 18279 26775
rect 18279 26741 18288 26775
rect 18236 26732 18288 26741
rect 20444 26732 20496 26784
rect 22008 26936 22060 26988
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 21916 26868 21968 26920
rect 21824 26800 21876 26852
rect 27712 26868 27764 26920
rect 30748 27081 30757 27115
rect 30757 27081 30791 27115
rect 30791 27081 30800 27115
rect 30748 27072 30800 27081
rect 30840 27072 30892 27124
rect 28816 27004 28868 27056
rect 38200 27004 38252 27056
rect 38292 26979 38344 26988
rect 32036 26868 32088 26920
rect 25872 26732 25924 26784
rect 28908 26800 28960 26852
rect 38292 26945 38301 26979
rect 38301 26945 38335 26979
rect 38335 26945 38344 26979
rect 38292 26936 38344 26945
rect 29000 26732 29052 26784
rect 29828 26732 29880 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3332 26528 3384 26580
rect 9312 26528 9364 26580
rect 10048 26528 10100 26580
rect 2964 26392 3016 26444
rect 4344 26460 4396 26512
rect 4896 26460 4948 26512
rect 5080 26460 5132 26512
rect 4160 26392 4212 26444
rect 4712 26392 4764 26444
rect 10140 26392 10192 26444
rect 10784 26392 10836 26444
rect 4896 26324 4948 26376
rect 5816 26367 5868 26376
rect 5816 26333 5825 26367
rect 5825 26333 5859 26367
rect 5859 26333 5868 26367
rect 5816 26324 5868 26333
rect 6184 26324 6236 26376
rect 1768 26231 1820 26240
rect 1768 26197 1777 26231
rect 1777 26197 1811 26231
rect 1811 26197 1820 26231
rect 1768 26188 1820 26197
rect 2780 26299 2832 26308
rect 2780 26265 2789 26299
rect 2789 26265 2823 26299
rect 2823 26265 2832 26299
rect 2780 26256 2832 26265
rect 2964 26188 3016 26240
rect 4160 26299 4212 26308
rect 4160 26265 4169 26299
rect 4169 26265 4203 26299
rect 4203 26265 4212 26299
rect 4160 26256 4212 26265
rect 5724 26256 5776 26308
rect 7012 26256 7064 26308
rect 6552 26188 6604 26240
rect 7932 26256 7984 26308
rect 8024 26256 8076 26308
rect 9036 26324 9088 26376
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 12440 26460 12492 26512
rect 11980 26435 12032 26444
rect 11980 26401 11989 26435
rect 11989 26401 12023 26435
rect 12023 26401 12032 26435
rect 11980 26392 12032 26401
rect 13268 26392 13320 26444
rect 14004 26460 14056 26512
rect 14648 26435 14700 26444
rect 14648 26401 14657 26435
rect 14657 26401 14691 26435
rect 14691 26401 14700 26435
rect 14648 26392 14700 26401
rect 9864 26324 9916 26333
rect 12716 26324 12768 26376
rect 9312 26299 9364 26308
rect 9312 26265 9321 26299
rect 9321 26265 9355 26299
rect 9355 26265 9364 26299
rect 9312 26256 9364 26265
rect 10692 26256 10744 26308
rect 11796 26256 11848 26308
rect 12440 26256 12492 26308
rect 12532 26256 12584 26308
rect 13268 26256 13320 26308
rect 13820 26256 13872 26308
rect 14372 26299 14424 26308
rect 14372 26265 14381 26299
rect 14381 26265 14415 26299
rect 14415 26265 14424 26299
rect 14372 26256 14424 26265
rect 14464 26299 14516 26308
rect 14464 26265 14473 26299
rect 14473 26265 14507 26299
rect 14507 26265 14516 26299
rect 15844 26460 15896 26512
rect 15660 26435 15712 26444
rect 15660 26401 15669 26435
rect 15669 26401 15703 26435
rect 15703 26401 15712 26435
rect 15660 26392 15712 26401
rect 16120 26392 16172 26444
rect 16580 26392 16632 26444
rect 17776 26392 17828 26444
rect 18144 26392 18196 26444
rect 18788 26392 18840 26444
rect 22192 26528 22244 26580
rect 22376 26571 22428 26580
rect 22376 26537 22385 26571
rect 22385 26537 22419 26571
rect 22419 26537 22428 26571
rect 22376 26528 22428 26537
rect 26424 26528 26476 26580
rect 20812 26460 20864 26512
rect 22100 26392 22152 26444
rect 22192 26392 22244 26444
rect 23204 26392 23256 26444
rect 17316 26324 17368 26376
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 22284 26367 22336 26376
rect 22284 26333 22293 26367
rect 22293 26333 22327 26367
rect 22327 26333 22336 26367
rect 22284 26324 22336 26333
rect 22928 26367 22980 26376
rect 22928 26333 22937 26367
rect 22937 26333 22971 26367
rect 22971 26333 22980 26367
rect 22928 26324 22980 26333
rect 25780 26392 25832 26444
rect 27620 26528 27672 26580
rect 28816 26571 28868 26580
rect 28816 26537 28825 26571
rect 28825 26537 28859 26571
rect 28859 26537 28868 26571
rect 28816 26528 28868 26537
rect 37740 26528 37792 26580
rect 38200 26503 38252 26512
rect 27712 26435 27764 26444
rect 27712 26401 27721 26435
rect 27721 26401 27755 26435
rect 27755 26401 27764 26435
rect 27712 26392 27764 26401
rect 38200 26469 38209 26503
rect 38209 26469 38243 26503
rect 38243 26469 38252 26503
rect 38200 26460 38252 26469
rect 28724 26367 28776 26376
rect 28724 26333 28733 26367
rect 28733 26333 28767 26367
rect 28767 26333 28776 26367
rect 28724 26324 28776 26333
rect 36544 26367 36596 26376
rect 36544 26333 36553 26367
rect 36553 26333 36587 26367
rect 36587 26333 36596 26367
rect 36544 26324 36596 26333
rect 14464 26256 14516 26265
rect 16580 26256 16632 26308
rect 19248 26256 19300 26308
rect 19984 26256 20036 26308
rect 9036 26188 9088 26240
rect 9496 26188 9548 26240
rect 13912 26188 13964 26240
rect 14004 26188 14056 26240
rect 17224 26231 17276 26240
rect 17224 26197 17233 26231
rect 17233 26197 17267 26231
rect 17267 26197 17276 26231
rect 17224 26188 17276 26197
rect 21364 26256 21416 26308
rect 30840 26256 30892 26308
rect 23388 26188 23440 26240
rect 25596 26188 25648 26240
rect 27252 26188 27304 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2228 25984 2280 26036
rect 2780 25984 2832 26036
rect 2320 25959 2372 25968
rect 2320 25925 2329 25959
rect 2329 25925 2363 25959
rect 2363 25925 2372 25959
rect 2320 25916 2372 25925
rect 3424 25916 3476 25968
rect 4068 25916 4120 25968
rect 5264 25984 5316 26036
rect 4252 25916 4304 25968
rect 2228 25823 2280 25832
rect 2228 25789 2237 25823
rect 2237 25789 2271 25823
rect 2271 25789 2280 25823
rect 2228 25780 2280 25789
rect 3332 25780 3384 25832
rect 4344 25823 4396 25832
rect 4344 25789 4353 25823
rect 4353 25789 4387 25823
rect 4387 25789 4396 25823
rect 4344 25780 4396 25789
rect 4804 25916 4856 25968
rect 8024 25959 8076 25968
rect 8024 25925 8033 25959
rect 8033 25925 8067 25959
rect 8067 25925 8076 25959
rect 8024 25916 8076 25925
rect 8300 25916 8352 25968
rect 8576 25916 8628 25968
rect 8852 25916 8904 25968
rect 10140 25959 10192 25968
rect 10140 25925 10149 25959
rect 10149 25925 10183 25959
rect 10183 25925 10192 25959
rect 10140 25916 10192 25925
rect 11336 25916 11388 25968
rect 12440 25984 12492 26036
rect 15844 25984 15896 26036
rect 16488 25984 16540 26036
rect 18328 25984 18380 26036
rect 22744 26027 22796 26036
rect 7288 25891 7340 25900
rect 5908 25823 5960 25832
rect 5908 25789 5917 25823
rect 5917 25789 5951 25823
rect 5951 25789 5960 25823
rect 5908 25780 5960 25789
rect 7288 25857 7297 25891
rect 7297 25857 7331 25891
rect 7331 25857 7340 25891
rect 7288 25848 7340 25857
rect 14004 25916 14056 25968
rect 15384 25916 15436 25968
rect 16028 25916 16080 25968
rect 20260 25916 20312 25968
rect 13912 25891 13964 25900
rect 13912 25857 13921 25891
rect 13921 25857 13955 25891
rect 13955 25857 13964 25891
rect 13912 25848 13964 25857
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 14832 25848 14884 25900
rect 15200 25891 15252 25900
rect 15200 25857 15209 25891
rect 15209 25857 15243 25891
rect 15243 25857 15252 25891
rect 15200 25848 15252 25857
rect 17684 25891 17736 25900
rect 17684 25857 17693 25891
rect 17693 25857 17727 25891
rect 17727 25857 17736 25891
rect 17684 25848 17736 25857
rect 18328 25891 18380 25900
rect 18328 25857 18337 25891
rect 18337 25857 18371 25891
rect 18371 25857 18380 25891
rect 18328 25848 18380 25857
rect 6920 25780 6972 25832
rect 8392 25823 8444 25832
rect 8392 25789 8401 25823
rect 8401 25789 8435 25823
rect 8435 25789 8444 25823
rect 8392 25780 8444 25789
rect 9128 25780 9180 25832
rect 9588 25780 9640 25832
rect 10324 25823 10376 25832
rect 10324 25789 10333 25823
rect 10333 25789 10367 25823
rect 10367 25789 10376 25823
rect 10324 25780 10376 25789
rect 12808 25823 12860 25832
rect 5356 25712 5408 25764
rect 5632 25712 5684 25764
rect 12808 25789 12817 25823
rect 12817 25789 12851 25823
rect 12851 25789 12860 25823
rect 12808 25780 12860 25789
rect 13728 25780 13780 25832
rect 15568 25780 15620 25832
rect 20812 25848 20864 25900
rect 21180 25848 21232 25900
rect 21824 25848 21876 25900
rect 22744 25993 22753 26027
rect 22753 25993 22787 26027
rect 22787 25993 22796 26027
rect 22744 25984 22796 25993
rect 23388 26027 23440 26036
rect 23388 25993 23397 26027
rect 23397 25993 23431 26027
rect 23431 25993 23440 26027
rect 23388 25984 23440 25993
rect 24124 25984 24176 26036
rect 28724 25984 28776 26036
rect 33876 25984 33928 26036
rect 25596 25959 25648 25968
rect 25596 25925 25605 25959
rect 25605 25925 25639 25959
rect 25639 25925 25648 25959
rect 25596 25916 25648 25925
rect 27344 25959 27396 25968
rect 27344 25925 27353 25959
rect 27353 25925 27387 25959
rect 27387 25925 27396 25959
rect 27344 25916 27396 25925
rect 28908 25916 28960 25968
rect 13636 25712 13688 25764
rect 13912 25712 13964 25764
rect 2964 25644 3016 25696
rect 5264 25644 5316 25696
rect 10140 25644 10192 25696
rect 13360 25687 13412 25696
rect 13360 25653 13369 25687
rect 13369 25653 13403 25687
rect 13403 25653 13412 25687
rect 13360 25644 13412 25653
rect 15384 25644 15436 25696
rect 15936 25687 15988 25696
rect 15936 25653 15945 25687
rect 15945 25653 15979 25687
rect 15979 25653 15988 25687
rect 15936 25644 15988 25653
rect 18880 25644 18932 25696
rect 19340 25712 19392 25764
rect 19524 25712 19576 25764
rect 21640 25780 21692 25832
rect 23112 25848 23164 25900
rect 24216 25848 24268 25900
rect 30840 25848 30892 25900
rect 23756 25780 23808 25832
rect 27252 25823 27304 25832
rect 21088 25712 21140 25764
rect 22652 25712 22704 25764
rect 26240 25712 26292 25764
rect 19432 25644 19484 25696
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 22192 25644 22244 25696
rect 24400 25644 24452 25696
rect 27252 25789 27261 25823
rect 27261 25789 27295 25823
rect 27295 25789 27304 25823
rect 27252 25780 27304 25789
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 1492 25440 1544 25492
rect 3332 25440 3384 25492
rect 5724 25440 5776 25492
rect 6276 25440 6328 25492
rect 6736 25440 6788 25492
rect 7288 25440 7340 25492
rect 9496 25440 9548 25492
rect 15476 25440 15528 25492
rect 16212 25440 16264 25492
rect 16488 25440 16540 25492
rect 19800 25440 19852 25492
rect 22284 25440 22336 25492
rect 27528 25440 27580 25492
rect 27620 25440 27672 25492
rect 29460 25440 29512 25492
rect 29920 25483 29972 25492
rect 29920 25449 29929 25483
rect 29929 25449 29963 25483
rect 29963 25449 29972 25483
rect 29920 25440 29972 25449
rect 6000 25372 6052 25424
rect 8116 25372 8168 25424
rect 9312 25372 9364 25424
rect 5264 25304 5316 25356
rect 1952 25279 2004 25288
rect 1952 25245 1961 25279
rect 1961 25245 1995 25279
rect 1995 25245 2004 25279
rect 1952 25236 2004 25245
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 4712 25236 4764 25288
rect 9128 25304 9180 25356
rect 10232 25304 10284 25356
rect 6276 25236 6328 25288
rect 3240 25211 3292 25220
rect 3240 25177 3249 25211
rect 3249 25177 3283 25211
rect 3283 25177 3292 25211
rect 3240 25168 3292 25177
rect 4988 25211 5040 25220
rect 4988 25177 4997 25211
rect 4997 25177 5031 25211
rect 5031 25177 5040 25211
rect 9496 25236 9548 25288
rect 14004 25304 14056 25356
rect 15200 25372 15252 25424
rect 11336 25279 11388 25288
rect 4988 25168 5040 25177
rect 4528 25100 4580 25152
rect 6828 25100 6880 25152
rect 8668 25168 8720 25220
rect 8116 25143 8168 25152
rect 8116 25109 8125 25143
rect 8125 25109 8159 25143
rect 8159 25109 8168 25143
rect 8116 25100 8168 25109
rect 8208 25100 8260 25152
rect 9496 25100 9548 25152
rect 11336 25245 11345 25279
rect 11345 25245 11379 25279
rect 11379 25245 11388 25279
rect 11336 25236 11388 25245
rect 13544 25279 13596 25288
rect 13544 25245 13553 25279
rect 13553 25245 13587 25279
rect 13587 25245 13596 25279
rect 13544 25236 13596 25245
rect 14832 25279 14884 25288
rect 14832 25245 14833 25279
rect 14833 25245 14867 25279
rect 14867 25245 14884 25279
rect 14832 25236 14884 25245
rect 15844 25236 15896 25288
rect 17960 25236 18012 25288
rect 18696 25279 18748 25288
rect 18696 25245 18705 25279
rect 18705 25245 18739 25279
rect 18739 25245 18748 25279
rect 18696 25236 18748 25245
rect 18972 25304 19024 25356
rect 19800 25347 19852 25356
rect 19800 25313 19809 25347
rect 19809 25313 19843 25347
rect 19843 25313 19852 25347
rect 19800 25304 19852 25313
rect 28632 25372 28684 25424
rect 22192 25304 22244 25356
rect 22376 25347 22428 25356
rect 22376 25313 22385 25347
rect 22385 25313 22419 25347
rect 22419 25313 22428 25347
rect 22376 25304 22428 25313
rect 26240 25347 26292 25356
rect 26240 25313 26249 25347
rect 26249 25313 26283 25347
rect 26283 25313 26292 25347
rect 26240 25304 26292 25313
rect 27252 25304 27304 25356
rect 36544 25304 36596 25356
rect 10876 25168 10928 25220
rect 11612 25211 11664 25220
rect 11612 25177 11621 25211
rect 11621 25177 11655 25211
rect 11655 25177 11664 25211
rect 11612 25168 11664 25177
rect 15936 25168 15988 25220
rect 12440 25100 12492 25152
rect 12532 25100 12584 25152
rect 13636 25143 13688 25152
rect 13636 25109 13645 25143
rect 13645 25109 13679 25143
rect 13679 25109 13688 25143
rect 13636 25100 13688 25109
rect 13820 25100 13872 25152
rect 16304 25211 16356 25220
rect 16304 25177 16313 25211
rect 16313 25177 16347 25211
rect 16347 25177 16356 25211
rect 16304 25168 16356 25177
rect 17500 25168 17552 25220
rect 16580 25100 16632 25152
rect 19524 25168 19576 25220
rect 18236 25100 18288 25152
rect 18788 25143 18840 25152
rect 18788 25109 18797 25143
rect 18797 25109 18831 25143
rect 18831 25109 18840 25143
rect 18788 25100 18840 25109
rect 19340 25100 19392 25152
rect 22284 25168 22336 25220
rect 22468 25168 22520 25220
rect 29092 25236 29144 25288
rect 26700 25168 26752 25220
rect 37648 25211 37700 25220
rect 25044 25100 25096 25152
rect 26056 25100 26108 25152
rect 37648 25177 37657 25211
rect 37657 25177 37691 25211
rect 37691 25177 37700 25211
rect 37648 25168 37700 25177
rect 27068 25100 27120 25152
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 1952 24896 2004 24948
rect 4436 24896 4488 24948
rect 4712 24896 4764 24948
rect 8208 24896 8260 24948
rect 8300 24896 8352 24948
rect 18788 24896 18840 24948
rect 1768 24828 1820 24880
rect 2320 24828 2372 24880
rect 3424 24828 3476 24880
rect 4620 24828 4672 24880
rect 5264 24828 5316 24880
rect 6000 24828 6052 24880
rect 7288 24828 7340 24880
rect 11244 24828 11296 24880
rect 11704 24828 11756 24880
rect 13728 24828 13780 24880
rect 14096 24871 14148 24880
rect 14096 24837 14105 24871
rect 14105 24837 14139 24871
rect 14139 24837 14148 24871
rect 14096 24828 14148 24837
rect 15752 24871 15804 24880
rect 15752 24837 15761 24871
rect 15761 24837 15795 24871
rect 15795 24837 15804 24871
rect 15752 24828 15804 24837
rect 17040 24871 17092 24880
rect 17040 24837 17049 24871
rect 17049 24837 17083 24871
rect 17083 24837 17092 24871
rect 17040 24828 17092 24837
rect 17500 24828 17552 24880
rect 20260 24896 20312 24948
rect 22284 24896 22336 24948
rect 23204 24896 23256 24948
rect 27344 24896 27396 24948
rect 19248 24828 19300 24880
rect 20812 24871 20864 24880
rect 20812 24837 20821 24871
rect 20821 24837 20855 24871
rect 20855 24837 20864 24871
rect 20812 24828 20864 24837
rect 20996 24828 21048 24880
rect 23480 24871 23532 24880
rect 3700 24760 3752 24812
rect 7748 24803 7800 24812
rect 7748 24769 7757 24803
rect 7757 24769 7791 24803
rect 7791 24769 7800 24803
rect 7748 24760 7800 24769
rect 10600 24760 10652 24812
rect 1860 24692 1912 24744
rect 4988 24692 5040 24744
rect 4620 24624 4672 24676
rect 3424 24599 3476 24608
rect 3424 24565 3433 24599
rect 3433 24565 3467 24599
rect 3467 24565 3476 24599
rect 3424 24556 3476 24565
rect 4528 24556 4580 24608
rect 5264 24556 5316 24608
rect 5908 24692 5960 24744
rect 8392 24735 8444 24744
rect 8392 24701 8401 24735
rect 8401 24701 8435 24735
rect 8435 24701 8444 24735
rect 8392 24692 8444 24701
rect 9128 24692 9180 24744
rect 7196 24667 7248 24676
rect 7196 24633 7205 24667
rect 7205 24633 7239 24667
rect 7239 24633 7248 24667
rect 7196 24624 7248 24633
rect 11336 24692 11388 24744
rect 8208 24556 8260 24608
rect 13728 24692 13780 24744
rect 15016 24735 15068 24744
rect 15016 24701 15025 24735
rect 15025 24701 15059 24735
rect 15059 24701 15068 24735
rect 15016 24692 15068 24701
rect 13268 24624 13320 24676
rect 15200 24624 15252 24676
rect 12992 24556 13044 24608
rect 17868 24760 17920 24812
rect 15660 24735 15712 24744
rect 15660 24701 15669 24735
rect 15669 24701 15703 24735
rect 15703 24701 15712 24735
rect 15660 24692 15712 24701
rect 16304 24735 16356 24744
rect 16304 24701 16313 24735
rect 16313 24701 16347 24735
rect 16347 24701 16356 24735
rect 16304 24692 16356 24701
rect 18052 24692 18104 24744
rect 18972 24692 19024 24744
rect 15752 24624 15804 24676
rect 20168 24692 20220 24744
rect 21640 24760 21692 24812
rect 21364 24667 21416 24676
rect 17500 24556 17552 24608
rect 18328 24556 18380 24608
rect 18696 24556 18748 24608
rect 21364 24633 21373 24667
rect 21373 24633 21407 24667
rect 21407 24633 21416 24667
rect 21364 24624 21416 24633
rect 21548 24692 21600 24744
rect 23480 24837 23489 24871
rect 23489 24837 23523 24871
rect 23523 24837 23532 24871
rect 23480 24828 23532 24837
rect 24400 24871 24452 24880
rect 24400 24837 24409 24871
rect 24409 24837 24443 24871
rect 24443 24837 24452 24871
rect 24400 24828 24452 24837
rect 25044 24871 25096 24880
rect 25044 24837 25053 24871
rect 25053 24837 25087 24871
rect 25087 24837 25096 24871
rect 25044 24828 25096 24837
rect 28264 24871 28316 24880
rect 28264 24837 28273 24871
rect 28273 24837 28307 24871
rect 28307 24837 28316 24871
rect 28264 24828 28316 24837
rect 28908 24828 28960 24880
rect 26056 24760 26108 24812
rect 26608 24760 26660 24812
rect 37556 24803 37608 24812
rect 37556 24769 37565 24803
rect 37565 24769 37599 24803
rect 37599 24769 37608 24803
rect 37556 24760 37608 24769
rect 23388 24735 23440 24744
rect 23388 24701 23397 24735
rect 23397 24701 23431 24735
rect 23431 24701 23440 24735
rect 23388 24692 23440 24701
rect 22744 24624 22796 24676
rect 26976 24692 27028 24744
rect 19984 24556 20036 24608
rect 21088 24556 21140 24608
rect 21640 24556 21692 24608
rect 22284 24556 22336 24608
rect 24584 24556 24636 24608
rect 37648 24599 37700 24608
rect 37648 24565 37657 24599
rect 37657 24565 37691 24599
rect 37691 24565 37700 24599
rect 37648 24556 37700 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4712 24352 4764 24404
rect 4896 24352 4948 24404
rect 5908 24352 5960 24404
rect 6000 24352 6052 24404
rect 7748 24352 7800 24404
rect 8668 24352 8720 24404
rect 9220 24352 9272 24404
rect 9496 24352 9548 24404
rect 13268 24352 13320 24404
rect 14648 24395 14700 24404
rect 14648 24361 14657 24395
rect 14657 24361 14691 24395
rect 14691 24361 14700 24395
rect 14648 24352 14700 24361
rect 15016 24352 15068 24404
rect 15660 24352 15712 24404
rect 17040 24352 17092 24404
rect 17776 24352 17828 24404
rect 19984 24352 20036 24404
rect 1860 24216 1912 24268
rect 3240 24216 3292 24268
rect 3424 24216 3476 24268
rect 6184 24216 6236 24268
rect 6736 24216 6788 24268
rect 8392 24216 8444 24268
rect 10968 24216 11020 24268
rect 11336 24216 11388 24268
rect 3700 24148 3752 24200
rect 4068 24148 4120 24200
rect 4620 24191 4672 24200
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 4620 24148 4672 24157
rect 6828 24191 6880 24200
rect 1584 24080 1636 24132
rect 3148 24080 3200 24132
rect 4804 24080 4856 24132
rect 2044 24012 2096 24064
rect 2136 24012 2188 24064
rect 5908 24012 5960 24064
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 17224 24284 17276 24336
rect 18880 24284 18932 24336
rect 19248 24284 19300 24336
rect 19708 24327 19760 24336
rect 19708 24293 19717 24327
rect 19717 24293 19751 24327
rect 19751 24293 19760 24327
rect 19708 24284 19760 24293
rect 13820 24216 13872 24268
rect 21180 24352 21232 24404
rect 21272 24352 21324 24404
rect 23204 24352 23256 24404
rect 28264 24352 28316 24404
rect 20536 24284 20588 24336
rect 20996 24284 21048 24336
rect 21548 24284 21600 24336
rect 21916 24284 21968 24336
rect 22376 24284 22428 24336
rect 25872 24284 25924 24336
rect 20720 24259 20772 24268
rect 20720 24225 20729 24259
rect 20729 24225 20763 24259
rect 20763 24225 20772 24259
rect 20720 24216 20772 24225
rect 23388 24216 23440 24268
rect 28908 24216 28960 24268
rect 38384 24216 38436 24268
rect 18696 24191 18748 24200
rect 7104 24123 7156 24132
rect 7104 24089 7113 24123
rect 7113 24089 7147 24123
rect 7147 24089 7156 24123
rect 7104 24080 7156 24089
rect 10048 24080 10100 24132
rect 7472 24012 7524 24064
rect 8760 24012 8812 24064
rect 11060 24012 11112 24064
rect 11244 24055 11296 24064
rect 11244 24021 11253 24055
rect 11253 24021 11287 24055
rect 11287 24021 11296 24055
rect 11244 24012 11296 24021
rect 11704 24080 11756 24132
rect 12072 24080 12124 24132
rect 12256 24080 12308 24132
rect 13268 24080 13320 24132
rect 14004 24080 14056 24132
rect 15108 24080 15160 24132
rect 13912 24012 13964 24064
rect 15016 24012 15068 24064
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 21824 24191 21876 24200
rect 16764 24123 16816 24132
rect 16764 24089 16773 24123
rect 16773 24089 16807 24123
rect 16807 24089 16816 24123
rect 16764 24080 16816 24089
rect 17592 24080 17644 24132
rect 17776 24123 17828 24132
rect 17776 24089 17785 24123
rect 17785 24089 17819 24123
rect 17819 24089 17828 24123
rect 17776 24080 17828 24089
rect 21824 24157 21833 24191
rect 21833 24157 21867 24191
rect 21867 24157 21876 24191
rect 21824 24148 21876 24157
rect 22100 24148 22152 24200
rect 22376 24148 22428 24200
rect 17040 24012 17092 24064
rect 17960 24012 18012 24064
rect 18052 24012 18104 24064
rect 20536 24080 20588 24132
rect 28172 24148 28224 24200
rect 33784 24148 33836 24200
rect 37464 24191 37516 24200
rect 37464 24157 37473 24191
rect 37473 24157 37507 24191
rect 37507 24157 37516 24191
rect 37464 24148 37516 24157
rect 37740 24191 37792 24200
rect 37740 24157 37749 24191
rect 37749 24157 37783 24191
rect 37783 24157 37792 24191
rect 37740 24148 37792 24157
rect 21916 24055 21968 24064
rect 21916 24021 21925 24055
rect 21925 24021 21959 24055
rect 21959 24021 21968 24055
rect 21916 24012 21968 24021
rect 22560 24055 22612 24064
rect 22560 24021 22569 24055
rect 22569 24021 22603 24055
rect 22603 24021 22612 24055
rect 22560 24012 22612 24021
rect 23664 24080 23716 24132
rect 24952 24080 25004 24132
rect 24676 24012 24728 24064
rect 29276 24080 29328 24132
rect 27344 24012 27396 24064
rect 30564 24012 30616 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 2964 23808 3016 23860
rect 4068 23808 4120 23860
rect 2872 23740 2924 23792
rect 4620 23808 4672 23860
rect 6276 23808 6328 23860
rect 6920 23740 6972 23792
rect 10232 23808 10284 23860
rect 11704 23808 11756 23860
rect 14188 23808 14240 23860
rect 14372 23808 14424 23860
rect 15200 23808 15252 23860
rect 15292 23808 15344 23860
rect 21824 23808 21876 23860
rect 23664 23851 23716 23860
rect 8944 23740 8996 23792
rect 10692 23740 10744 23792
rect 12072 23740 12124 23792
rect 13452 23740 13504 23792
rect 17868 23740 17920 23792
rect 19248 23740 19300 23792
rect 19432 23740 19484 23792
rect 19800 23783 19852 23792
rect 19800 23749 19809 23783
rect 19809 23749 19843 23783
rect 19843 23749 19852 23783
rect 19800 23740 19852 23749
rect 19892 23740 19944 23792
rect 21640 23740 21692 23792
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 3424 23604 3476 23656
rect 5080 23604 5132 23656
rect 5264 23604 5316 23656
rect 7932 23715 7984 23724
rect 7932 23681 7941 23715
rect 7941 23681 7975 23715
rect 7975 23681 7984 23715
rect 7932 23672 7984 23681
rect 11060 23672 11112 23724
rect 14188 23672 14240 23724
rect 6920 23604 6972 23656
rect 8300 23604 8352 23656
rect 8392 23604 8444 23656
rect 8852 23647 8904 23656
rect 8852 23613 8861 23647
rect 8861 23613 8895 23647
rect 8895 23613 8904 23647
rect 8852 23604 8904 23613
rect 8944 23604 8996 23656
rect 7288 23536 7340 23588
rect 7656 23536 7708 23588
rect 8116 23536 8168 23588
rect 10968 23604 11020 23656
rect 11428 23536 11480 23588
rect 11520 23536 11572 23588
rect 12164 23604 12216 23656
rect 12624 23604 12676 23656
rect 13820 23647 13872 23656
rect 13820 23613 13829 23647
rect 13829 23613 13863 23647
rect 13863 23613 13872 23647
rect 13820 23604 13872 23613
rect 14372 23647 14424 23656
rect 14372 23613 14381 23647
rect 14381 23613 14415 23647
rect 14415 23613 14424 23647
rect 14372 23604 14424 23613
rect 14556 23604 14608 23656
rect 13452 23536 13504 23588
rect 16028 23536 16080 23588
rect 2228 23468 2280 23520
rect 5632 23468 5684 23520
rect 6736 23468 6788 23520
rect 7104 23468 7156 23520
rect 7196 23468 7248 23520
rect 7748 23468 7800 23520
rect 9496 23468 9548 23520
rect 17224 23647 17276 23656
rect 17224 23613 17233 23647
rect 17233 23613 17267 23647
rect 17267 23613 17276 23647
rect 17224 23604 17276 23613
rect 17500 23647 17552 23656
rect 17500 23613 17509 23647
rect 17509 23613 17543 23647
rect 17543 23613 17552 23647
rect 17500 23604 17552 23613
rect 19800 23604 19852 23656
rect 16764 23536 16816 23588
rect 17868 23536 17920 23588
rect 17960 23536 18012 23588
rect 19432 23536 19484 23588
rect 20904 23604 20956 23656
rect 21088 23647 21140 23656
rect 21088 23613 21097 23647
rect 21097 23613 21131 23647
rect 21131 23613 21140 23647
rect 22284 23740 22336 23792
rect 23204 23740 23256 23792
rect 23664 23817 23673 23851
rect 23673 23817 23707 23851
rect 23707 23817 23716 23851
rect 23664 23808 23716 23817
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 25228 23808 25280 23860
rect 23940 23740 23992 23792
rect 27344 23783 27396 23792
rect 23572 23715 23624 23724
rect 23572 23681 23581 23715
rect 23581 23681 23615 23715
rect 23615 23681 23624 23715
rect 23572 23672 23624 23681
rect 27344 23749 27353 23783
rect 27353 23749 27387 23783
rect 27387 23749 27396 23783
rect 27344 23740 27396 23749
rect 28632 23783 28684 23792
rect 28632 23749 28641 23783
rect 28641 23749 28675 23783
rect 28675 23749 28684 23783
rect 28632 23740 28684 23749
rect 24492 23672 24544 23724
rect 21088 23604 21140 23613
rect 22744 23604 22796 23656
rect 22376 23536 22428 23588
rect 25044 23672 25096 23724
rect 26608 23672 26660 23724
rect 30564 23783 30616 23792
rect 30564 23749 30573 23783
rect 30573 23749 30607 23783
rect 30607 23749 30616 23783
rect 30564 23740 30616 23749
rect 30748 23740 30800 23792
rect 26516 23604 26568 23656
rect 27252 23647 27304 23656
rect 27252 23613 27261 23647
rect 27261 23613 27295 23647
rect 27295 23613 27304 23647
rect 27252 23604 27304 23613
rect 27896 23647 27948 23656
rect 27896 23613 27905 23647
rect 27905 23613 27939 23647
rect 27939 23613 27948 23647
rect 27896 23604 27948 23613
rect 28908 23604 28960 23656
rect 30656 23604 30708 23656
rect 30840 23647 30892 23656
rect 30840 23613 30849 23647
rect 30849 23613 30883 23647
rect 30883 23613 30892 23647
rect 30840 23604 30892 23613
rect 29736 23536 29788 23588
rect 16396 23468 16448 23520
rect 21272 23468 21324 23520
rect 23664 23468 23716 23520
rect 24952 23468 25004 23520
rect 26240 23511 26292 23520
rect 26240 23477 26249 23511
rect 26249 23477 26283 23511
rect 26283 23477 26292 23511
rect 26240 23468 26292 23477
rect 36084 23468 36136 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2228 23264 2280 23316
rect 2412 23264 2464 23316
rect 1860 23128 1912 23180
rect 1952 23128 2004 23180
rect 2412 23128 2464 23180
rect 5816 23264 5868 23316
rect 4252 23128 4304 23180
rect 4620 23128 4672 23180
rect 5448 23128 5500 23180
rect 8576 23196 8628 23248
rect 8668 23196 8720 23248
rect 8944 23196 8996 23248
rect 8024 23128 8076 23180
rect 8392 23128 8444 23180
rect 11244 23128 11296 23180
rect 11336 23128 11388 23180
rect 11980 23128 12032 23180
rect 12072 23128 12124 23180
rect 13268 23128 13320 23180
rect 20812 23264 20864 23316
rect 23388 23264 23440 23316
rect 30564 23264 30616 23316
rect 14372 23196 14424 23248
rect 14832 23196 14884 23248
rect 15476 23196 15528 23248
rect 16856 23196 16908 23248
rect 9312 23103 9364 23112
rect 1768 22992 1820 23044
rect 3608 22992 3660 23044
rect 9312 23069 9321 23103
rect 9321 23069 9355 23103
rect 9355 23069 9364 23103
rect 9312 23060 9364 23069
rect 10968 23060 11020 23112
rect 17224 23128 17276 23180
rect 17408 23171 17460 23180
rect 17408 23137 17417 23171
rect 17417 23137 17451 23171
rect 17451 23137 17460 23171
rect 17408 23128 17460 23137
rect 3332 22967 3384 22976
rect 3332 22933 3341 22967
rect 3341 22933 3375 22967
rect 3375 22933 3384 22967
rect 3332 22924 3384 22933
rect 6920 22992 6972 23044
rect 8392 22992 8444 23044
rect 11244 22992 11296 23044
rect 12256 22992 12308 23044
rect 13636 22992 13688 23044
rect 14096 22992 14148 23044
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 15016 22992 15068 23044
rect 16212 22992 16264 23044
rect 6552 22924 6604 22976
rect 9772 22924 9824 22976
rect 11612 22924 11664 22976
rect 15200 22924 15252 22976
rect 16488 22924 16540 22976
rect 16672 23035 16724 23044
rect 16672 23001 16681 23035
rect 16681 23001 16715 23035
rect 16715 23001 16724 23035
rect 16672 22992 16724 23001
rect 21456 23196 21508 23248
rect 21548 23196 21600 23248
rect 19892 23171 19944 23180
rect 19892 23137 19901 23171
rect 19901 23137 19935 23171
rect 19935 23137 19944 23171
rect 19892 23128 19944 23137
rect 20352 23128 20404 23180
rect 22008 23128 22060 23180
rect 24676 23171 24728 23180
rect 24676 23137 24685 23171
rect 24685 23137 24719 23171
rect 24719 23137 24728 23171
rect 24676 23128 24728 23137
rect 28540 23196 28592 23248
rect 27896 23128 27948 23180
rect 28632 23171 28684 23180
rect 28632 23137 28641 23171
rect 28641 23137 28675 23171
rect 28675 23137 28684 23171
rect 28632 23128 28684 23137
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 30288 23060 30340 23112
rect 18328 23035 18380 23044
rect 18328 23001 18337 23035
rect 18337 23001 18371 23035
rect 18371 23001 18380 23035
rect 18880 23035 18932 23044
rect 18328 22992 18380 23001
rect 18880 23001 18889 23035
rect 18889 23001 18923 23035
rect 18923 23001 18932 23035
rect 18880 22992 18932 23001
rect 20904 23035 20956 23044
rect 20904 23001 20913 23035
rect 20913 23001 20947 23035
rect 20947 23001 20956 23035
rect 20904 22992 20956 23001
rect 21548 22992 21600 23044
rect 21916 23035 21968 23044
rect 21916 23001 21925 23035
rect 21925 23001 21959 23035
rect 21959 23001 21968 23035
rect 21916 22992 21968 23001
rect 22560 22992 22612 23044
rect 22744 22992 22796 23044
rect 23572 22992 23624 23044
rect 24952 22992 25004 23044
rect 25504 22992 25556 23044
rect 27988 22992 28040 23044
rect 28356 23035 28408 23044
rect 28356 23001 28365 23035
rect 28365 23001 28399 23035
rect 28399 23001 28408 23035
rect 28356 22992 28408 23001
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 1676 22720 1728 22772
rect 4160 22720 4212 22772
rect 5724 22720 5776 22772
rect 6460 22720 6512 22772
rect 1308 22652 1360 22704
rect 3516 22652 3568 22704
rect 4528 22652 4580 22704
rect 6644 22652 6696 22704
rect 4160 22627 4212 22636
rect 4160 22593 4169 22627
rect 4169 22593 4203 22627
rect 4203 22593 4212 22627
rect 4160 22584 4212 22593
rect 5540 22584 5592 22636
rect 7288 22627 7340 22636
rect 7288 22593 7297 22627
rect 7297 22593 7331 22627
rect 7331 22593 7340 22627
rect 10968 22720 11020 22772
rect 11244 22720 11296 22772
rect 12440 22720 12492 22772
rect 12808 22720 12860 22772
rect 14004 22720 14056 22772
rect 9588 22652 9640 22704
rect 9772 22652 9824 22704
rect 10048 22652 10100 22704
rect 12256 22652 12308 22704
rect 12624 22652 12676 22704
rect 13544 22652 13596 22704
rect 17684 22720 17736 22772
rect 14280 22695 14332 22704
rect 14280 22661 14289 22695
rect 14289 22661 14323 22695
rect 14323 22661 14332 22695
rect 14280 22652 14332 22661
rect 14648 22652 14700 22704
rect 15936 22652 15988 22704
rect 7288 22584 7340 22593
rect 9312 22584 9364 22636
rect 9956 22584 10008 22636
rect 10232 22627 10284 22636
rect 10232 22593 10241 22627
rect 10241 22593 10275 22627
rect 10275 22593 10284 22627
rect 10232 22584 10284 22593
rect 15292 22584 15344 22636
rect 15752 22584 15804 22636
rect 16672 22584 16724 22636
rect 16764 22584 16816 22636
rect 1676 22516 1728 22568
rect 2136 22559 2188 22568
rect 2136 22525 2145 22559
rect 2145 22525 2179 22559
rect 2179 22525 2188 22559
rect 2136 22516 2188 22525
rect 2780 22516 2832 22568
rect 7380 22516 7432 22568
rect 8024 22559 8076 22568
rect 8024 22525 8033 22559
rect 8033 22525 8067 22559
rect 8067 22525 8076 22559
rect 8024 22516 8076 22525
rect 8576 22516 8628 22568
rect 9220 22516 9272 22568
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 3240 22448 3292 22500
rect 5540 22448 5592 22500
rect 7472 22448 7524 22500
rect 9128 22448 9180 22500
rect 13176 22516 13228 22568
rect 13544 22516 13596 22568
rect 13912 22516 13964 22568
rect 14556 22559 14608 22568
rect 1952 22380 2004 22432
rect 7288 22380 7340 22432
rect 14096 22380 14148 22432
rect 14556 22525 14565 22559
rect 14565 22525 14599 22559
rect 14599 22525 14608 22559
rect 14556 22516 14608 22525
rect 14464 22448 14516 22500
rect 16856 22448 16908 22500
rect 18880 22720 18932 22772
rect 22100 22720 22152 22772
rect 18328 22652 18380 22704
rect 18696 22652 18748 22704
rect 18696 22516 18748 22568
rect 20352 22584 20404 22636
rect 20812 22652 20864 22704
rect 23664 22652 23716 22704
rect 23940 22695 23992 22704
rect 23940 22661 23949 22695
rect 23949 22661 23983 22695
rect 23983 22661 23992 22695
rect 23940 22652 23992 22661
rect 17132 22448 17184 22500
rect 17592 22448 17644 22500
rect 14648 22380 14700 22432
rect 14832 22380 14884 22432
rect 16304 22380 16356 22432
rect 16580 22380 16632 22432
rect 22376 22516 22428 22568
rect 22560 22559 22612 22568
rect 22560 22525 22569 22559
rect 22569 22525 22603 22559
rect 22603 22525 22612 22559
rect 22560 22516 22612 22525
rect 25964 22695 26016 22704
rect 25964 22661 25973 22695
rect 25973 22661 26007 22695
rect 26007 22661 26016 22695
rect 25964 22652 26016 22661
rect 26240 22652 26292 22704
rect 26700 22720 26752 22772
rect 28080 22763 28132 22772
rect 28080 22729 28089 22763
rect 28089 22729 28123 22763
rect 28123 22729 28132 22763
rect 28080 22720 28132 22729
rect 28356 22652 28408 22704
rect 29368 22695 29420 22704
rect 29368 22661 29377 22695
rect 29377 22661 29411 22695
rect 29411 22661 29420 22695
rect 29368 22652 29420 22661
rect 27068 22584 27120 22636
rect 29000 22584 29052 22636
rect 37556 22584 37608 22636
rect 38016 22627 38068 22636
rect 38016 22593 38025 22627
rect 38025 22593 38059 22627
rect 38059 22593 38068 22627
rect 38016 22584 38068 22593
rect 24860 22559 24912 22568
rect 24860 22525 24869 22559
rect 24869 22525 24903 22559
rect 24903 22525 24912 22559
rect 29276 22559 29328 22568
rect 24860 22516 24912 22525
rect 20812 22448 20864 22500
rect 21916 22448 21968 22500
rect 22192 22448 22244 22500
rect 26516 22491 26568 22500
rect 20628 22380 20680 22432
rect 21272 22380 21324 22432
rect 21456 22380 21508 22432
rect 26516 22457 26525 22491
rect 26525 22457 26559 22491
rect 26559 22457 26568 22491
rect 26516 22448 26568 22457
rect 29276 22525 29285 22559
rect 29285 22525 29319 22559
rect 29319 22525 29328 22559
rect 29276 22516 29328 22525
rect 29552 22559 29604 22568
rect 29552 22525 29561 22559
rect 29561 22525 29595 22559
rect 29595 22525 29604 22559
rect 29552 22516 29604 22525
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 23388 22380 23440 22432
rect 26608 22380 26660 22432
rect 29184 22380 29236 22432
rect 29552 22380 29604 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2412 22176 2464 22228
rect 6184 22176 6236 22228
rect 5632 22108 5684 22160
rect 9128 22176 9180 22228
rect 9220 22176 9272 22228
rect 11152 22176 11204 22228
rect 1676 22083 1728 22092
rect 1676 22049 1685 22083
rect 1685 22049 1719 22083
rect 1719 22049 1728 22083
rect 1676 22040 1728 22049
rect 1952 22083 2004 22092
rect 1952 22049 1961 22083
rect 1961 22049 1995 22083
rect 1995 22049 2004 22083
rect 1952 22040 2004 22049
rect 3516 22040 3568 22092
rect 3976 22054 4028 22106
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 5908 22040 5960 22092
rect 5632 21972 5684 22024
rect 4436 21904 4488 21956
rect 6276 22083 6328 22092
rect 6276 22049 6285 22083
rect 6285 22049 6319 22083
rect 6319 22049 6328 22083
rect 6276 22040 6328 22049
rect 7012 22040 7064 22092
rect 8668 22040 8720 22092
rect 10508 22108 10560 22160
rect 14464 22176 14516 22228
rect 9680 22040 9732 22092
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 7564 21972 7616 22024
rect 6276 21904 6328 21956
rect 8208 21904 8260 21956
rect 9404 21904 9456 21956
rect 11612 22083 11664 22092
rect 11612 22049 11621 22083
rect 11621 22049 11655 22083
rect 11655 22049 11664 22083
rect 11612 22040 11664 22049
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10968 21972 11020 22024
rect 12716 21972 12768 22024
rect 13176 22040 13228 22092
rect 14188 22040 14240 22092
rect 13820 21972 13872 22024
rect 15016 21972 15068 22024
rect 3240 21836 3292 21888
rect 5816 21879 5868 21888
rect 5816 21845 5825 21879
rect 5825 21845 5859 21879
rect 5859 21845 5868 21879
rect 5816 21836 5868 21845
rect 7196 21836 7248 21888
rect 8668 21836 8720 21888
rect 11612 21904 11664 21956
rect 16764 22176 16816 22228
rect 15200 22108 15252 22160
rect 16028 22040 16080 22092
rect 16488 22108 16540 22160
rect 17500 22176 17552 22228
rect 18604 22176 18656 22228
rect 20076 22219 20128 22228
rect 20076 22185 20085 22219
rect 20085 22185 20119 22219
rect 20119 22185 20128 22219
rect 20076 22176 20128 22185
rect 20444 22176 20496 22228
rect 22928 22176 22980 22228
rect 23940 22176 23992 22228
rect 17224 22108 17276 22160
rect 26424 22108 26476 22160
rect 27068 22108 27120 22160
rect 30656 22108 30708 22160
rect 17224 21972 17276 22024
rect 17960 21972 18012 22024
rect 19432 22040 19484 22092
rect 21364 22083 21416 22092
rect 21364 22049 21373 22083
rect 21373 22049 21407 22083
rect 21407 22049 21416 22083
rect 21364 22040 21416 22049
rect 22284 22083 22336 22092
rect 22284 22049 22293 22083
rect 22293 22049 22327 22083
rect 22327 22049 22336 22083
rect 22284 22040 22336 22049
rect 23572 22040 23624 22092
rect 23756 22040 23808 22092
rect 26516 22040 26568 22092
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 15384 21947 15436 21956
rect 12440 21836 12492 21888
rect 15384 21913 15404 21947
rect 15404 21913 15436 21947
rect 15384 21904 15436 21913
rect 15936 21947 15988 21956
rect 15936 21913 15945 21947
rect 15945 21913 15979 21947
rect 15979 21913 15988 21947
rect 15936 21904 15988 21913
rect 16488 21947 16540 21956
rect 16488 21913 16497 21947
rect 16497 21913 16531 21947
rect 16531 21913 16540 21947
rect 16488 21904 16540 21913
rect 16580 21947 16632 21956
rect 16580 21913 16589 21947
rect 16589 21913 16623 21947
rect 16623 21913 16632 21947
rect 16580 21904 16632 21913
rect 16764 21904 16816 21956
rect 22192 22015 22244 22024
rect 22192 21981 22201 22015
rect 22201 21981 22235 22015
rect 22235 21981 22244 22015
rect 22192 21972 22244 21981
rect 24492 21972 24544 22024
rect 21272 21904 21324 21956
rect 22100 21904 22152 21956
rect 23204 21904 23256 21956
rect 23388 21947 23440 21956
rect 23388 21913 23397 21947
rect 23397 21913 23431 21947
rect 23431 21913 23440 21947
rect 23388 21904 23440 21913
rect 24216 21904 24268 21956
rect 26884 22015 26936 22024
rect 26884 21981 26893 22015
rect 26893 21981 26927 22015
rect 26927 21981 26936 22015
rect 26884 21972 26936 21981
rect 28632 22040 28684 22092
rect 33784 21972 33836 22024
rect 38292 22015 38344 22024
rect 38292 21981 38301 22015
rect 38301 21981 38335 22015
rect 38335 21981 38344 22015
rect 38292 21972 38344 21981
rect 13176 21836 13228 21888
rect 15660 21836 15712 21888
rect 15844 21836 15896 21888
rect 16948 21836 17000 21888
rect 17040 21836 17092 21888
rect 17408 21836 17460 21888
rect 18788 21879 18840 21888
rect 18788 21845 18797 21879
rect 18797 21845 18831 21879
rect 18831 21845 18840 21879
rect 18788 21836 18840 21845
rect 22652 21836 22704 21888
rect 32680 21904 32732 21956
rect 33600 21836 33652 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2504 21632 2556 21684
rect 3240 21632 3292 21684
rect 3332 21632 3384 21684
rect 5080 21632 5132 21684
rect 5356 21632 5408 21684
rect 6460 21632 6512 21684
rect 1860 21564 1912 21616
rect 1584 21539 1636 21548
rect 1584 21505 1593 21539
rect 1593 21505 1627 21539
rect 1627 21505 1636 21539
rect 1584 21496 1636 21505
rect 5172 21564 5224 21616
rect 6644 21564 6696 21616
rect 7012 21564 7064 21616
rect 9220 21632 9272 21684
rect 7196 21496 7248 21548
rect 8852 21564 8904 21616
rect 11244 21632 11296 21684
rect 11612 21632 11664 21684
rect 1952 21428 2004 21480
rect 2504 21428 2556 21480
rect 4528 21428 4580 21480
rect 4712 21428 4764 21480
rect 5172 21428 5224 21480
rect 4436 21360 4488 21412
rect 7472 21428 7524 21480
rect 6828 21360 6880 21412
rect 8392 21428 8444 21480
rect 9956 21564 10008 21616
rect 15384 21632 15436 21684
rect 10232 21496 10284 21548
rect 10600 21496 10652 21548
rect 11980 21564 12032 21616
rect 12256 21564 12308 21616
rect 14096 21564 14148 21616
rect 18696 21632 18748 21684
rect 18788 21632 18840 21684
rect 21272 21675 21324 21684
rect 15844 21564 15896 21616
rect 15016 21496 15068 21548
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 17132 21539 17184 21548
rect 16304 21496 16356 21505
rect 17132 21505 17141 21539
rect 17141 21505 17175 21539
rect 17175 21505 17184 21539
rect 17132 21496 17184 21505
rect 9956 21428 10008 21480
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 12900 21428 12952 21480
rect 12992 21428 13044 21480
rect 14096 21428 14148 21480
rect 14832 21428 14884 21480
rect 15844 21428 15896 21480
rect 16028 21428 16080 21480
rect 18144 21564 18196 21616
rect 18512 21607 18564 21616
rect 18512 21573 18521 21607
rect 18521 21573 18555 21607
rect 18555 21573 18564 21607
rect 18512 21564 18564 21573
rect 17776 21539 17828 21548
rect 17776 21505 17785 21539
rect 17785 21505 17819 21539
rect 17819 21505 17828 21539
rect 17776 21496 17828 21505
rect 20168 21564 20220 21616
rect 21272 21641 21281 21675
rect 21281 21641 21315 21675
rect 21315 21641 21324 21675
rect 21272 21632 21324 21641
rect 23480 21632 23532 21684
rect 24216 21675 24268 21684
rect 24216 21641 24225 21675
rect 24225 21641 24259 21675
rect 24259 21641 24268 21675
rect 24216 21632 24268 21641
rect 24860 21632 24912 21684
rect 30748 21632 30800 21684
rect 38200 21675 38252 21684
rect 38200 21641 38209 21675
rect 38209 21641 38243 21675
rect 38243 21641 38252 21675
rect 38200 21632 38252 21641
rect 21916 21564 21968 21616
rect 21180 21539 21232 21548
rect 19340 21428 19392 21480
rect 5632 21292 5684 21344
rect 10508 21360 10560 21412
rect 13912 21360 13964 21412
rect 11796 21292 11848 21344
rect 12440 21292 12492 21344
rect 12532 21292 12584 21344
rect 18788 21360 18840 21412
rect 18144 21292 18196 21344
rect 21180 21505 21189 21539
rect 21189 21505 21223 21539
rect 21223 21505 21232 21539
rect 21180 21496 21232 21505
rect 21548 21496 21600 21548
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 23020 21496 23072 21548
rect 23480 21539 23532 21548
rect 23480 21505 23489 21539
rect 23489 21505 23523 21539
rect 23523 21505 23532 21539
rect 23480 21496 23532 21505
rect 23848 21496 23900 21548
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 24216 21496 24268 21548
rect 28908 21607 28960 21616
rect 28908 21573 28917 21607
rect 28917 21573 28951 21607
rect 28951 21573 28960 21607
rect 28908 21564 28960 21573
rect 29000 21564 29052 21616
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 37556 21496 37608 21548
rect 38108 21539 38160 21548
rect 38108 21505 38117 21539
rect 38117 21505 38151 21539
rect 38151 21505 38160 21539
rect 38108 21496 38160 21505
rect 20260 21471 20312 21480
rect 20260 21437 20269 21471
rect 20269 21437 20303 21471
rect 20303 21437 20312 21471
rect 20260 21428 20312 21437
rect 20720 21428 20772 21480
rect 22100 21428 22152 21480
rect 22192 21428 22244 21480
rect 21088 21292 21140 21344
rect 22192 21292 22244 21344
rect 22468 21292 22520 21344
rect 25320 21292 25372 21344
rect 27436 21428 27488 21480
rect 28356 21428 28408 21480
rect 29276 21360 29328 21412
rect 28816 21292 28868 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1124 21088 1176 21140
rect 3332 21063 3384 21072
rect 3332 21029 3341 21063
rect 3341 21029 3375 21063
rect 3375 21029 3384 21063
rect 3332 21020 3384 21029
rect 1860 20952 1912 21004
rect 5356 21088 5408 21140
rect 4068 20952 4120 21004
rect 6368 20952 6420 21004
rect 6460 20952 6512 21004
rect 8208 20952 8260 21004
rect 8392 21088 8444 21140
rect 9128 21020 9180 21072
rect 10416 21020 10468 21072
rect 12440 21088 12492 21140
rect 16304 21088 16356 21140
rect 16580 21088 16632 21140
rect 3792 20816 3844 20868
rect 5080 20816 5132 20868
rect 6552 20816 6604 20868
rect 7012 20816 7064 20868
rect 7564 20816 7616 20868
rect 8668 20884 8720 20936
rect 10324 20952 10376 21004
rect 10600 20884 10652 20936
rect 10968 20927 11020 20936
rect 10968 20893 10977 20927
rect 10977 20893 11011 20927
rect 11011 20893 11020 20927
rect 10968 20884 11020 20893
rect 12532 20884 12584 20936
rect 13728 21020 13780 21072
rect 13636 20952 13688 21004
rect 17132 21020 17184 21072
rect 18696 21020 18748 21072
rect 19340 21020 19392 21072
rect 19432 21020 19484 21072
rect 20536 21088 20588 21140
rect 21456 21088 21508 21140
rect 22192 21088 22244 21140
rect 25504 21088 25556 21140
rect 28816 21088 28868 21140
rect 29368 21088 29420 21140
rect 13728 20884 13780 20936
rect 15476 20884 15528 20936
rect 16120 20884 16172 20936
rect 16396 20884 16448 20936
rect 18512 20952 18564 21004
rect 17960 20884 18012 20936
rect 2780 20748 2832 20800
rect 3976 20748 4028 20800
rect 8852 20816 8904 20868
rect 9036 20816 9088 20868
rect 9220 20859 9272 20868
rect 9220 20825 9229 20859
rect 9229 20825 9263 20859
rect 9263 20825 9272 20859
rect 9220 20816 9272 20825
rect 8116 20748 8168 20800
rect 10324 20816 10376 20868
rect 11152 20816 11204 20868
rect 11704 20816 11756 20868
rect 12716 20816 12768 20868
rect 9772 20748 9824 20800
rect 9956 20748 10008 20800
rect 10048 20748 10100 20800
rect 10876 20748 10928 20800
rect 11428 20748 11480 20800
rect 12532 20748 12584 20800
rect 13084 20748 13136 20800
rect 14188 20816 14240 20868
rect 14464 20859 14516 20868
rect 14464 20825 14473 20859
rect 14473 20825 14507 20859
rect 14507 20825 14516 20859
rect 14464 20816 14516 20825
rect 15292 20816 15344 20868
rect 15384 20859 15436 20868
rect 15384 20825 15393 20859
rect 15393 20825 15427 20859
rect 15427 20825 15436 20859
rect 15384 20816 15436 20825
rect 16856 20816 16908 20868
rect 17132 20859 17184 20868
rect 17132 20825 17141 20859
rect 17141 20825 17175 20859
rect 17175 20825 17184 20859
rect 17132 20816 17184 20825
rect 17868 20816 17920 20868
rect 19800 20952 19852 21004
rect 20720 20952 20772 21004
rect 21916 20952 21968 21004
rect 22928 20952 22980 21004
rect 22100 20884 22152 20936
rect 22560 20884 22612 20936
rect 22836 20927 22888 20936
rect 22836 20893 22845 20927
rect 22845 20893 22879 20927
rect 22879 20893 22888 20927
rect 22836 20884 22888 20893
rect 23848 21020 23900 21072
rect 24492 21020 24544 21072
rect 25780 21063 25832 21072
rect 25780 21029 25789 21063
rect 25789 21029 25823 21063
rect 25823 21029 25832 21063
rect 25780 21020 25832 21029
rect 25964 21020 26016 21072
rect 27252 20952 27304 21004
rect 28632 20952 28684 21004
rect 29644 20952 29696 21004
rect 26240 20884 26292 20936
rect 27804 20927 27856 20936
rect 27804 20893 27813 20927
rect 27813 20893 27847 20927
rect 27847 20893 27856 20927
rect 27804 20884 27856 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 14832 20748 14884 20800
rect 19156 20748 19208 20800
rect 19524 20816 19576 20868
rect 19800 20816 19852 20868
rect 20352 20816 20404 20868
rect 23020 20816 23072 20868
rect 24860 20816 24912 20868
rect 25320 20859 25372 20868
rect 25320 20825 25329 20859
rect 25329 20825 25363 20859
rect 25363 20825 25372 20859
rect 25320 20816 25372 20825
rect 25964 20816 26016 20868
rect 21456 20748 21508 20800
rect 22192 20748 22244 20800
rect 22376 20748 22428 20800
rect 24768 20748 24820 20800
rect 30380 20816 30432 20868
rect 29276 20748 29328 20800
rect 29552 20748 29604 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1216 20544 1268 20596
rect 3884 20476 3936 20528
rect 1860 20451 1912 20460
rect 1860 20417 1869 20451
rect 1869 20417 1903 20451
rect 1903 20417 1912 20451
rect 1860 20408 1912 20417
rect 3332 20340 3384 20392
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 4068 20544 4120 20596
rect 4988 20519 5040 20528
rect 4988 20485 4997 20519
rect 4997 20485 5031 20519
rect 5031 20485 5040 20519
rect 4988 20476 5040 20485
rect 5448 20476 5500 20528
rect 7196 20476 7248 20528
rect 9404 20476 9456 20528
rect 10232 20544 10284 20596
rect 12900 20544 12952 20596
rect 14832 20544 14884 20596
rect 15292 20544 15344 20596
rect 10784 20476 10836 20528
rect 11980 20476 12032 20528
rect 13360 20476 13412 20528
rect 13452 20476 13504 20528
rect 13912 20476 13964 20528
rect 16580 20544 16632 20596
rect 17132 20544 17184 20596
rect 18696 20544 18748 20596
rect 19248 20544 19300 20596
rect 19432 20544 19484 20596
rect 19892 20544 19944 20596
rect 18788 20519 18840 20528
rect 18788 20485 18797 20519
rect 18797 20485 18831 20519
rect 18831 20485 18840 20519
rect 18788 20476 18840 20485
rect 20076 20476 20128 20528
rect 6920 20408 6972 20460
rect 7288 20340 7340 20392
rect 8300 20340 8352 20392
rect 9220 20408 9272 20460
rect 3516 20272 3568 20324
rect 9956 20340 10008 20392
rect 10968 20340 11020 20392
rect 12072 20340 12124 20392
rect 12532 20340 12584 20392
rect 17960 20451 18012 20460
rect 13820 20340 13872 20392
rect 14648 20340 14700 20392
rect 15292 20383 15344 20392
rect 15292 20349 15301 20383
rect 15301 20349 15335 20383
rect 15335 20349 15344 20383
rect 15292 20340 15344 20349
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 16304 20340 16356 20392
rect 17224 20340 17276 20392
rect 17960 20417 17969 20451
rect 17969 20417 18003 20451
rect 18003 20417 18012 20451
rect 17960 20408 18012 20417
rect 19616 20408 19668 20460
rect 26332 20544 26384 20596
rect 28908 20544 28960 20596
rect 20444 20476 20496 20528
rect 22376 20519 22428 20528
rect 22376 20485 22385 20519
rect 22385 20485 22419 20519
rect 22419 20485 22428 20519
rect 22376 20476 22428 20485
rect 22468 20476 22520 20528
rect 20352 20398 20404 20450
rect 17500 20340 17552 20392
rect 18696 20383 18748 20392
rect 18696 20349 18705 20383
rect 18705 20349 18739 20383
rect 18739 20349 18748 20383
rect 18696 20340 18748 20349
rect 18788 20340 18840 20392
rect 21732 20408 21784 20460
rect 23020 20408 23072 20460
rect 23480 20408 23532 20460
rect 1768 20204 1820 20256
rect 3884 20204 3936 20256
rect 11612 20272 11664 20324
rect 6000 20204 6052 20256
rect 19984 20272 20036 20324
rect 21180 20340 21232 20392
rect 21824 20340 21876 20392
rect 22008 20340 22060 20392
rect 22284 20383 22336 20392
rect 22284 20349 22293 20383
rect 22293 20349 22327 20383
rect 22327 20349 22336 20383
rect 22284 20340 22336 20349
rect 24124 20408 24176 20460
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 26148 20476 26200 20528
rect 27804 20476 27856 20528
rect 27896 20476 27948 20528
rect 29460 20476 29512 20528
rect 23848 20340 23900 20392
rect 25688 20383 25740 20392
rect 25688 20349 25697 20383
rect 25697 20349 25731 20383
rect 25731 20349 25740 20383
rect 25688 20340 25740 20349
rect 25964 20340 26016 20392
rect 27068 20408 27120 20460
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 29736 20408 29788 20460
rect 28448 20340 28500 20392
rect 22836 20315 22888 20324
rect 22836 20281 22845 20315
rect 22845 20281 22879 20315
rect 22879 20281 22888 20315
rect 22836 20272 22888 20281
rect 22928 20272 22980 20324
rect 25780 20272 25832 20324
rect 30012 20272 30064 20324
rect 15844 20204 15896 20256
rect 17868 20204 17920 20256
rect 17960 20204 18012 20256
rect 18512 20204 18564 20256
rect 19064 20204 19116 20256
rect 19248 20204 19300 20256
rect 20720 20204 20772 20256
rect 21272 20204 21324 20256
rect 23020 20204 23072 20256
rect 23480 20247 23532 20256
rect 23480 20213 23489 20247
rect 23489 20213 23523 20247
rect 23523 20213 23532 20247
rect 23480 20204 23532 20213
rect 24308 20204 24360 20256
rect 24492 20204 24544 20256
rect 27068 20204 27120 20256
rect 27344 20204 27396 20256
rect 29736 20247 29788 20256
rect 29736 20213 29745 20247
rect 29745 20213 29779 20247
rect 29779 20213 29788 20247
rect 29736 20204 29788 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2964 20000 3016 20052
rect 3700 20000 3752 20052
rect 3884 20000 3936 20052
rect 11704 20000 11756 20052
rect 12900 20000 12952 20052
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 13636 20000 13688 20009
rect 13912 20000 13964 20052
rect 16764 20000 16816 20052
rect 16948 20000 17000 20052
rect 18788 20000 18840 20052
rect 18880 20000 18932 20052
rect 19616 20000 19668 20052
rect 21088 20043 21140 20052
rect 1860 19864 1912 19916
rect 2872 19864 2924 19916
rect 3424 19864 3476 19916
rect 5356 19864 5408 19916
rect 6920 19864 6972 19916
rect 9220 19864 9272 19916
rect 10232 19907 10284 19916
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 10232 19873 10241 19907
rect 10241 19873 10275 19907
rect 10275 19873 10284 19907
rect 10232 19864 10284 19873
rect 10876 19907 10928 19916
rect 10876 19873 10885 19907
rect 10885 19873 10919 19907
rect 10919 19873 10928 19907
rect 10876 19864 10928 19873
rect 12440 19932 12492 19984
rect 12532 19932 12584 19984
rect 10600 19796 10652 19848
rect 12716 19864 12768 19916
rect 16948 19864 17000 19916
rect 17316 19864 17368 19916
rect 19432 19932 19484 19984
rect 19892 19932 19944 19984
rect 20352 19932 20404 19984
rect 20812 19932 20864 19984
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 22468 20000 22520 20052
rect 23388 20000 23440 20052
rect 23664 20043 23716 20052
rect 23664 20009 23673 20043
rect 23673 20009 23707 20043
rect 23707 20009 23716 20043
rect 23664 20000 23716 20009
rect 24308 19932 24360 19984
rect 25596 19932 25648 19984
rect 27712 19975 27764 19984
rect 27712 19941 27721 19975
rect 27721 19941 27755 19975
rect 27755 19941 27764 19975
rect 27712 19932 27764 19941
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 13728 19796 13780 19848
rect 19616 19864 19668 19916
rect 20076 19864 20128 19916
rect 2596 19728 2648 19780
rect 2688 19660 2740 19712
rect 4620 19728 4672 19780
rect 5448 19728 5500 19780
rect 5816 19728 5868 19780
rect 7840 19728 7892 19780
rect 9036 19728 9088 19780
rect 4712 19660 4764 19712
rect 8668 19660 8720 19712
rect 9404 19728 9456 19780
rect 10876 19728 10928 19780
rect 11244 19728 11296 19780
rect 9496 19660 9548 19712
rect 12716 19728 12768 19780
rect 13360 19728 13412 19780
rect 13452 19728 13504 19780
rect 13912 19728 13964 19780
rect 14096 19728 14148 19780
rect 14924 19728 14976 19780
rect 15568 19728 15620 19780
rect 15844 19728 15896 19780
rect 18420 19796 18472 19848
rect 17592 19771 17644 19780
rect 17592 19737 17601 19771
rect 17601 19737 17635 19771
rect 17635 19737 17644 19771
rect 17592 19728 17644 19737
rect 17684 19771 17736 19780
rect 17684 19737 17693 19771
rect 17693 19737 17727 19771
rect 17727 19737 17736 19771
rect 17684 19728 17736 19737
rect 12532 19660 12584 19712
rect 13636 19660 13688 19712
rect 13728 19660 13780 19712
rect 18788 19703 18840 19712
rect 18788 19669 18797 19703
rect 18797 19669 18831 19703
rect 18831 19669 18840 19703
rect 18788 19660 18840 19669
rect 18972 19728 19024 19780
rect 19340 19728 19392 19780
rect 25688 19864 25740 19916
rect 26424 19864 26476 19916
rect 20904 19796 20956 19848
rect 21180 19796 21232 19848
rect 21640 19839 21692 19848
rect 21272 19728 21324 19780
rect 21640 19805 21649 19839
rect 21649 19805 21683 19839
rect 21683 19805 21692 19839
rect 21640 19796 21692 19805
rect 23756 19796 23808 19848
rect 24216 19796 24268 19848
rect 24492 19796 24544 19848
rect 22468 19771 22520 19780
rect 21180 19660 21232 19712
rect 22468 19737 22477 19771
rect 22477 19737 22511 19771
rect 22511 19737 22520 19771
rect 22468 19728 22520 19737
rect 22560 19771 22612 19780
rect 22560 19737 22569 19771
rect 22569 19737 22603 19771
rect 22603 19737 22612 19771
rect 22560 19728 22612 19737
rect 22928 19728 22980 19780
rect 23664 19728 23716 19780
rect 25044 19796 25096 19848
rect 27252 19796 27304 19848
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 37832 19796 37884 19848
rect 38292 19839 38344 19848
rect 38292 19805 38301 19839
rect 38301 19805 38335 19839
rect 38335 19805 38344 19839
rect 38292 19796 38344 19805
rect 24860 19728 24912 19780
rect 29920 19771 29972 19780
rect 29920 19737 29929 19771
rect 29929 19737 29963 19771
rect 29963 19737 29972 19771
rect 29920 19728 29972 19737
rect 30012 19771 30064 19780
rect 30012 19737 30021 19771
rect 30021 19737 30055 19771
rect 30055 19737 30064 19771
rect 30012 19728 30064 19737
rect 30380 19728 30432 19780
rect 31392 19728 31444 19780
rect 23388 19660 23440 19712
rect 25780 19703 25832 19712
rect 25780 19669 25789 19703
rect 25789 19669 25823 19703
rect 25823 19669 25832 19703
rect 25780 19660 25832 19669
rect 26424 19703 26476 19712
rect 26424 19669 26433 19703
rect 26433 19669 26467 19703
rect 26467 19669 26476 19703
rect 26424 19660 26476 19669
rect 27068 19703 27120 19712
rect 27068 19669 27077 19703
rect 27077 19669 27111 19703
rect 27111 19669 27120 19703
rect 27068 19660 27120 19669
rect 27804 19660 27856 19712
rect 28540 19660 28592 19712
rect 29092 19660 29144 19712
rect 31484 19660 31536 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1952 19456 2004 19508
rect 11244 19456 11296 19508
rect 6736 19388 6788 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 5356 19320 5408 19372
rect 7748 19388 7800 19440
rect 9496 19431 9548 19440
rect 9496 19397 9505 19431
rect 9505 19397 9539 19431
rect 9539 19397 9548 19431
rect 9496 19388 9548 19397
rect 10140 19431 10192 19440
rect 10140 19397 10149 19431
rect 10149 19397 10183 19431
rect 10183 19397 10192 19431
rect 10140 19388 10192 19397
rect 10232 19388 10284 19440
rect 10600 19388 10652 19440
rect 11612 19388 11664 19440
rect 13176 19456 13228 19508
rect 13452 19456 13504 19508
rect 12256 19431 12308 19440
rect 12256 19397 12265 19431
rect 12265 19397 12299 19431
rect 12299 19397 12308 19431
rect 12256 19388 12308 19397
rect 12440 19388 12492 19440
rect 13544 19388 13596 19440
rect 14924 19456 14976 19508
rect 13820 19431 13872 19440
rect 13820 19397 13829 19431
rect 13829 19397 13863 19431
rect 13863 19397 13872 19431
rect 13820 19388 13872 19397
rect 14556 19388 14608 19440
rect 14832 19388 14884 19440
rect 16028 19456 16080 19508
rect 16488 19456 16540 19508
rect 15568 19388 15620 19440
rect 16948 19431 17000 19440
rect 16948 19397 16957 19431
rect 16957 19397 16991 19431
rect 16991 19397 17000 19431
rect 16948 19388 17000 19397
rect 18512 19456 18564 19508
rect 17224 19388 17276 19440
rect 18972 19456 19024 19508
rect 18788 19388 18840 19440
rect 19984 19456 20036 19508
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 20444 19456 20496 19508
rect 6920 19320 6972 19372
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 6000 19252 6052 19304
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 5816 19184 5868 19236
rect 6276 19184 6328 19236
rect 11244 19320 11296 19372
rect 9036 19252 9088 19304
rect 9680 19252 9732 19304
rect 9864 19252 9916 19304
rect 10416 19252 10468 19304
rect 13084 19320 13136 19372
rect 18144 19320 18196 19372
rect 9956 19184 10008 19236
rect 10784 19184 10836 19236
rect 12440 19252 12492 19304
rect 13452 19252 13504 19304
rect 17132 19252 17184 19304
rect 17592 19295 17644 19304
rect 17592 19261 17601 19295
rect 17601 19261 17635 19295
rect 17635 19261 17644 19295
rect 17592 19252 17644 19261
rect 17868 19252 17920 19304
rect 5908 19116 5960 19168
rect 8300 19116 8352 19168
rect 8484 19116 8536 19168
rect 12532 19184 12584 19236
rect 11244 19116 11296 19168
rect 18144 19184 18196 19236
rect 18880 19295 18932 19304
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 18972 19252 19024 19304
rect 19616 19388 19668 19440
rect 20628 19456 20680 19508
rect 22192 19456 22244 19508
rect 20260 19320 20312 19372
rect 22468 19431 22520 19440
rect 22468 19397 22477 19431
rect 22477 19397 22511 19431
rect 22511 19397 22520 19431
rect 22468 19388 22520 19397
rect 23940 19456 23992 19508
rect 24032 19431 24084 19440
rect 20628 19320 20680 19372
rect 19616 19252 19668 19304
rect 20444 19252 20496 19304
rect 20536 19252 20588 19304
rect 21272 19252 21324 19304
rect 24032 19397 24041 19431
rect 24041 19397 24075 19431
rect 24075 19397 24084 19431
rect 24032 19388 24084 19397
rect 25596 19431 25648 19440
rect 19708 19184 19760 19236
rect 21640 19184 21692 19236
rect 12900 19116 12952 19168
rect 20444 19116 20496 19168
rect 20720 19116 20772 19168
rect 24676 19252 24728 19304
rect 25136 19252 25188 19304
rect 25320 19252 25372 19304
rect 24492 19184 24544 19236
rect 25596 19397 25605 19431
rect 25605 19397 25639 19431
rect 25639 19397 25648 19431
rect 25596 19388 25648 19397
rect 26424 19388 26476 19440
rect 26976 19388 27028 19440
rect 27344 19431 27396 19440
rect 27344 19397 27353 19431
rect 27353 19397 27387 19431
rect 27387 19397 27396 19431
rect 27344 19388 27396 19397
rect 27620 19388 27672 19440
rect 28816 19431 28868 19440
rect 28816 19397 28825 19431
rect 28825 19397 28859 19431
rect 28859 19397 28868 19431
rect 28816 19388 28868 19397
rect 29920 19456 29972 19508
rect 37924 19456 37976 19508
rect 29828 19431 29880 19440
rect 29828 19397 29837 19431
rect 29837 19397 29871 19431
rect 29871 19397 29880 19431
rect 29828 19388 29880 19397
rect 30196 19388 30248 19440
rect 30380 19431 30432 19440
rect 30380 19397 30389 19431
rect 30389 19397 30423 19431
rect 30423 19397 30432 19431
rect 30380 19388 30432 19397
rect 30564 19388 30616 19440
rect 31484 19363 31536 19372
rect 31484 19329 31493 19363
rect 31493 19329 31527 19363
rect 31527 19329 31536 19363
rect 31484 19320 31536 19329
rect 37832 19363 37884 19372
rect 37832 19329 37841 19363
rect 37841 19329 37875 19363
rect 37875 19329 37884 19363
rect 37832 19320 37884 19329
rect 25596 19252 25648 19304
rect 29460 19252 29512 19304
rect 30104 19252 30156 19304
rect 30656 19295 30708 19304
rect 30656 19261 30665 19295
rect 30665 19261 30699 19295
rect 30699 19261 30708 19295
rect 30656 19252 30708 19261
rect 26884 19184 26936 19236
rect 27068 19184 27120 19236
rect 28080 19184 28132 19236
rect 26792 19116 26844 19168
rect 28264 19116 28316 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2044 18912 2096 18964
rect 14924 18912 14976 18964
rect 15476 18912 15528 18964
rect 15844 18912 15896 18964
rect 16856 18912 16908 18964
rect 17868 18912 17920 18964
rect 8116 18844 8168 18896
rect 9864 18844 9916 18896
rect 11980 18844 12032 18896
rect 12256 18844 12308 18896
rect 1860 18776 1912 18828
rect 3976 18819 4028 18828
rect 3976 18785 3985 18819
rect 3985 18785 4019 18819
rect 4019 18785 4028 18819
rect 3976 18776 4028 18785
rect 4804 18776 4856 18828
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 11152 18776 11204 18828
rect 14096 18844 14148 18896
rect 12532 18776 12584 18828
rect 13452 18776 13504 18828
rect 13820 18776 13872 18828
rect 17224 18844 17276 18896
rect 17408 18844 17460 18896
rect 18972 18912 19024 18964
rect 18144 18844 18196 18896
rect 19984 18912 20036 18964
rect 26424 18912 26476 18964
rect 26884 18955 26936 18964
rect 26884 18921 26893 18955
rect 26893 18921 26927 18955
rect 26927 18921 26936 18955
rect 26884 18912 26936 18921
rect 27068 18912 27120 18964
rect 22008 18844 22060 18896
rect 24952 18844 25004 18896
rect 30012 18844 30064 18896
rect 5356 18708 5408 18760
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 2872 18640 2924 18692
rect 8760 18640 8812 18692
rect 9220 18751 9272 18760
rect 9220 18717 9229 18751
rect 9229 18717 9263 18751
rect 9263 18717 9272 18751
rect 9220 18708 9272 18717
rect 9680 18708 9732 18760
rect 10048 18640 10100 18692
rect 8484 18572 8536 18624
rect 11428 18572 11480 18624
rect 11888 18640 11940 18692
rect 13176 18640 13228 18692
rect 13820 18572 13872 18624
rect 14188 18640 14240 18692
rect 17960 18776 18012 18828
rect 15476 18708 15528 18760
rect 18236 18776 18288 18828
rect 19340 18776 19392 18828
rect 19616 18776 19668 18828
rect 20536 18819 20588 18828
rect 20536 18785 20545 18819
rect 20545 18785 20579 18819
rect 20579 18785 20588 18819
rect 20536 18776 20588 18785
rect 21272 18776 21324 18828
rect 22468 18776 22520 18828
rect 22928 18819 22980 18828
rect 22928 18785 22937 18819
rect 22937 18785 22971 18819
rect 22971 18785 22980 18819
rect 22928 18776 22980 18785
rect 15384 18683 15436 18692
rect 15384 18649 15393 18683
rect 15393 18649 15427 18683
rect 15427 18649 15436 18683
rect 15384 18640 15436 18649
rect 15568 18640 15620 18692
rect 15660 18572 15712 18624
rect 16856 18640 16908 18692
rect 17408 18640 17460 18692
rect 18972 18708 19024 18760
rect 17960 18572 18012 18624
rect 18052 18572 18104 18624
rect 19248 18640 19300 18692
rect 19708 18640 19760 18692
rect 19977 18683 20029 18692
rect 19977 18649 19986 18683
rect 19986 18649 20020 18683
rect 20020 18649 20029 18683
rect 19977 18640 20029 18649
rect 18972 18572 19024 18624
rect 19340 18572 19392 18624
rect 20720 18572 20772 18624
rect 20996 18572 21048 18624
rect 21272 18640 21324 18692
rect 23480 18708 23532 18760
rect 25504 18776 25556 18828
rect 25688 18819 25740 18828
rect 25688 18785 25697 18819
rect 25697 18785 25731 18819
rect 25731 18785 25740 18819
rect 25688 18776 25740 18785
rect 25964 18776 26016 18828
rect 26148 18751 26200 18760
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 26792 18751 26844 18760
rect 26792 18717 26801 18751
rect 26801 18717 26835 18751
rect 26835 18717 26844 18751
rect 26792 18708 26844 18717
rect 24676 18640 24728 18692
rect 25136 18683 25188 18692
rect 25136 18649 25145 18683
rect 25145 18649 25179 18683
rect 25179 18649 25188 18683
rect 25136 18640 25188 18649
rect 25964 18640 26016 18692
rect 29092 18776 29144 18828
rect 29920 18776 29972 18828
rect 30196 18844 30248 18896
rect 31392 18776 31444 18828
rect 28632 18751 28684 18760
rect 28632 18717 28641 18751
rect 28641 18717 28675 18751
rect 28675 18717 28684 18751
rect 28632 18708 28684 18717
rect 32680 18751 32732 18760
rect 32680 18717 32689 18751
rect 32689 18717 32723 18751
rect 32723 18717 32732 18751
rect 32680 18708 32732 18717
rect 38292 18751 38344 18760
rect 38292 18717 38301 18751
rect 38301 18717 38335 18751
rect 38335 18717 38344 18751
rect 38292 18708 38344 18717
rect 27804 18640 27856 18692
rect 24032 18572 24084 18624
rect 26332 18572 26384 18624
rect 29368 18640 29420 18692
rect 29920 18683 29972 18692
rect 29920 18649 29929 18683
rect 29929 18649 29963 18683
rect 29963 18649 29972 18683
rect 31300 18683 31352 18692
rect 29920 18640 29972 18649
rect 31300 18649 31309 18683
rect 31309 18649 31343 18683
rect 31343 18649 31352 18683
rect 31300 18640 31352 18649
rect 28724 18615 28776 18624
rect 28724 18581 28733 18615
rect 28733 18581 28767 18615
rect 28767 18581 28776 18615
rect 28724 18572 28776 18581
rect 28816 18572 28868 18624
rect 34520 18572 34572 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1860 18368 1912 18420
rect 2228 18343 2280 18352
rect 2228 18309 2237 18343
rect 2237 18309 2271 18343
rect 2271 18309 2280 18343
rect 2228 18300 2280 18309
rect 4160 18300 4212 18352
rect 12348 18368 12400 18420
rect 10140 18300 10192 18352
rect 6460 18232 6512 18284
rect 8208 18232 8260 18284
rect 12532 18300 12584 18352
rect 13268 18300 13320 18352
rect 18880 18368 18932 18420
rect 19432 18368 19484 18420
rect 20812 18368 20864 18420
rect 2320 18164 2372 18216
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 4252 18164 4304 18216
rect 6828 18207 6880 18216
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 7840 18164 7892 18216
rect 8576 18164 8628 18216
rect 9220 18164 9272 18216
rect 11612 18232 11664 18284
rect 5448 18096 5500 18148
rect 10876 18164 10928 18216
rect 11888 18164 11940 18216
rect 12716 18164 12768 18216
rect 12992 18164 13044 18216
rect 4620 18028 4672 18080
rect 5356 18028 5408 18080
rect 6092 18028 6144 18080
rect 6920 18028 6972 18080
rect 7104 18028 7156 18080
rect 12072 18096 12124 18148
rect 13452 18300 13504 18352
rect 16948 18343 17000 18352
rect 14188 18164 14240 18216
rect 14924 18164 14976 18216
rect 15476 18164 15528 18216
rect 9588 18071 9640 18080
rect 9588 18037 9612 18071
rect 9612 18037 9640 18071
rect 9588 18028 9640 18037
rect 11244 18028 11296 18080
rect 12440 18028 12492 18080
rect 16672 18232 16724 18284
rect 16488 18164 16540 18216
rect 16948 18309 16957 18343
rect 16957 18309 16991 18343
rect 16991 18309 17000 18343
rect 16948 18300 17000 18309
rect 17960 18300 18012 18352
rect 18512 18300 18564 18352
rect 19248 18300 19300 18352
rect 19616 18343 19668 18352
rect 19616 18309 19625 18343
rect 19625 18309 19659 18343
rect 19659 18309 19668 18343
rect 19616 18300 19668 18309
rect 20352 18300 20404 18352
rect 21456 18368 21508 18420
rect 18420 18232 18472 18284
rect 18696 18232 18748 18284
rect 17960 18207 18012 18216
rect 17960 18173 17969 18207
rect 17969 18173 18003 18207
rect 18003 18173 18012 18207
rect 17960 18164 18012 18173
rect 18972 18164 19024 18216
rect 20628 18232 20680 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 21456 18164 21508 18216
rect 21640 18164 21692 18216
rect 22100 18164 22152 18216
rect 22468 18300 22520 18352
rect 24032 18300 24084 18352
rect 24860 18343 24912 18352
rect 24860 18309 24869 18343
rect 24869 18309 24903 18343
rect 24903 18309 24912 18343
rect 24860 18300 24912 18309
rect 25320 18368 25372 18420
rect 25964 18343 26016 18352
rect 25964 18309 25973 18343
rect 25973 18309 26007 18343
rect 26007 18309 26016 18343
rect 25964 18300 26016 18309
rect 27528 18300 27580 18352
rect 25688 18232 25740 18284
rect 26700 18232 26752 18284
rect 29920 18368 29972 18420
rect 29736 18300 29788 18352
rect 30104 18275 30156 18284
rect 30104 18241 30113 18275
rect 30113 18241 30147 18275
rect 30147 18241 30156 18275
rect 30104 18232 30156 18241
rect 30564 18232 30616 18284
rect 30840 18232 30892 18284
rect 24032 18164 24084 18216
rect 16948 18096 17000 18148
rect 19156 18096 19208 18148
rect 16396 18028 16448 18080
rect 18236 18028 18288 18080
rect 18420 18028 18472 18080
rect 18880 18028 18932 18080
rect 19524 18028 19576 18080
rect 20444 18096 20496 18148
rect 20168 18028 20220 18080
rect 21088 18096 21140 18148
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 20812 18028 20864 18080
rect 23480 18096 23532 18148
rect 24492 18164 24544 18216
rect 26332 18207 26384 18216
rect 25044 18096 25096 18148
rect 26332 18173 26341 18207
rect 26341 18173 26375 18207
rect 26375 18173 26384 18207
rect 26332 18164 26384 18173
rect 29000 18164 29052 18216
rect 26516 18096 26568 18148
rect 27252 18139 27304 18148
rect 27252 18105 27261 18139
rect 27261 18105 27295 18139
rect 27295 18105 27304 18139
rect 27252 18096 27304 18105
rect 30012 18164 30064 18216
rect 29460 18096 29512 18148
rect 27620 18028 27672 18080
rect 28080 18028 28132 18080
rect 29184 18028 29236 18080
rect 30196 18071 30248 18080
rect 30196 18037 30205 18071
rect 30205 18037 30239 18071
rect 30239 18037 30248 18071
rect 30196 18028 30248 18037
rect 30380 18028 30432 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2320 17688 2372 17740
rect 4988 17688 5040 17740
rect 6368 17756 6420 17808
rect 8300 17824 8352 17876
rect 14832 17824 14884 17876
rect 8760 17756 8812 17808
rect 5540 17688 5592 17740
rect 6460 17731 6512 17740
rect 6460 17697 6469 17731
rect 6469 17697 6503 17731
rect 6503 17697 6512 17731
rect 6460 17688 6512 17697
rect 6828 17688 6880 17740
rect 5356 17620 5408 17672
rect 3700 17552 3752 17604
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 6736 17595 6788 17604
rect 6736 17561 6745 17595
rect 6745 17561 6779 17595
rect 6779 17561 6788 17595
rect 6736 17552 6788 17561
rect 8208 17552 8260 17604
rect 8576 17688 8628 17740
rect 9404 17756 9456 17808
rect 11888 17756 11940 17808
rect 12900 17756 12952 17808
rect 16580 17824 16632 17876
rect 16856 17824 16908 17876
rect 17960 17824 18012 17876
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 9956 17688 10008 17740
rect 14372 17688 14424 17740
rect 15752 17688 15804 17740
rect 18420 17756 18472 17808
rect 17040 17731 17092 17740
rect 17040 17697 17049 17731
rect 17049 17697 17083 17731
rect 17083 17697 17092 17731
rect 17040 17688 17092 17697
rect 18788 17688 18840 17740
rect 19616 17824 19668 17876
rect 19892 17824 19944 17876
rect 24124 17824 24176 17876
rect 24676 17824 24728 17876
rect 24860 17824 24912 17876
rect 25964 17824 26016 17876
rect 30748 17824 30800 17876
rect 18972 17756 19024 17808
rect 20444 17756 20496 17808
rect 21364 17799 21416 17808
rect 21364 17765 21373 17799
rect 21373 17765 21407 17799
rect 21407 17765 21416 17799
rect 21364 17756 21416 17765
rect 21916 17756 21968 17808
rect 29828 17756 29880 17808
rect 20812 17731 20864 17740
rect 9404 17620 9456 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 12532 17620 12584 17672
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 18420 17620 18472 17672
rect 9772 17552 9824 17604
rect 10508 17552 10560 17604
rect 12164 17552 12216 17604
rect 1032 17484 1084 17536
rect 2688 17484 2740 17536
rect 3884 17484 3936 17536
rect 4344 17484 4396 17536
rect 11796 17484 11848 17536
rect 12256 17484 12308 17536
rect 14188 17552 14240 17604
rect 14372 17595 14424 17604
rect 14372 17561 14381 17595
rect 14381 17561 14415 17595
rect 14415 17561 14424 17595
rect 14372 17552 14424 17561
rect 12532 17484 12584 17536
rect 14648 17552 14700 17604
rect 15568 17552 15620 17604
rect 14832 17484 14884 17536
rect 17776 17595 17828 17604
rect 17776 17561 17778 17595
rect 17778 17561 17812 17595
rect 17812 17561 17828 17595
rect 17776 17552 17828 17561
rect 17868 17552 17920 17604
rect 20812 17697 20821 17731
rect 20821 17697 20855 17731
rect 20855 17697 20864 17731
rect 20812 17688 20864 17697
rect 27252 17688 27304 17740
rect 27896 17688 27948 17740
rect 22284 17620 22336 17672
rect 22560 17663 22612 17672
rect 22560 17629 22569 17663
rect 22569 17629 22603 17663
rect 22603 17629 22612 17663
rect 22560 17620 22612 17629
rect 23112 17620 23164 17672
rect 23296 17620 23348 17672
rect 23848 17663 23900 17672
rect 23848 17629 23857 17663
rect 23857 17629 23891 17663
rect 23891 17629 23900 17663
rect 23848 17620 23900 17629
rect 19524 17595 19576 17604
rect 19524 17561 19533 17595
rect 19533 17561 19567 17595
rect 19567 17561 19576 17595
rect 19524 17552 19576 17561
rect 16580 17484 16632 17536
rect 17316 17484 17368 17536
rect 17960 17484 18012 17536
rect 19984 17484 20036 17536
rect 20812 17552 20864 17604
rect 21180 17552 21232 17604
rect 24492 17552 24544 17604
rect 24676 17595 24728 17604
rect 24676 17561 24685 17595
rect 24685 17561 24719 17595
rect 24719 17561 24728 17595
rect 24676 17552 24728 17561
rect 24768 17595 24820 17604
rect 24768 17561 24777 17595
rect 24777 17561 24811 17595
rect 24811 17561 24820 17595
rect 24768 17552 24820 17561
rect 25412 17552 25464 17604
rect 22100 17484 22152 17536
rect 23296 17527 23348 17536
rect 23296 17493 23305 17527
rect 23305 17493 23339 17527
rect 23339 17493 23348 17527
rect 23296 17484 23348 17493
rect 23940 17527 23992 17536
rect 23940 17493 23949 17527
rect 23949 17493 23983 17527
rect 23983 17493 23992 17527
rect 23940 17484 23992 17493
rect 24124 17484 24176 17536
rect 26792 17620 26844 17672
rect 27068 17620 27120 17672
rect 27252 17595 27304 17604
rect 27252 17561 27261 17595
rect 27261 17561 27295 17595
rect 27295 17561 27304 17595
rect 27252 17552 27304 17561
rect 30196 17688 30248 17740
rect 37372 17688 37424 17740
rect 31116 17663 31168 17672
rect 27436 17484 27488 17536
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 34520 17620 34572 17672
rect 29828 17595 29880 17604
rect 29828 17561 29837 17595
rect 29837 17561 29871 17595
rect 29871 17561 29880 17595
rect 29828 17552 29880 17561
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 30012 17552 30064 17604
rect 30472 17595 30524 17604
rect 30472 17561 30481 17595
rect 30481 17561 30515 17595
rect 30515 17561 30524 17595
rect 30472 17552 30524 17561
rect 28816 17484 28868 17493
rect 30380 17484 30432 17536
rect 30656 17484 30708 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 2688 17280 2740 17332
rect 572 17212 624 17264
rect 4344 17255 4396 17264
rect 4344 17221 4353 17255
rect 4353 17221 4387 17255
rect 4387 17221 4396 17255
rect 4344 17212 4396 17221
rect 4896 17255 4948 17264
rect 4896 17221 4905 17255
rect 4905 17221 4939 17255
rect 4939 17221 4948 17255
rect 4896 17212 4948 17221
rect 11428 17280 11480 17332
rect 11704 17280 11756 17332
rect 8760 17212 8812 17264
rect 2320 17187 2372 17196
rect 2320 17153 2329 17187
rect 2329 17153 2363 17187
rect 2363 17153 2372 17187
rect 2320 17144 2372 17153
rect 6460 17144 6512 17196
rect 9036 17212 9088 17264
rect 9128 17255 9180 17264
rect 9128 17221 9137 17255
rect 9137 17221 9171 17255
rect 9171 17221 9180 17255
rect 9128 17212 9180 17221
rect 9404 17212 9456 17264
rect 11980 17255 12032 17264
rect 11980 17221 11989 17255
rect 11989 17221 12023 17255
rect 12023 17221 12032 17255
rect 11980 17212 12032 17221
rect 10600 17144 10652 17196
rect 10968 17144 11020 17196
rect 5172 17119 5224 17128
rect 5172 17085 5181 17119
rect 5181 17085 5215 17119
rect 5215 17085 5224 17119
rect 5172 17076 5224 17085
rect 8576 17008 8628 17060
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 2412 16940 2464 16992
rect 4896 16940 4948 16992
rect 5080 16940 5132 16992
rect 8760 16940 8812 16992
rect 10140 16940 10192 16992
rect 10784 17076 10836 17128
rect 11428 17076 11480 17128
rect 13360 17076 13412 17128
rect 13728 17076 13780 17128
rect 16580 17280 16632 17332
rect 15384 17255 15436 17264
rect 15384 17221 15393 17255
rect 15393 17221 15427 17255
rect 15427 17221 15436 17255
rect 15384 17212 15436 17221
rect 17040 17255 17092 17264
rect 17040 17221 17049 17255
rect 17049 17221 17083 17255
rect 17083 17221 17092 17255
rect 17040 17212 17092 17221
rect 17592 17280 17644 17332
rect 18512 17280 18564 17332
rect 18604 17280 18656 17332
rect 23940 17280 23992 17332
rect 24032 17323 24084 17332
rect 24032 17289 24041 17323
rect 24041 17289 24075 17323
rect 24075 17289 24084 17323
rect 24032 17280 24084 17289
rect 25136 17280 25188 17332
rect 27436 17280 27488 17332
rect 27528 17280 27580 17332
rect 19064 17212 19116 17264
rect 20076 17212 20128 17264
rect 20904 17212 20956 17264
rect 22192 17255 22244 17264
rect 22192 17221 22201 17255
rect 22201 17221 22235 17255
rect 22235 17221 22244 17255
rect 22192 17212 22244 17221
rect 23112 17212 23164 17264
rect 24952 17212 25004 17264
rect 28540 17212 28592 17264
rect 16580 17076 16632 17128
rect 11980 16940 12032 16992
rect 12072 16940 12124 16992
rect 14372 16940 14424 16992
rect 15200 17008 15252 17060
rect 15476 17008 15528 17060
rect 17868 17076 17920 17128
rect 17960 17119 18012 17128
rect 17960 17085 17969 17119
rect 17969 17085 18003 17119
rect 18003 17085 18012 17119
rect 17960 17076 18012 17085
rect 18512 17076 18564 17128
rect 18880 17076 18932 17128
rect 20168 17144 20220 17196
rect 17132 17008 17184 17060
rect 17592 17008 17644 17060
rect 17776 17008 17828 17060
rect 21916 17144 21968 17196
rect 22836 17187 22888 17196
rect 22836 17153 22845 17187
rect 22845 17153 22879 17187
rect 22879 17153 22888 17187
rect 22836 17144 22888 17153
rect 23204 17144 23256 17196
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 30564 17280 30616 17332
rect 31576 17212 31628 17264
rect 22652 17076 22704 17128
rect 25136 17076 25188 17128
rect 26240 17076 26292 17128
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 27528 17119 27580 17128
rect 27528 17085 27537 17119
rect 27537 17085 27571 17119
rect 27571 17085 27580 17119
rect 27528 17076 27580 17085
rect 27712 17076 27764 17128
rect 31116 17144 31168 17196
rect 29000 17076 29052 17128
rect 30104 17076 30156 17128
rect 24032 16940 24084 16992
rect 28908 17008 28960 17060
rect 30748 17008 30800 17060
rect 37464 17119 37516 17128
rect 37464 17085 37473 17119
rect 37473 17085 37507 17119
rect 37507 17085 37516 17119
rect 37464 17076 37516 17085
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5816 16736 5868 16788
rect 6092 16736 6144 16788
rect 1584 16600 1636 16652
rect 2320 16600 2372 16652
rect 2688 16600 2740 16652
rect 4620 16600 4672 16652
rect 5356 16600 5408 16652
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7564 16600 7616 16652
rect 9864 16736 9916 16788
rect 8300 16668 8352 16720
rect 8760 16600 8812 16652
rect 9680 16600 9732 16652
rect 11980 16668 12032 16720
rect 16948 16736 17000 16788
rect 17040 16736 17092 16788
rect 22928 16736 22980 16788
rect 23112 16736 23164 16788
rect 23204 16736 23256 16788
rect 24032 16736 24084 16788
rect 27252 16736 27304 16788
rect 27436 16736 27488 16788
rect 28356 16736 28408 16788
rect 33508 16736 33560 16788
rect 15384 16668 15436 16720
rect 28816 16668 28868 16720
rect 29644 16668 29696 16720
rect 3424 16532 3476 16584
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 15568 16600 15620 16652
rect 16580 16600 16632 16652
rect 17500 16600 17552 16652
rect 17592 16600 17644 16652
rect 17776 16600 17828 16652
rect 1768 16396 1820 16448
rect 4068 16464 4120 16516
rect 4344 16464 4396 16516
rect 3240 16396 3292 16448
rect 6736 16464 6788 16516
rect 8208 16464 8260 16516
rect 8668 16464 8720 16516
rect 9036 16464 9088 16516
rect 9772 16464 9824 16516
rect 10140 16464 10192 16516
rect 10508 16464 10560 16516
rect 10784 16464 10836 16516
rect 10876 16507 10928 16516
rect 10876 16473 10885 16507
rect 10885 16473 10919 16507
rect 10919 16473 10928 16507
rect 10876 16464 10928 16473
rect 12164 16464 12216 16516
rect 12348 16532 12400 16584
rect 12440 16464 12492 16516
rect 12808 16464 12860 16516
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 13912 16532 13964 16584
rect 14096 16532 14148 16584
rect 14648 16532 14700 16584
rect 13636 16464 13688 16516
rect 15200 16507 15252 16516
rect 15200 16473 15209 16507
rect 15209 16473 15243 16507
rect 15243 16473 15252 16507
rect 15200 16464 15252 16473
rect 17316 16464 17368 16516
rect 19708 16600 19760 16652
rect 19800 16600 19852 16652
rect 20536 16600 20588 16652
rect 18604 16532 18656 16584
rect 20720 16643 20772 16652
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 22284 16600 22336 16652
rect 19064 16464 19116 16516
rect 4712 16396 4764 16448
rect 4988 16396 5040 16448
rect 6184 16396 6236 16448
rect 8852 16396 8904 16448
rect 14464 16396 14516 16448
rect 15016 16396 15068 16448
rect 16304 16396 16356 16448
rect 16488 16396 16540 16448
rect 18880 16396 18932 16448
rect 22744 16600 22796 16652
rect 22836 16532 22888 16584
rect 23388 16532 23440 16584
rect 23664 16532 23716 16584
rect 27896 16600 27948 16652
rect 19524 16507 19576 16516
rect 19524 16473 19533 16507
rect 19533 16473 19567 16507
rect 19567 16473 19576 16507
rect 19524 16464 19576 16473
rect 19984 16464 20036 16516
rect 20352 16464 20404 16516
rect 21088 16464 21140 16516
rect 24676 16507 24728 16516
rect 22100 16396 22152 16448
rect 24676 16473 24685 16507
rect 24685 16473 24719 16507
rect 24719 16473 24728 16507
rect 24676 16464 24728 16473
rect 27620 16532 27672 16584
rect 27712 16575 27764 16584
rect 27712 16541 27721 16575
rect 27721 16541 27755 16575
rect 27755 16541 27764 16575
rect 27712 16532 27764 16541
rect 28448 16575 28500 16584
rect 28448 16541 28457 16575
rect 28457 16541 28491 16575
rect 28491 16541 28500 16575
rect 28448 16532 28500 16541
rect 29092 16575 29144 16584
rect 29092 16541 29101 16575
rect 29101 16541 29135 16575
rect 29135 16541 29144 16575
rect 30840 16668 30892 16720
rect 30288 16600 30340 16652
rect 37188 16600 37240 16652
rect 29092 16532 29144 16541
rect 26056 16464 26108 16516
rect 26240 16507 26292 16516
rect 26240 16473 26249 16507
rect 26249 16473 26283 16507
rect 26283 16473 26292 16507
rect 26240 16464 26292 16473
rect 22836 16396 22888 16448
rect 25872 16396 25924 16448
rect 27068 16464 27120 16516
rect 38108 16507 38160 16516
rect 38108 16473 38117 16507
rect 38117 16473 38151 16507
rect 38151 16473 38160 16507
rect 38108 16464 38160 16473
rect 27804 16439 27856 16448
rect 27804 16405 27813 16439
rect 27813 16405 27847 16439
rect 27847 16405 27856 16439
rect 27804 16396 27856 16405
rect 28080 16396 28132 16448
rect 29736 16396 29788 16448
rect 30472 16439 30524 16448
rect 30472 16405 30481 16439
rect 30481 16405 30515 16439
rect 30515 16405 30524 16439
rect 30472 16396 30524 16405
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 5172 16192 5224 16244
rect 7104 16235 7156 16244
rect 7104 16201 7113 16235
rect 7113 16201 7147 16235
rect 7147 16201 7156 16235
rect 7104 16192 7156 16201
rect 4344 16124 4396 16176
rect 7656 16124 7708 16176
rect 10508 16192 10560 16244
rect 9588 16124 9640 16176
rect 10968 16167 11020 16176
rect 10968 16133 10977 16167
rect 10977 16133 11011 16167
rect 11011 16133 11020 16167
rect 10968 16124 11020 16133
rect 11060 16124 11112 16176
rect 11336 16124 11388 16176
rect 11980 16124 12032 16176
rect 12440 16124 12492 16176
rect 13544 16192 13596 16244
rect 16396 16192 16448 16244
rect 15016 16124 15068 16176
rect 15384 16167 15436 16176
rect 15384 16133 15393 16167
rect 15393 16133 15427 16167
rect 15427 16133 15436 16167
rect 15384 16124 15436 16133
rect 16764 16124 16816 16176
rect 27252 16235 27304 16244
rect 27252 16201 27261 16235
rect 27261 16201 27295 16235
rect 27295 16201 27304 16235
rect 27252 16192 27304 16201
rect 17408 16124 17460 16176
rect 18604 16124 18656 16176
rect 18788 16167 18840 16176
rect 18788 16133 18797 16167
rect 18797 16133 18831 16167
rect 18831 16133 18840 16167
rect 18788 16124 18840 16133
rect 19248 16124 19300 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2688 16099 2740 16108
rect 2688 16065 2697 16099
rect 2697 16065 2731 16099
rect 2731 16065 2740 16099
rect 2688 16056 2740 16065
rect 3700 15852 3752 15904
rect 4252 16056 4304 16108
rect 7012 16099 7064 16108
rect 7012 16065 7021 16099
rect 7021 16065 7055 16099
rect 7055 16065 7064 16099
rect 7012 16056 7064 16065
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 6552 15988 6604 16040
rect 8668 15988 8720 16040
rect 9496 16056 9548 16108
rect 10048 16056 10100 16108
rect 10140 16056 10192 16108
rect 19800 16124 19852 16176
rect 19984 16124 20036 16176
rect 20904 16124 20956 16176
rect 22100 16167 22152 16176
rect 22100 16133 22109 16167
rect 22109 16133 22143 16167
rect 22143 16133 22152 16167
rect 22100 16124 22152 16133
rect 23204 16124 23256 16176
rect 24308 16167 24360 16176
rect 24308 16133 24317 16167
rect 24317 16133 24351 16167
rect 24351 16133 24360 16167
rect 24308 16124 24360 16133
rect 24768 16124 24820 16176
rect 27804 16124 27856 16176
rect 11520 16056 11572 16108
rect 13912 16056 13964 16108
rect 19432 16056 19484 16108
rect 19616 16056 19668 16108
rect 20444 16056 20496 16108
rect 20720 16056 20772 16108
rect 11060 15988 11112 16040
rect 11336 15988 11388 16040
rect 13636 15988 13688 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 14372 16031 14424 16040
rect 13728 15988 13780 15997
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 16948 16031 17000 16040
rect 5264 15852 5316 15904
rect 6184 15852 6236 15904
rect 6644 15852 6696 15904
rect 10968 15920 11020 15972
rect 14004 15920 14056 15972
rect 14832 15920 14884 15972
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 17408 15988 17460 16040
rect 17868 15988 17920 16040
rect 17960 16031 18012 16040
rect 17960 15997 17969 16031
rect 17969 15997 18003 16031
rect 18003 15997 18012 16031
rect 17960 15988 18012 15997
rect 18880 15988 18932 16040
rect 17224 15920 17276 15972
rect 20904 15988 20956 16040
rect 21640 15988 21692 16040
rect 21916 15988 21968 16040
rect 22100 15988 22152 16040
rect 23388 16056 23440 16108
rect 24860 16099 24912 16108
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 23112 15988 23164 15997
rect 13176 15852 13228 15904
rect 13268 15852 13320 15904
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 21824 15920 21876 15972
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 25044 16056 25096 16108
rect 26148 16099 26200 16108
rect 26148 16065 26157 16099
rect 26157 16065 26191 16099
rect 26191 16065 26200 16099
rect 26148 16056 26200 16065
rect 27252 16056 27304 16108
rect 24676 15988 24728 16040
rect 31116 16192 31168 16244
rect 31576 16235 31628 16244
rect 31576 16201 31585 16235
rect 31585 16201 31619 16235
rect 31619 16201 31628 16235
rect 31576 16192 31628 16201
rect 38016 16192 38068 16244
rect 28264 16167 28316 16176
rect 28264 16133 28273 16167
rect 28273 16133 28307 16167
rect 28307 16133 28316 16167
rect 28264 16124 28316 16133
rect 29184 16167 29236 16176
rect 29184 16133 29193 16167
rect 29193 16133 29227 16167
rect 29227 16133 29236 16167
rect 29184 16124 29236 16133
rect 29552 16124 29604 16176
rect 30472 16124 30524 16176
rect 30840 16099 30892 16108
rect 30840 16065 30849 16099
rect 30849 16065 30883 16099
rect 30883 16065 30892 16099
rect 30840 16056 30892 16065
rect 31116 16056 31168 16108
rect 35900 16056 35952 16108
rect 29000 15988 29052 16040
rect 30012 16031 30064 16040
rect 30012 15997 30021 16031
rect 30021 15997 30055 16031
rect 30055 15997 30064 16031
rect 30012 15988 30064 15997
rect 24492 15920 24544 15972
rect 25872 15920 25924 15972
rect 28080 15920 28132 15972
rect 23664 15895 23716 15904
rect 23664 15861 23673 15895
rect 23673 15861 23707 15895
rect 23707 15861 23716 15895
rect 24952 15895 25004 15904
rect 23664 15852 23716 15861
rect 24952 15861 24961 15895
rect 24961 15861 24995 15895
rect 24995 15861 25004 15895
rect 24952 15852 25004 15861
rect 25136 15852 25188 15904
rect 29092 15920 29144 15972
rect 29184 15920 29236 15972
rect 28448 15852 28500 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 940 15648 992 15700
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 4252 15580 4304 15632
rect 1584 15512 1636 15521
rect 5724 15512 5776 15564
rect 6368 15512 6420 15564
rect 9220 15580 9272 15632
rect 11428 15648 11480 15700
rect 12348 15648 12400 15700
rect 13636 15648 13688 15700
rect 22100 15648 22152 15700
rect 22192 15648 22244 15700
rect 26148 15648 26200 15700
rect 26424 15648 26476 15700
rect 27160 15691 27212 15700
rect 27160 15657 27169 15691
rect 27169 15657 27203 15691
rect 27203 15657 27212 15691
rect 27160 15648 27212 15657
rect 27620 15648 27672 15700
rect 33508 15648 33560 15700
rect 13084 15580 13136 15632
rect 7288 15512 7340 15564
rect 7932 15512 7984 15564
rect 8668 15512 8720 15564
rect 9680 15512 9732 15564
rect 10048 15512 10100 15564
rect 5356 15487 5408 15496
rect 5356 15453 5365 15487
rect 5365 15453 5399 15487
rect 5399 15453 5408 15487
rect 5356 15444 5408 15453
rect 4068 15376 4120 15428
rect 4620 15376 4672 15428
rect 5908 15376 5960 15428
rect 7656 15376 7708 15428
rect 8116 15376 8168 15428
rect 8392 15376 8444 15428
rect 8760 15444 8812 15496
rect 8668 15376 8720 15428
rect 9496 15376 9548 15428
rect 3240 15308 3292 15360
rect 3700 15308 3752 15360
rect 6368 15308 6420 15360
rect 6644 15308 6696 15360
rect 9680 15308 9732 15360
rect 10048 15376 10100 15428
rect 11060 15512 11112 15564
rect 11336 15512 11388 15564
rect 11520 15555 11572 15564
rect 11520 15521 11529 15555
rect 11529 15521 11563 15555
rect 11563 15521 11572 15555
rect 11520 15512 11572 15521
rect 16304 15580 16356 15632
rect 16396 15580 16448 15632
rect 22744 15580 22796 15632
rect 24584 15580 24636 15632
rect 26976 15580 27028 15632
rect 27804 15580 27856 15632
rect 31392 15580 31444 15632
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17500 15512 17552 15564
rect 17224 15444 17276 15453
rect 17592 15444 17644 15496
rect 18972 15512 19024 15564
rect 20260 15444 20312 15496
rect 20536 15444 20588 15496
rect 20812 15444 20864 15496
rect 22284 15512 22336 15564
rect 22652 15444 22704 15496
rect 27528 15512 27580 15564
rect 28356 15555 28408 15564
rect 28356 15521 28365 15555
rect 28365 15521 28399 15555
rect 28399 15521 28408 15555
rect 28356 15512 28408 15521
rect 26332 15444 26384 15496
rect 26976 15444 27028 15496
rect 11796 15419 11848 15428
rect 11796 15385 11805 15419
rect 11805 15385 11839 15419
rect 11839 15385 11848 15419
rect 11796 15376 11848 15385
rect 11888 15376 11940 15428
rect 11152 15308 11204 15360
rect 14004 15376 14056 15428
rect 14648 15376 14700 15428
rect 16580 15419 16632 15428
rect 16580 15385 16589 15419
rect 16589 15385 16623 15419
rect 16623 15385 16632 15419
rect 16580 15376 16632 15385
rect 16396 15308 16448 15360
rect 20076 15376 20128 15428
rect 18880 15308 18932 15360
rect 19156 15308 19208 15360
rect 19892 15308 19944 15360
rect 21272 15308 21324 15360
rect 21456 15419 21508 15428
rect 21456 15385 21465 15419
rect 21465 15385 21499 15419
rect 21499 15385 21508 15419
rect 21456 15376 21508 15385
rect 22560 15376 22612 15428
rect 22928 15419 22980 15428
rect 22928 15385 22937 15419
rect 22937 15385 22971 15419
rect 22971 15385 22980 15419
rect 22928 15376 22980 15385
rect 23020 15419 23072 15428
rect 23020 15385 23029 15419
rect 23029 15385 23063 15419
rect 23063 15385 23072 15419
rect 23020 15376 23072 15385
rect 23204 15376 23256 15428
rect 25136 15376 25188 15428
rect 22008 15308 22060 15360
rect 22192 15308 22244 15360
rect 26240 15376 26292 15428
rect 26424 15308 26476 15360
rect 26608 15376 26660 15428
rect 29276 15444 29328 15496
rect 29828 15444 29880 15496
rect 37740 15512 37792 15564
rect 37372 15444 37424 15496
rect 28172 15376 28224 15428
rect 28448 15419 28500 15428
rect 28448 15385 28457 15419
rect 28457 15385 28491 15419
rect 28491 15385 28500 15419
rect 28448 15376 28500 15385
rect 28816 15376 28868 15428
rect 27988 15308 28040 15360
rect 30564 15308 30616 15360
rect 38200 15351 38252 15360
rect 38200 15317 38209 15351
rect 38209 15317 38243 15351
rect 38243 15317 38252 15351
rect 38200 15308 38252 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 5356 15104 5408 15156
rect 664 15036 716 15088
rect 2136 15036 2188 15088
rect 3700 15036 3752 15088
rect 5816 15036 5868 15088
rect 6368 15036 6420 15088
rect 6460 15036 6512 15088
rect 7840 15104 7892 15156
rect 1584 15011 1636 15020
rect 1584 14977 1593 15011
rect 1593 14977 1627 15011
rect 1627 14977 1636 15011
rect 1584 14968 1636 14977
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 9496 15036 9548 15088
rect 3700 14764 3752 14816
rect 5080 14900 5132 14952
rect 11060 15104 11112 15156
rect 15752 15104 15804 15156
rect 16396 15104 16448 15156
rect 17040 15104 17092 15156
rect 17684 15104 17736 15156
rect 11888 15036 11940 15088
rect 12072 15036 12124 15088
rect 12440 15036 12492 15088
rect 15108 15036 15160 15088
rect 17500 15036 17552 15088
rect 18144 15104 18196 15156
rect 19156 15104 19208 15156
rect 11520 14968 11572 15020
rect 13912 14968 13964 15020
rect 16672 14968 16724 15020
rect 17132 14968 17184 15020
rect 18972 15036 19024 15088
rect 19432 15036 19484 15088
rect 19616 15036 19668 15088
rect 20536 15036 20588 15088
rect 20812 15079 20864 15088
rect 20812 15045 20821 15079
rect 20821 15045 20855 15079
rect 20855 15045 20864 15079
rect 20812 15036 20864 15045
rect 20904 15036 20956 15088
rect 21916 15036 21968 15088
rect 22192 15079 22244 15088
rect 22192 15045 22201 15079
rect 22201 15045 22235 15079
rect 22235 15045 22244 15079
rect 22192 15036 22244 15045
rect 23112 15079 23164 15088
rect 23112 15045 23121 15079
rect 23121 15045 23155 15079
rect 23155 15045 23164 15079
rect 23112 15036 23164 15045
rect 23296 15036 23348 15088
rect 24952 15036 25004 15088
rect 26608 15104 26660 15156
rect 27528 15104 27580 15156
rect 9864 14900 9916 14952
rect 6920 14832 6972 14884
rect 5724 14764 5776 14816
rect 6184 14764 6236 14816
rect 9956 14764 10008 14816
rect 10600 14900 10652 14952
rect 13452 14900 13504 14952
rect 13544 14900 13596 14952
rect 15384 14900 15436 14952
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 16304 14900 16356 14952
rect 17316 14900 17368 14952
rect 17868 14900 17920 14952
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 19064 14968 19116 15020
rect 19156 14968 19208 15020
rect 20076 14968 20128 15020
rect 10508 14832 10560 14884
rect 11152 14832 11204 14884
rect 11612 14832 11664 14884
rect 15108 14832 15160 14884
rect 18788 14900 18840 14952
rect 19248 14900 19300 14952
rect 18328 14832 18380 14884
rect 18696 14832 18748 14884
rect 19708 14832 19760 14884
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 20352 14900 20404 14952
rect 21640 14968 21692 15020
rect 25504 15036 25556 15088
rect 28356 15036 28408 15088
rect 28724 15079 28776 15088
rect 28724 15045 28733 15079
rect 28733 15045 28767 15079
rect 28767 15045 28776 15079
rect 28724 15036 28776 15045
rect 25320 14968 25372 15020
rect 26240 14968 26292 15020
rect 27344 14968 27396 15020
rect 20536 14832 20588 14884
rect 21824 14900 21876 14952
rect 22376 14900 22428 14952
rect 24308 14900 24360 14952
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 26148 14900 26200 14952
rect 26608 14900 26660 14952
rect 27712 14900 27764 14952
rect 29184 14943 29236 14952
rect 29184 14909 29193 14943
rect 29193 14909 29227 14943
rect 29227 14909 29236 14943
rect 29184 14900 29236 14909
rect 27344 14832 27396 14884
rect 30380 14968 30432 15020
rect 31116 15011 31168 15020
rect 31116 14977 31125 15011
rect 31125 14977 31159 15011
rect 31159 14977 31168 15011
rect 31116 14968 31168 14977
rect 37740 14968 37792 15020
rect 18972 14764 19024 14816
rect 23388 14764 23440 14816
rect 23572 14764 23624 14816
rect 24492 14764 24544 14816
rect 25688 14764 25740 14816
rect 26884 14764 26936 14816
rect 27068 14764 27120 14816
rect 29828 14764 29880 14816
rect 31208 14807 31260 14816
rect 31208 14773 31217 14807
rect 31217 14773 31251 14807
rect 31251 14773 31260 14807
rect 31208 14764 31260 14773
rect 38016 14764 38068 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 7564 14560 7616 14612
rect 10784 14560 10836 14612
rect 11428 14560 11480 14612
rect 11612 14560 11664 14612
rect 15108 14560 15160 14612
rect 15200 14560 15252 14612
rect 18696 14560 18748 14612
rect 18788 14560 18840 14612
rect 21548 14560 21600 14612
rect 22100 14603 22152 14612
rect 22100 14569 22109 14603
rect 22109 14569 22143 14603
rect 22143 14569 22152 14603
rect 22100 14560 22152 14569
rect 23296 14560 23348 14612
rect 26424 14560 26476 14612
rect 27712 14603 27764 14612
rect 27712 14569 27721 14603
rect 27721 14569 27755 14603
rect 27755 14569 27764 14603
rect 27712 14560 27764 14569
rect 37372 14603 37424 14612
rect 37372 14569 37381 14603
rect 37381 14569 37415 14603
rect 37415 14569 37424 14603
rect 37372 14560 37424 14569
rect 5356 14492 5408 14544
rect 7932 14492 7984 14544
rect 10508 14492 10560 14544
rect 1584 14424 1636 14476
rect 3148 14424 3200 14476
rect 6000 14467 6052 14476
rect 6000 14433 6009 14467
rect 6009 14433 6043 14467
rect 6043 14433 6052 14467
rect 6000 14424 6052 14433
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 7380 14424 7432 14476
rect 9956 14424 10008 14476
rect 10600 14424 10652 14476
rect 11520 14424 11572 14476
rect 14004 14492 14056 14544
rect 14280 14492 14332 14544
rect 17408 14492 17460 14544
rect 17500 14492 17552 14544
rect 12992 14424 13044 14476
rect 15108 14424 15160 14476
rect 15384 14424 15436 14476
rect 16396 14424 16448 14476
rect 16580 14424 16632 14476
rect 16764 14424 16816 14476
rect 17592 14424 17644 14476
rect 17960 14492 18012 14544
rect 18052 14492 18104 14544
rect 19892 14492 19944 14544
rect 19984 14492 20036 14544
rect 20444 14492 20496 14544
rect 5356 14356 5408 14408
rect 3884 14288 3936 14340
rect 6828 14331 6880 14340
rect 2780 14220 2832 14272
rect 6828 14297 6837 14331
rect 6837 14297 6871 14331
rect 6871 14297 6880 14331
rect 6828 14288 6880 14297
rect 8116 14288 8168 14340
rect 5540 14220 5592 14272
rect 6092 14220 6144 14272
rect 8760 14356 8812 14408
rect 12808 14356 12860 14408
rect 13912 14356 13964 14408
rect 9588 14331 9640 14340
rect 9588 14297 9597 14331
rect 9597 14297 9631 14331
rect 9631 14297 9640 14331
rect 9588 14288 9640 14297
rect 11244 14288 11296 14340
rect 13636 14288 13688 14340
rect 10324 14220 10376 14272
rect 10508 14220 10560 14272
rect 17224 14356 17276 14408
rect 14280 14331 14332 14340
rect 14280 14297 14289 14331
rect 14289 14297 14323 14331
rect 14323 14297 14332 14331
rect 14280 14288 14332 14297
rect 14464 14288 14516 14340
rect 14372 14220 14424 14272
rect 15660 14220 15712 14272
rect 16856 14220 16908 14272
rect 17040 14288 17092 14340
rect 17684 14331 17736 14340
rect 17684 14297 17693 14331
rect 17693 14297 17727 14331
rect 17727 14297 17736 14331
rect 17684 14288 17736 14297
rect 17500 14220 17552 14272
rect 17776 14220 17828 14272
rect 19340 14220 19392 14272
rect 20260 14220 20312 14272
rect 20536 14467 20588 14476
rect 20536 14433 20545 14467
rect 20545 14433 20579 14467
rect 20579 14433 20588 14467
rect 20536 14424 20588 14433
rect 21640 14356 21692 14408
rect 22100 14356 22152 14408
rect 27620 14492 27672 14544
rect 22652 14424 22704 14476
rect 24032 14424 24084 14476
rect 22744 14356 22796 14408
rect 23664 14399 23716 14408
rect 21548 14331 21600 14340
rect 21548 14297 21557 14331
rect 21557 14297 21591 14331
rect 21591 14297 21600 14331
rect 21548 14288 21600 14297
rect 22284 14288 22336 14340
rect 22376 14288 22428 14340
rect 23664 14365 23673 14399
rect 23673 14365 23707 14399
rect 23707 14365 23716 14399
rect 23664 14356 23716 14365
rect 21088 14220 21140 14272
rect 21180 14220 21232 14272
rect 21824 14220 21876 14272
rect 22744 14220 22796 14272
rect 22836 14220 22888 14272
rect 23296 14220 23348 14272
rect 24584 14220 24636 14272
rect 24860 14288 24912 14340
rect 25412 14356 25464 14408
rect 25688 14424 25740 14476
rect 29552 14424 29604 14476
rect 30288 14424 30340 14476
rect 31392 14467 31444 14476
rect 31392 14433 31401 14467
rect 31401 14433 31435 14467
rect 31435 14433 31444 14467
rect 31392 14424 31444 14433
rect 25872 14331 25924 14340
rect 25872 14297 25881 14331
rect 25881 14297 25915 14331
rect 25915 14297 25924 14331
rect 25872 14288 25924 14297
rect 26516 14331 26568 14340
rect 25688 14220 25740 14272
rect 26516 14297 26525 14331
rect 26525 14297 26559 14331
rect 26559 14297 26568 14331
rect 26516 14288 26568 14297
rect 26608 14288 26660 14340
rect 27160 14356 27212 14408
rect 27620 14401 27672 14408
rect 27620 14367 27629 14401
rect 27629 14367 27663 14401
rect 27663 14367 27672 14401
rect 27620 14356 27672 14367
rect 27712 14220 27764 14272
rect 27896 14220 27948 14272
rect 28448 14356 28500 14408
rect 29920 14356 29972 14408
rect 37188 14356 37240 14408
rect 37924 14356 37976 14408
rect 28172 14288 28224 14340
rect 28356 14220 28408 14272
rect 28908 14220 28960 14272
rect 31116 14288 31168 14340
rect 31208 14331 31260 14340
rect 31208 14297 31217 14331
rect 31217 14297 31251 14331
rect 31251 14297 31260 14331
rect 31208 14288 31260 14297
rect 29736 14263 29788 14272
rect 29736 14229 29745 14263
rect 29745 14229 29779 14263
rect 29779 14229 29788 14263
rect 29736 14220 29788 14229
rect 30472 14263 30524 14272
rect 30472 14229 30481 14263
rect 30481 14229 30515 14263
rect 30515 14229 30524 14263
rect 30472 14220 30524 14229
rect 38200 14263 38252 14272
rect 38200 14229 38209 14263
rect 38209 14229 38243 14263
rect 38243 14229 38252 14263
rect 38200 14220 38252 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4528 13991 4580 14000
rect 4528 13957 4537 13991
rect 4537 13957 4571 13991
rect 4571 13957 4580 13991
rect 4528 13948 4580 13957
rect 9864 14016 9916 14068
rect 1860 13880 1912 13932
rect 3884 13880 3936 13932
rect 6092 13880 6144 13932
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 4068 13812 4120 13864
rect 4712 13812 4764 13864
rect 7932 13948 7984 14000
rect 10508 13948 10560 14000
rect 10600 13991 10652 14000
rect 10600 13957 10609 13991
rect 10609 13957 10643 13991
rect 10643 13957 10652 13991
rect 10600 13948 10652 13957
rect 11980 13991 12032 14000
rect 11980 13957 11989 13991
rect 11989 13957 12023 13991
rect 12023 13957 12032 13991
rect 11980 13948 12032 13957
rect 6276 13880 6328 13932
rect 8392 13812 8444 13864
rect 9312 13812 9364 13864
rect 10048 13812 10100 13864
rect 11704 13855 11756 13864
rect 6552 13744 6604 13796
rect 10324 13744 10376 13796
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 15016 13948 15068 14000
rect 16304 13948 16356 14000
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 3792 13676 3844 13728
rect 6920 13676 6972 13728
rect 11612 13676 11664 13728
rect 11796 13676 11848 13728
rect 13360 13812 13412 13864
rect 14648 13812 14700 13864
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 16948 13991 17000 14000
rect 16948 13957 16957 13991
rect 16957 13957 16991 13991
rect 16991 13957 17000 13991
rect 16948 13948 17000 13957
rect 20076 14016 20128 14068
rect 21180 14059 21232 14068
rect 21180 14025 21189 14059
rect 21189 14025 21223 14059
rect 21223 14025 21232 14059
rect 21180 14016 21232 14025
rect 22284 14016 22336 14068
rect 22560 14016 22612 14068
rect 23296 14016 23348 14068
rect 17868 13948 17920 14000
rect 18328 13948 18380 14000
rect 18512 13948 18564 14000
rect 19064 13948 19116 14000
rect 19156 13948 19208 14000
rect 19892 13948 19944 14000
rect 20628 13948 20680 14000
rect 21548 13948 21600 14000
rect 21916 13948 21968 14000
rect 22192 13991 22244 14000
rect 22192 13957 22201 13991
rect 22201 13957 22235 13991
rect 22235 13957 22244 13991
rect 22192 13948 22244 13957
rect 26608 14016 26660 14068
rect 18052 13923 18104 13932
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 18144 13923 18196 13932
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13880 18196 13889
rect 18420 13880 18472 13932
rect 20444 13880 20496 13932
rect 20996 13880 21048 13932
rect 21824 13880 21876 13932
rect 22744 13880 22796 13932
rect 23112 13880 23164 13932
rect 17316 13812 17368 13864
rect 17592 13812 17644 13864
rect 19156 13812 19208 13864
rect 20904 13812 20956 13864
rect 22100 13855 22152 13864
rect 22100 13821 22109 13855
rect 22109 13821 22143 13855
rect 22143 13821 22152 13855
rect 22100 13812 22152 13821
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 16212 13744 16264 13796
rect 18052 13744 18104 13796
rect 18420 13744 18472 13796
rect 19432 13744 19484 13796
rect 19524 13744 19576 13796
rect 17776 13676 17828 13728
rect 17868 13676 17920 13728
rect 18328 13676 18380 13728
rect 18512 13676 18564 13728
rect 21916 13676 21968 13728
rect 24584 13880 24636 13932
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 27712 13880 27764 13932
rect 28908 14016 28960 14068
rect 29736 14016 29788 14068
rect 30288 14016 30340 14068
rect 37188 14016 37240 14068
rect 30472 13948 30524 14000
rect 37740 13880 37792 13932
rect 38292 13923 38344 13932
rect 38292 13889 38301 13923
rect 38301 13889 38335 13923
rect 38335 13889 38344 13923
rect 38292 13880 38344 13889
rect 24308 13812 24360 13864
rect 25412 13812 25464 13864
rect 25872 13855 25924 13864
rect 25872 13821 25881 13855
rect 25881 13821 25915 13855
rect 25915 13821 25924 13855
rect 25872 13812 25924 13821
rect 27068 13812 27120 13864
rect 29368 13855 29420 13864
rect 29368 13821 29377 13855
rect 29377 13821 29411 13855
rect 29411 13821 29420 13855
rect 29368 13812 29420 13821
rect 23112 13744 23164 13796
rect 24860 13744 24912 13796
rect 23940 13676 23992 13728
rect 30564 13744 30616 13796
rect 27252 13719 27304 13728
rect 27252 13685 27261 13719
rect 27261 13685 27295 13719
rect 27295 13685 27304 13719
rect 27252 13676 27304 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4804 13472 4856 13524
rect 5816 13472 5868 13524
rect 11152 13472 11204 13524
rect 10600 13404 10652 13456
rect 20812 13472 20864 13524
rect 20904 13472 20956 13524
rect 21456 13472 21508 13524
rect 23388 13472 23440 13524
rect 13268 13404 13320 13456
rect 20536 13404 20588 13456
rect 23664 13404 23716 13456
rect 29368 13472 29420 13524
rect 26516 13404 26568 13456
rect 2044 13336 2096 13388
rect 2504 13336 2556 13388
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 11428 13336 11480 13388
rect 12624 13336 12676 13388
rect 13176 13336 13228 13388
rect 13636 13336 13688 13388
rect 13820 13336 13872 13388
rect 15568 13336 15620 13388
rect 8944 13268 8996 13320
rect 9128 13268 9180 13320
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 16396 13336 16448 13388
rect 16672 13379 16724 13388
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 16764 13336 16816 13388
rect 17224 13336 17276 13388
rect 16948 13268 17000 13320
rect 19156 13336 19208 13388
rect 19248 13336 19300 13388
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 20260 13268 20312 13320
rect 4436 13200 4488 13252
rect 5816 13200 5868 13252
rect 6092 13243 6144 13252
rect 6092 13209 6101 13243
rect 6101 13209 6135 13243
rect 6135 13209 6144 13243
rect 6092 13200 6144 13209
rect 6736 13200 6788 13252
rect 6828 13243 6880 13252
rect 6828 13209 6837 13243
rect 6837 13209 6871 13243
rect 6871 13209 6880 13243
rect 6828 13200 6880 13209
rect 7104 13200 7156 13252
rect 8392 13200 8444 13252
rect 9036 13200 9088 13252
rect 10876 13200 10928 13252
rect 12072 13200 12124 13252
rect 12992 13200 13044 13252
rect 2964 13132 3016 13184
rect 3516 13132 3568 13184
rect 4988 13132 5040 13184
rect 14280 13132 14332 13184
rect 14464 13243 14516 13252
rect 14464 13209 14473 13243
rect 14473 13209 14507 13243
rect 14507 13209 14516 13243
rect 14464 13200 14516 13209
rect 15660 13200 15712 13252
rect 16396 13243 16448 13252
rect 16396 13209 16405 13243
rect 16405 13209 16439 13243
rect 16439 13209 16448 13243
rect 16396 13200 16448 13209
rect 16028 13132 16080 13184
rect 16304 13132 16356 13184
rect 16672 13200 16724 13252
rect 17960 13200 18012 13252
rect 18236 13243 18288 13252
rect 18236 13209 18245 13243
rect 18245 13209 18279 13243
rect 18279 13209 18288 13243
rect 18236 13200 18288 13209
rect 18604 13200 18656 13252
rect 18696 13200 18748 13252
rect 18972 13200 19024 13252
rect 19064 13200 19116 13252
rect 19340 13200 19392 13252
rect 19524 13243 19576 13252
rect 19524 13209 19533 13243
rect 19533 13209 19567 13243
rect 19567 13209 19576 13243
rect 19524 13200 19576 13209
rect 16580 13132 16632 13184
rect 19892 13200 19944 13252
rect 20996 13336 21048 13388
rect 21640 13379 21692 13388
rect 21640 13345 21649 13379
rect 21649 13345 21683 13379
rect 21683 13345 21692 13379
rect 21640 13336 21692 13345
rect 22100 13336 22152 13388
rect 22284 13336 22336 13388
rect 23572 13336 23624 13388
rect 20812 13268 20864 13320
rect 22744 13268 22796 13320
rect 20536 13200 20588 13252
rect 20904 13132 20956 13184
rect 22560 13200 22612 13252
rect 23296 13200 23348 13252
rect 22468 13132 22520 13184
rect 23848 13268 23900 13320
rect 24676 13243 24728 13252
rect 24676 13209 24685 13243
rect 24685 13209 24719 13243
rect 24719 13209 24728 13243
rect 24676 13200 24728 13209
rect 25688 13200 25740 13252
rect 25504 13132 25556 13184
rect 28172 13311 28224 13320
rect 28172 13277 28181 13311
rect 28181 13277 28215 13311
rect 28215 13277 28224 13311
rect 28172 13268 28224 13277
rect 28448 13268 28500 13320
rect 28632 13268 28684 13320
rect 29736 13311 29788 13320
rect 29736 13277 29745 13311
rect 29745 13277 29779 13311
rect 29779 13277 29788 13311
rect 29736 13268 29788 13277
rect 29920 13268 29972 13320
rect 27068 13243 27120 13252
rect 27068 13209 27077 13243
rect 27077 13209 27111 13243
rect 27111 13209 27120 13243
rect 27068 13200 27120 13209
rect 28908 13175 28960 13184
rect 28908 13141 28917 13175
rect 28917 13141 28951 13175
rect 28951 13141 28960 13175
rect 28908 13132 28960 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 4436 12928 4488 12980
rect 8484 12928 8536 12980
rect 940 12860 992 12912
rect 4160 12903 4212 12912
rect 4160 12869 4169 12903
rect 4169 12869 4203 12903
rect 4203 12869 4212 12903
rect 4160 12860 4212 12869
rect 6920 12903 6972 12912
rect 6920 12869 6929 12903
rect 6929 12869 6963 12903
rect 6963 12869 6972 12903
rect 6920 12860 6972 12869
rect 8208 12860 8260 12912
rect 2044 12792 2096 12844
rect 4528 12792 4580 12844
rect 3608 12724 3660 12776
rect 5540 12724 5592 12776
rect 6000 12792 6052 12844
rect 8944 12792 8996 12844
rect 11244 12928 11296 12980
rect 11888 12928 11940 12980
rect 9496 12860 9548 12912
rect 10784 12860 10836 12912
rect 13452 12860 13504 12912
rect 13728 12860 13780 12912
rect 14096 12860 14148 12912
rect 15752 12860 15804 12912
rect 16396 12928 16448 12980
rect 22284 12928 22336 12980
rect 22560 12928 22612 12980
rect 16764 12860 16816 12912
rect 17040 12903 17092 12912
rect 17040 12869 17049 12903
rect 17049 12869 17083 12903
rect 17083 12869 17092 12903
rect 17040 12860 17092 12869
rect 17868 12860 17920 12912
rect 13176 12792 13228 12844
rect 13360 12792 13412 12844
rect 15844 12835 15896 12844
rect 5816 12724 5868 12776
rect 6552 12724 6604 12776
rect 4068 12656 4120 12708
rect 10600 12724 10652 12776
rect 10968 12724 11020 12776
rect 11244 12724 11296 12776
rect 11704 12724 11756 12776
rect 13636 12724 13688 12776
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 14648 12724 14700 12776
rect 16304 12792 16356 12844
rect 18236 12860 18288 12912
rect 16120 12767 16172 12776
rect 16120 12733 16129 12767
rect 16129 12733 16163 12767
rect 16163 12733 16172 12767
rect 16120 12724 16172 12733
rect 17040 12724 17092 12776
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 17868 12724 17920 12776
rect 8484 12656 8536 12708
rect 9036 12656 9088 12708
rect 13084 12656 13136 12708
rect 13728 12656 13780 12708
rect 16488 12656 16540 12708
rect 19064 12767 19116 12776
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 19156 12724 19208 12776
rect 19708 12724 19760 12776
rect 18420 12656 18472 12708
rect 11888 12588 11940 12640
rect 12440 12588 12492 12640
rect 16212 12588 16264 12640
rect 17040 12588 17092 12640
rect 18144 12588 18196 12640
rect 18328 12588 18380 12640
rect 18604 12588 18656 12640
rect 18788 12588 18840 12640
rect 18972 12656 19024 12708
rect 19800 12656 19852 12708
rect 20536 12860 20588 12912
rect 20628 12860 20680 12912
rect 21456 12860 21508 12912
rect 21916 12860 21968 12912
rect 22744 12860 22796 12912
rect 23020 12928 23072 12980
rect 24032 12928 24084 12980
rect 24584 12928 24636 12980
rect 21732 12792 21784 12844
rect 23020 12792 23072 12844
rect 21180 12724 21232 12776
rect 22376 12724 22428 12776
rect 22928 12724 22980 12776
rect 23480 12792 23532 12844
rect 24768 12792 24820 12844
rect 24860 12792 24912 12844
rect 25228 12792 25280 12844
rect 27528 12792 27580 12844
rect 25964 12767 26016 12776
rect 20720 12656 20772 12708
rect 20812 12656 20864 12708
rect 21640 12656 21692 12708
rect 22284 12656 22336 12708
rect 25688 12656 25740 12708
rect 25964 12733 25973 12767
rect 25973 12733 26007 12767
rect 26007 12733 26016 12767
rect 25964 12724 26016 12733
rect 29184 12928 29236 12980
rect 30380 12928 30432 12980
rect 27988 12903 28040 12912
rect 27988 12869 27997 12903
rect 27997 12869 28031 12903
rect 28031 12869 28040 12903
rect 27988 12860 28040 12869
rect 30840 12903 30892 12912
rect 30840 12869 30849 12903
rect 30849 12869 30883 12903
rect 30883 12869 30892 12903
rect 30840 12860 30892 12869
rect 33968 12792 34020 12844
rect 36452 12792 36504 12844
rect 26240 12656 26292 12708
rect 28080 12724 28132 12776
rect 30748 12767 30800 12776
rect 30748 12733 30757 12767
rect 30757 12733 30791 12767
rect 30791 12733 30800 12767
rect 30748 12724 30800 12733
rect 31668 12767 31720 12776
rect 31668 12733 31677 12767
rect 31677 12733 31711 12767
rect 31711 12733 31720 12767
rect 31668 12724 31720 12733
rect 31024 12656 31076 12708
rect 26148 12588 26200 12640
rect 27068 12588 27120 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3884 12384 3936 12436
rect 4068 12384 4120 12436
rect 5724 12384 5776 12436
rect 8300 12384 8352 12436
rect 8484 12384 8536 12436
rect 7840 12316 7892 12368
rect 9036 12316 9088 12368
rect 10784 12316 10836 12368
rect 12900 12316 12952 12368
rect 13084 12316 13136 12368
rect 13912 12316 13964 12368
rect 1584 12248 1636 12300
rect 2044 12248 2096 12300
rect 5172 12248 5224 12300
rect 5632 12180 5684 12232
rect 3608 12112 3660 12164
rect 4160 12155 4212 12164
rect 4160 12121 4169 12155
rect 4169 12121 4203 12155
rect 4203 12121 4212 12155
rect 4160 12112 4212 12121
rect 4712 12112 4764 12164
rect 4896 12112 4948 12164
rect 1860 12044 1912 12096
rect 2872 12044 2924 12096
rect 6736 12248 6788 12300
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 13820 12248 13872 12300
rect 23480 12384 23532 12436
rect 26148 12384 26200 12436
rect 36452 12384 36504 12436
rect 14556 12316 14608 12368
rect 14740 12316 14792 12368
rect 15476 12316 15528 12368
rect 17684 12316 17736 12368
rect 17868 12316 17920 12368
rect 15292 12248 15344 12300
rect 8300 12180 8352 12232
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 9220 12180 9272 12232
rect 9588 12180 9640 12232
rect 10232 12180 10284 12232
rect 16580 12248 16632 12300
rect 17040 12248 17092 12300
rect 20904 12316 20956 12368
rect 21180 12316 21232 12368
rect 18052 12248 18104 12300
rect 5816 12044 5868 12096
rect 8116 12112 8168 12164
rect 8392 12155 8444 12164
rect 8392 12121 8401 12155
rect 8401 12121 8435 12155
rect 8435 12121 8444 12155
rect 8392 12112 8444 12121
rect 9680 12112 9732 12164
rect 10140 12112 10192 12164
rect 13360 12112 13412 12164
rect 14280 12155 14332 12164
rect 14280 12121 14289 12155
rect 14289 12121 14323 12155
rect 14323 12121 14332 12155
rect 14280 12112 14332 12121
rect 15016 12155 15068 12164
rect 15016 12121 15025 12155
rect 15025 12121 15059 12155
rect 15059 12121 15068 12155
rect 15016 12112 15068 12121
rect 16396 12180 16448 12232
rect 17868 12180 17920 12232
rect 7288 12044 7340 12096
rect 10232 12044 10284 12096
rect 10784 12044 10836 12096
rect 17316 12112 17368 12164
rect 17684 12112 17736 12164
rect 18512 12112 18564 12164
rect 22284 12248 22336 12300
rect 27988 12316 28040 12368
rect 37280 12316 37332 12368
rect 21364 12180 21416 12232
rect 18788 12112 18840 12164
rect 20904 12112 20956 12164
rect 22008 12112 22060 12164
rect 23020 12112 23072 12164
rect 23204 12155 23256 12164
rect 23204 12121 23213 12155
rect 23213 12121 23247 12155
rect 23247 12121 23256 12155
rect 23204 12112 23256 12121
rect 23848 12248 23900 12300
rect 24952 12248 25004 12300
rect 26056 12248 26108 12300
rect 24308 12180 24360 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 24676 12180 24728 12232
rect 27344 12223 27396 12232
rect 25136 12112 25188 12164
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 30748 12248 30800 12300
rect 31668 12180 31720 12232
rect 34060 12180 34112 12232
rect 26424 12112 26476 12164
rect 26976 12112 27028 12164
rect 21916 12044 21968 12096
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 23940 12044 23992 12096
rect 27160 12044 27212 12096
rect 27712 12044 27764 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 756 11840 808 11892
rect 2412 11772 2464 11824
rect 3240 11840 3292 11892
rect 3516 11840 3568 11892
rect 3792 11840 3844 11892
rect 3884 11840 3936 11892
rect 5172 11840 5224 11892
rect 4160 11772 4212 11824
rect 6828 11840 6880 11892
rect 8668 11840 8720 11892
rect 9312 11840 9364 11892
rect 9036 11772 9088 11824
rect 11520 11772 11572 11824
rect 13452 11772 13504 11824
rect 14556 11815 14608 11824
rect 14556 11781 14565 11815
rect 14565 11781 14599 11815
rect 14599 11781 14608 11815
rect 14556 11772 14608 11781
rect 15384 11772 15436 11824
rect 1584 11747 1636 11756
rect 1584 11713 1593 11747
rect 1593 11713 1627 11747
rect 1627 11713 1636 11747
rect 1584 11704 1636 11713
rect 6460 11704 6512 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 10508 11704 10560 11756
rect 10784 11704 10836 11756
rect 11244 11704 11296 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 2872 11636 2924 11688
rect 3792 11636 3844 11688
rect 4896 11636 4948 11688
rect 5632 11636 5684 11688
rect 6184 11636 6236 11688
rect 9128 11679 9180 11688
rect 5264 11568 5316 11620
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 11704 11636 11756 11688
rect 13544 11704 13596 11756
rect 13820 11704 13872 11756
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 16488 11636 16540 11688
rect 4068 11500 4120 11552
rect 5816 11500 5868 11552
rect 10784 11568 10836 11620
rect 11060 11500 11112 11552
rect 11244 11568 11296 11620
rect 13268 11568 13320 11620
rect 14556 11568 14608 11620
rect 15384 11568 15436 11620
rect 15844 11568 15896 11620
rect 14832 11500 14884 11552
rect 15108 11500 15160 11552
rect 16488 11500 16540 11552
rect 16856 11840 16908 11892
rect 17500 11840 17552 11892
rect 17960 11772 18012 11824
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 18328 11840 18380 11892
rect 18972 11840 19024 11892
rect 19064 11840 19116 11892
rect 19616 11840 19668 11892
rect 20168 11840 20220 11892
rect 20996 11883 21048 11892
rect 20996 11849 21005 11883
rect 21005 11849 21039 11883
rect 21039 11849 21048 11883
rect 20996 11840 21048 11849
rect 21916 11840 21968 11892
rect 24032 11840 24084 11892
rect 18328 11704 18380 11756
rect 19340 11772 19392 11824
rect 19800 11772 19852 11824
rect 21088 11772 21140 11824
rect 22100 11815 22152 11824
rect 22100 11781 22109 11815
rect 22109 11781 22143 11815
rect 22143 11781 22152 11815
rect 22100 11772 22152 11781
rect 22284 11772 22336 11824
rect 23480 11772 23532 11824
rect 23940 11772 23992 11824
rect 34060 11883 34112 11892
rect 34060 11849 34069 11883
rect 34069 11849 34103 11883
rect 34103 11849 34112 11883
rect 34060 11840 34112 11849
rect 19524 11704 19576 11756
rect 19616 11747 19668 11756
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 20628 11704 20680 11756
rect 21732 11704 21784 11756
rect 21916 11704 21968 11756
rect 25320 11772 25372 11824
rect 25688 11772 25740 11824
rect 27068 11772 27120 11824
rect 17592 11636 17644 11645
rect 18236 11636 18288 11688
rect 22468 11636 22520 11688
rect 22928 11636 22980 11688
rect 23112 11679 23164 11688
rect 23112 11645 23121 11679
rect 23121 11645 23155 11679
rect 23155 11645 23164 11679
rect 23112 11636 23164 11645
rect 26700 11704 26752 11756
rect 27252 11704 27304 11756
rect 34796 11772 34848 11824
rect 24584 11679 24636 11688
rect 18972 11568 19024 11620
rect 24584 11645 24593 11679
rect 24593 11645 24627 11679
rect 24627 11645 24636 11679
rect 24584 11636 24636 11645
rect 25136 11636 25188 11688
rect 26332 11636 26384 11688
rect 31668 11636 31720 11688
rect 37464 11679 37516 11688
rect 37464 11645 37473 11679
rect 37473 11645 37507 11679
rect 37507 11645 37516 11679
rect 37464 11636 37516 11645
rect 26976 11568 27028 11620
rect 27160 11568 27212 11620
rect 28540 11568 28592 11620
rect 18144 11500 18196 11552
rect 18420 11500 18472 11552
rect 23756 11500 23808 11552
rect 24032 11500 24084 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 9680 11296 9732 11348
rect 14280 11296 14332 11348
rect 3424 11271 3476 11280
rect 3424 11237 3433 11271
rect 3433 11237 3467 11271
rect 3467 11237 3476 11271
rect 3424 11228 3476 11237
rect 1584 11160 1636 11212
rect 5264 11228 5316 11280
rect 4804 11160 4856 11212
rect 5816 11160 5868 11212
rect 6276 11160 6328 11212
rect 6828 11160 6880 11212
rect 7472 11160 7524 11212
rect 7932 11160 7984 11212
rect 3976 11092 4028 11144
rect 5264 11092 5316 11144
rect 6920 11092 6972 11144
rect 10140 11228 10192 11280
rect 12256 11228 12308 11280
rect 12532 11228 12584 11280
rect 12624 11228 12676 11280
rect 13912 11228 13964 11280
rect 15108 11296 15160 11348
rect 15292 11296 15344 11348
rect 16304 11296 16356 11348
rect 16580 11296 16632 11348
rect 19340 11296 19392 11348
rect 19708 11296 19760 11348
rect 15752 11228 15804 11280
rect 16764 11228 16816 11280
rect 9128 11160 9180 11212
rect 11888 11160 11940 11212
rect 15016 11160 15068 11212
rect 15844 11160 15896 11212
rect 19800 11228 19852 11280
rect 17040 11160 17092 11212
rect 17316 11160 17368 11212
rect 20904 11296 20956 11348
rect 21180 11296 21232 11348
rect 22192 11296 22244 11348
rect 24860 11296 24912 11348
rect 25412 11296 25464 11348
rect 26608 11339 26660 11348
rect 26608 11305 26617 11339
rect 26617 11305 26651 11339
rect 26651 11305 26660 11339
rect 26608 11296 26660 11305
rect 27068 11296 27120 11348
rect 19984 11228 20036 11280
rect 22560 11228 22612 11280
rect 4620 11024 4672 11076
rect 4804 11024 4856 11076
rect 5816 11067 5868 11076
rect 5816 11033 5825 11067
rect 5825 11033 5859 11067
rect 5859 11033 5868 11067
rect 5816 11024 5868 11033
rect 7380 11024 7432 11076
rect 8392 11067 8444 11076
rect 8392 11033 8401 11067
rect 8401 11033 8435 11067
rect 8435 11033 8444 11067
rect 8392 11024 8444 11033
rect 8668 11024 8720 11076
rect 9680 11092 9732 11144
rect 12440 11092 12492 11144
rect 13268 11092 13320 11144
rect 13820 11092 13872 11144
rect 18788 11092 18840 11144
rect 19248 11092 19300 11144
rect 19616 11092 19668 11144
rect 20628 11160 20680 11212
rect 23756 11228 23808 11280
rect 21364 11092 21416 11144
rect 22192 11092 22244 11144
rect 23664 11203 23716 11212
rect 23664 11169 23673 11203
rect 23673 11169 23707 11203
rect 23707 11169 23716 11203
rect 23664 11160 23716 11169
rect 25136 11160 25188 11212
rect 27712 11160 27764 11212
rect 23204 11092 23256 11144
rect 24124 11092 24176 11144
rect 24584 11092 24636 11144
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 25412 11092 25464 11144
rect 26056 11092 26108 11144
rect 26516 11135 26568 11144
rect 26516 11101 26525 11135
rect 26525 11101 26559 11135
rect 26559 11101 26568 11135
rect 26516 11092 26568 11101
rect 27160 11135 27212 11144
rect 27160 11101 27169 11135
rect 27169 11101 27203 11135
rect 27203 11101 27212 11135
rect 27160 11092 27212 11101
rect 7288 10956 7340 11008
rect 9312 10956 9364 11008
rect 9496 10956 9548 11008
rect 10416 10956 10468 11008
rect 11060 11024 11112 11076
rect 12808 11024 12860 11076
rect 14004 11024 14056 11076
rect 14556 11067 14608 11076
rect 14556 11033 14565 11067
rect 14565 11033 14599 11067
rect 14599 11033 14608 11067
rect 14556 11024 14608 11033
rect 14832 11024 14884 11076
rect 15844 11024 15896 11076
rect 16580 11024 16632 11076
rect 17500 11024 17552 11076
rect 18052 11067 18104 11076
rect 18052 11033 18061 11067
rect 18061 11033 18095 11067
rect 18095 11033 18104 11067
rect 18052 11024 18104 11033
rect 18236 11024 18288 11076
rect 13544 10956 13596 11008
rect 18972 11024 19024 11076
rect 19524 11024 19576 11076
rect 19984 11024 20036 11076
rect 20168 11067 20220 11076
rect 20168 11033 20177 11067
rect 20177 11033 20211 11067
rect 20211 11033 20220 11067
rect 20168 11024 20220 11033
rect 20260 11067 20312 11076
rect 20260 11033 20269 11067
rect 20269 11033 20303 11067
rect 20303 11033 20312 11067
rect 20260 11024 20312 11033
rect 20720 11024 20772 11076
rect 23112 11024 23164 11076
rect 23480 11067 23532 11076
rect 23480 11033 23489 11067
rect 23489 11033 23523 11067
rect 23523 11033 23532 11067
rect 23480 11024 23532 11033
rect 28356 11024 28408 11076
rect 34796 11024 34848 11076
rect 35900 11024 35952 11076
rect 18512 10956 18564 11008
rect 22008 10956 22060 11008
rect 24584 10999 24636 11008
rect 24584 10965 24593 10999
rect 24593 10965 24627 10999
rect 24627 10965 24636 10999
rect 24584 10956 24636 10965
rect 24860 10956 24912 11008
rect 25872 10956 25924 11008
rect 27896 10999 27948 11008
rect 27896 10965 27905 10999
rect 27905 10965 27939 10999
rect 27939 10965 27948 10999
rect 27896 10956 27948 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1584 10752 1636 10804
rect 3976 10752 4028 10804
rect 1952 10684 2004 10736
rect 3608 10684 3660 10736
rect 6644 10752 6696 10804
rect 13544 10752 13596 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 3976 10659 4028 10668
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4620 10548 4672 10600
rect 8024 10616 8076 10668
rect 8300 10616 8352 10668
rect 9312 10684 9364 10736
rect 9680 10684 9732 10736
rect 11704 10684 11756 10736
rect 12072 10684 12124 10736
rect 12624 10684 12676 10736
rect 13728 10684 13780 10736
rect 14464 10727 14516 10736
rect 14464 10693 14473 10727
rect 14473 10693 14507 10727
rect 14507 10693 14516 10727
rect 14464 10684 14516 10693
rect 17684 10752 17736 10804
rect 17868 10752 17920 10804
rect 15200 10684 15252 10736
rect 15476 10684 15528 10736
rect 15844 10684 15896 10736
rect 16304 10727 16356 10736
rect 16304 10693 16313 10727
rect 16313 10693 16347 10727
rect 16347 10693 16356 10727
rect 16304 10684 16356 10693
rect 16948 10727 17000 10736
rect 16948 10693 16957 10727
rect 16957 10693 16991 10727
rect 16991 10693 17000 10727
rect 16948 10684 17000 10693
rect 18512 10752 18564 10804
rect 18880 10684 18932 10736
rect 19248 10684 19300 10736
rect 19340 10684 19392 10736
rect 20168 10684 20220 10736
rect 10784 10616 10836 10668
rect 10968 10616 11020 10668
rect 11888 10659 11940 10668
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 9128 10591 9180 10600
rect 9128 10557 9137 10591
rect 9137 10557 9171 10591
rect 9171 10557 9180 10591
rect 9128 10548 9180 10557
rect 10048 10548 10100 10600
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 17960 10616 18012 10668
rect 18236 10616 18288 10668
rect 18328 10616 18380 10668
rect 20720 10684 20772 10736
rect 21548 10684 21600 10736
rect 22008 10752 22060 10804
rect 22744 10752 22796 10804
rect 23480 10752 23532 10804
rect 26148 10795 26200 10804
rect 25044 10727 25096 10736
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 22468 10616 22520 10668
rect 17224 10591 17276 10600
rect 11704 10480 11756 10532
rect 11888 10480 11940 10532
rect 16580 10480 16632 10532
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 17316 10548 17368 10600
rect 18420 10548 18472 10600
rect 18512 10548 18564 10600
rect 19064 10591 19116 10600
rect 19064 10557 19073 10591
rect 19073 10557 19107 10591
rect 19107 10557 19116 10591
rect 19064 10548 19116 10557
rect 19984 10548 20036 10600
rect 20628 10548 20680 10600
rect 20996 10548 21048 10600
rect 23112 10616 23164 10668
rect 25044 10693 25053 10727
rect 25053 10693 25087 10727
rect 25087 10693 25096 10727
rect 25044 10684 25096 10693
rect 26148 10761 26157 10795
rect 26157 10761 26191 10795
rect 26191 10761 26200 10795
rect 26148 10752 26200 10761
rect 28172 10684 28224 10736
rect 38384 10684 38436 10736
rect 25688 10616 25740 10668
rect 26700 10616 26752 10668
rect 38108 10659 38160 10668
rect 38108 10625 38117 10659
rect 38117 10625 38151 10659
rect 38151 10625 38160 10659
rect 38108 10616 38160 10625
rect 24032 10548 24084 10600
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 25136 10548 25188 10600
rect 25412 10548 25464 10600
rect 26148 10548 26200 10600
rect 14188 10412 14240 10464
rect 25872 10480 25924 10532
rect 27160 10480 27212 10532
rect 20352 10412 20404 10464
rect 22468 10412 22520 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2136 10208 2188 10260
rect 3884 10208 3936 10260
rect 4620 10208 4672 10260
rect 7104 10208 7156 10260
rect 14832 10208 14884 10260
rect 14924 10208 14976 10260
rect 17224 10208 17276 10260
rect 1584 10072 1636 10124
rect 3240 10072 3292 10124
rect 4620 10072 4672 10124
rect 6644 10072 6696 10124
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 8760 10140 8812 10192
rect 10508 10140 10560 10192
rect 11060 10140 11112 10192
rect 11520 10140 11572 10192
rect 13176 10140 13228 10192
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 12440 10072 12492 10124
rect 12716 10072 12768 10124
rect 13544 10072 13596 10124
rect 13912 10140 13964 10192
rect 14188 10140 14240 10192
rect 15660 10140 15712 10192
rect 17684 10208 17736 10260
rect 17776 10208 17828 10260
rect 17960 10208 18012 10260
rect 18236 10208 18288 10260
rect 21640 10208 21692 10260
rect 22376 10208 22428 10260
rect 23020 10208 23072 10260
rect 25320 10251 25372 10260
rect 25320 10217 25329 10251
rect 25329 10217 25363 10251
rect 25363 10217 25372 10251
rect 25320 10208 25372 10217
rect 30104 10208 30156 10260
rect 17408 10140 17460 10192
rect 14832 10072 14884 10124
rect 16304 10072 16356 10124
rect 16488 10072 16540 10124
rect 17776 10072 17828 10124
rect 18512 10072 18564 10124
rect 19064 10140 19116 10192
rect 23204 10140 23256 10192
rect 23940 10183 23992 10192
rect 23940 10149 23949 10183
rect 23949 10149 23983 10183
rect 23983 10149 23992 10183
rect 23940 10140 23992 10149
rect 27804 10140 27856 10192
rect 19156 10072 19208 10124
rect 11520 10004 11572 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 15292 10004 15344 10056
rect 17316 10004 17368 10056
rect 17500 10004 17552 10056
rect 5632 9936 5684 9988
rect 7472 9936 7524 9988
rect 7932 9979 7984 9988
rect 7932 9945 7941 9979
rect 7941 9945 7975 9979
rect 7975 9945 7984 9979
rect 7932 9936 7984 9945
rect 8116 9936 8168 9988
rect 11060 9936 11112 9988
rect 11612 9936 11664 9988
rect 12256 9936 12308 9988
rect 13728 9979 13780 9988
rect 13728 9945 13737 9979
rect 13737 9945 13771 9979
rect 13771 9945 13780 9979
rect 13728 9936 13780 9945
rect 14372 9936 14424 9988
rect 15200 9936 15252 9988
rect 15936 9936 15988 9988
rect 16304 9936 16356 9988
rect 16672 9979 16724 9988
rect 16672 9945 16681 9979
rect 16681 9945 16715 9979
rect 16715 9945 16724 9979
rect 16672 9936 16724 9945
rect 20444 10072 20496 10124
rect 16028 9868 16080 9920
rect 16212 9868 16264 9920
rect 17224 9868 17276 9920
rect 17408 9868 17460 9920
rect 17960 9868 18012 9920
rect 18052 9868 18104 9920
rect 18512 9936 18564 9988
rect 19892 10004 19944 10056
rect 22284 10072 22336 10124
rect 20812 10004 20864 10056
rect 21088 10004 21140 10056
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 22376 10004 22428 10056
rect 27252 10072 27304 10124
rect 25504 10004 25556 10056
rect 25872 10047 25924 10056
rect 25872 10013 25881 10047
rect 25881 10013 25915 10047
rect 25915 10013 25924 10047
rect 25872 10004 25924 10013
rect 34428 10004 34480 10056
rect 37188 10004 37240 10056
rect 37740 10047 37792 10056
rect 37740 10013 37749 10047
rect 37749 10013 37783 10047
rect 37783 10013 37792 10047
rect 37740 10004 37792 10013
rect 21824 9936 21876 9988
rect 19156 9868 19208 9920
rect 21180 9868 21232 9920
rect 23296 9868 23348 9920
rect 24032 9936 24084 9988
rect 27896 9936 27948 9988
rect 25412 9868 25464 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3792 9664 3844 9716
rect 1400 9596 1452 9648
rect 2136 9596 2188 9648
rect 3976 9596 4028 9648
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 6276 9528 6328 9580
rect 8484 9596 8536 9648
rect 13728 9664 13780 9716
rect 24676 9664 24728 9716
rect 25044 9664 25096 9716
rect 10416 9596 10468 9648
rect 12256 9596 12308 9648
rect 13636 9596 13688 9648
rect 4436 9460 4488 9512
rect 4712 9460 4764 9512
rect 2228 9324 2280 9376
rect 2504 9324 2556 9376
rect 6092 9324 6144 9376
rect 7840 9460 7892 9512
rect 9128 9528 9180 9580
rect 10140 9460 10192 9512
rect 10232 9460 10284 9512
rect 9128 9392 9180 9444
rect 11704 9460 11756 9512
rect 14648 9596 14700 9648
rect 8300 9367 8352 9376
rect 8300 9333 8309 9367
rect 8309 9333 8343 9367
rect 8343 9333 8352 9367
rect 8300 9324 8352 9333
rect 8576 9324 8628 9376
rect 8668 9324 8720 9376
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 11980 9324 12032 9376
rect 12348 9324 12400 9376
rect 12532 9324 12584 9376
rect 14372 9324 14424 9376
rect 15108 9392 15160 9444
rect 16028 9596 16080 9648
rect 16304 9639 16356 9648
rect 16304 9605 16313 9639
rect 16313 9605 16347 9639
rect 16347 9605 16356 9639
rect 16304 9596 16356 9605
rect 16764 9596 16816 9648
rect 18236 9596 18288 9648
rect 18328 9596 18380 9648
rect 19248 9596 19300 9648
rect 19340 9596 19392 9648
rect 19708 9596 19760 9648
rect 16488 9528 16540 9580
rect 15660 9460 15712 9512
rect 16028 9460 16080 9512
rect 16856 9528 16908 9580
rect 17224 9528 17276 9580
rect 15292 9392 15344 9444
rect 18236 9460 18288 9512
rect 18420 9460 18472 9512
rect 18604 9460 18656 9512
rect 18880 9460 18932 9512
rect 19708 9503 19760 9512
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 21180 9596 21232 9648
rect 20904 9528 20956 9580
rect 21548 9596 21600 9648
rect 21916 9596 21968 9648
rect 22284 9596 22336 9648
rect 25412 9596 25464 9648
rect 28724 9596 28776 9648
rect 21640 9528 21692 9580
rect 25596 9528 25648 9580
rect 19708 9460 19760 9469
rect 21548 9460 21600 9512
rect 24492 9460 24544 9512
rect 24676 9460 24728 9512
rect 18328 9392 18380 9444
rect 19616 9392 19668 9444
rect 19800 9392 19852 9444
rect 22284 9392 22336 9444
rect 23204 9392 23256 9444
rect 24584 9392 24636 9444
rect 26148 9460 26200 9512
rect 28816 9528 28868 9580
rect 29736 9460 29788 9512
rect 20904 9324 20956 9376
rect 21548 9324 21600 9376
rect 22192 9324 22244 9376
rect 22652 9324 22704 9376
rect 27344 9324 27396 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1676 9120 1728 9172
rect 8300 9120 8352 9172
rect 12624 9120 12676 9172
rect 12808 9120 12860 9172
rect 13636 9120 13688 9172
rect 13912 9120 13964 9172
rect 14556 9120 14608 9172
rect 14740 9120 14792 9172
rect 15660 9120 15712 9172
rect 3056 9052 3108 9104
rect 3700 9052 3752 9104
rect 5540 9052 5592 9104
rect 6828 9052 6880 9104
rect 10784 9052 10836 9104
rect 4252 8984 4304 9036
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 7564 8984 7616 9036
rect 9496 8984 9548 9036
rect 10692 8984 10744 9036
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 3976 8848 4028 8900
rect 4160 8848 4212 8900
rect 4344 8848 4396 8900
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 6000 8848 6052 8857
rect 7564 8848 7616 8900
rect 9312 8891 9364 8900
rect 9312 8857 9321 8891
rect 9321 8857 9355 8891
rect 9355 8857 9364 8891
rect 9312 8848 9364 8857
rect 9496 8848 9548 8900
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 13912 8984 13964 9036
rect 14740 8984 14792 9036
rect 16764 8984 16816 9036
rect 17408 9052 17460 9104
rect 18328 9052 18380 9104
rect 18696 9120 18748 9172
rect 19616 9120 19668 9172
rect 20628 9120 20680 9172
rect 20720 9120 20772 9172
rect 21180 9120 21232 9172
rect 21916 9120 21968 9172
rect 22192 9120 22244 9172
rect 21548 9052 21600 9104
rect 12532 8916 12584 8968
rect 13084 8916 13136 8968
rect 15476 8916 15528 8968
rect 17592 8984 17644 9036
rect 18788 9027 18840 9036
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 18972 8984 19024 9036
rect 11520 8891 11572 8900
rect 11520 8857 11529 8891
rect 11529 8857 11563 8891
rect 11563 8857 11572 8891
rect 11520 8848 11572 8857
rect 12072 8848 12124 8900
rect 14372 8848 14424 8900
rect 14740 8848 14792 8900
rect 8116 8780 8168 8832
rect 8576 8780 8628 8832
rect 16120 8780 16172 8832
rect 16488 8848 16540 8900
rect 19524 8916 19576 8968
rect 19984 8916 20036 8968
rect 21364 8916 21416 8968
rect 17684 8848 17736 8900
rect 18972 8848 19024 8900
rect 19064 8848 19116 8900
rect 19340 8848 19392 8900
rect 20260 8891 20312 8900
rect 20260 8857 20269 8891
rect 20269 8857 20303 8891
rect 20303 8857 20312 8891
rect 20812 8891 20864 8900
rect 20260 8848 20312 8857
rect 20812 8857 20821 8891
rect 20821 8857 20855 8891
rect 20855 8857 20864 8891
rect 20812 8848 20864 8857
rect 21180 8848 21232 8900
rect 23204 8916 23256 8968
rect 25780 9052 25832 9104
rect 37556 9052 37608 9104
rect 26976 8984 27028 9036
rect 38016 8959 38068 8968
rect 22560 8891 22612 8900
rect 22560 8857 22569 8891
rect 22569 8857 22603 8891
rect 22603 8857 22612 8891
rect 22560 8848 22612 8857
rect 22652 8891 22704 8900
rect 22652 8857 22661 8891
rect 22661 8857 22695 8891
rect 22695 8857 22704 8891
rect 38016 8925 38025 8959
rect 38025 8925 38059 8959
rect 38059 8925 38068 8959
rect 38016 8916 38068 8925
rect 27252 8891 27304 8900
rect 22652 8848 22704 8857
rect 21364 8780 21416 8832
rect 21640 8780 21692 8832
rect 27252 8857 27261 8891
rect 27261 8857 27295 8891
rect 27295 8857 27304 8891
rect 27252 8848 27304 8857
rect 27344 8891 27396 8900
rect 27344 8857 27353 8891
rect 27353 8857 27387 8891
rect 27387 8857 27396 8891
rect 27344 8848 27396 8857
rect 23756 8823 23808 8832
rect 23756 8789 23765 8823
rect 23765 8789 23799 8823
rect 23799 8789 23808 8823
rect 23756 8780 23808 8789
rect 25596 8823 25648 8832
rect 25596 8789 25605 8823
rect 25605 8789 25639 8823
rect 25639 8789 25648 8823
rect 25596 8780 25648 8789
rect 25688 8780 25740 8832
rect 27620 8780 27672 8832
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4620 8508 4672 8560
rect 9220 8576 9272 8628
rect 7196 8508 7248 8560
rect 8576 8508 8628 8560
rect 13268 8576 13320 8628
rect 14004 8576 14056 8628
rect 14832 8576 14884 8628
rect 10048 8508 10100 8560
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 5632 8440 5684 8492
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 4160 8372 4212 8424
rect 6920 8415 6972 8424
rect 4068 8304 4120 8356
rect 5632 8304 5684 8356
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 11888 8508 11940 8560
rect 12532 8508 12584 8560
rect 11336 8440 11388 8492
rect 15292 8508 15344 8560
rect 16488 8576 16540 8628
rect 17132 8576 17184 8628
rect 15476 8508 15528 8560
rect 17316 8508 17368 8560
rect 18236 8551 18288 8560
rect 18236 8517 18245 8551
rect 18245 8517 18279 8551
rect 18279 8517 18288 8551
rect 18236 8508 18288 8517
rect 18512 8508 18564 8560
rect 19248 8576 19300 8628
rect 20260 8576 20312 8628
rect 21364 8576 21416 8628
rect 29000 8619 29052 8628
rect 29000 8585 29009 8619
rect 29009 8585 29043 8619
rect 29043 8585 29052 8619
rect 29000 8576 29052 8585
rect 20352 8508 20404 8560
rect 3884 8236 3936 8288
rect 4988 8236 5040 8288
rect 6828 8236 6880 8288
rect 7748 8236 7800 8288
rect 9864 8236 9916 8288
rect 10140 8236 10192 8288
rect 10876 8236 10928 8288
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 13360 8440 13412 8492
rect 14004 8440 14056 8492
rect 14280 8440 14332 8492
rect 14464 8440 14516 8492
rect 20812 8440 20864 8492
rect 21916 8440 21968 8492
rect 12992 8304 13044 8356
rect 13636 8304 13688 8356
rect 15844 8372 15896 8424
rect 16396 8372 16448 8424
rect 16580 8372 16632 8424
rect 17316 8372 17368 8424
rect 14188 8236 14240 8288
rect 14832 8236 14884 8288
rect 17592 8304 17644 8356
rect 17868 8372 17920 8424
rect 18696 8372 18748 8424
rect 19064 8372 19116 8424
rect 21548 8372 21600 8424
rect 22376 8508 22428 8560
rect 23020 8508 23072 8560
rect 23572 8508 23624 8560
rect 23664 8440 23716 8492
rect 23848 8483 23900 8492
rect 23848 8449 23857 8483
rect 23857 8449 23891 8483
rect 23891 8449 23900 8483
rect 23848 8440 23900 8449
rect 24584 8440 24636 8492
rect 25044 8483 25096 8492
rect 25044 8449 25053 8483
rect 25053 8449 25087 8483
rect 25087 8449 25096 8483
rect 25044 8440 25096 8449
rect 25504 8483 25556 8492
rect 25504 8449 25513 8483
rect 25513 8449 25547 8483
rect 25547 8449 25556 8483
rect 25504 8440 25556 8449
rect 29736 8440 29788 8492
rect 18512 8236 18564 8288
rect 18696 8236 18748 8288
rect 19340 8236 19392 8288
rect 19800 8304 19852 8356
rect 22192 8304 22244 8356
rect 21088 8236 21140 8288
rect 22744 8372 22796 8424
rect 23388 8415 23440 8424
rect 23388 8381 23397 8415
rect 23397 8381 23431 8415
rect 23431 8381 23440 8415
rect 23388 8372 23440 8381
rect 23480 8372 23532 8424
rect 23112 8304 23164 8356
rect 24676 8304 24728 8356
rect 23388 8236 23440 8288
rect 23572 8236 23624 8288
rect 30840 8236 30892 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3148 8032 3200 8084
rect 8668 8032 8720 8084
rect 11704 8032 11756 8084
rect 13176 8032 13228 8084
rect 13728 8032 13780 8084
rect 14372 8032 14424 8084
rect 14648 8032 14700 8084
rect 17776 8032 17828 8084
rect 18420 8032 18472 8084
rect 3700 7964 3752 8016
rect 4988 7964 5040 8016
rect 6920 7964 6972 8016
rect 7104 7964 7156 8016
rect 3332 7896 3384 7948
rect 3884 7896 3936 7948
rect 4620 7896 4672 7948
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6276 7896 6328 7948
rect 7380 7896 7432 7948
rect 7748 7896 7800 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 4804 7828 4856 7880
rect 5448 7828 5500 7880
rect 11612 7964 11664 8016
rect 11336 7896 11388 7948
rect 12900 7964 12952 8016
rect 9128 7828 9180 7880
rect 11888 7896 11940 7948
rect 13452 7896 13504 7948
rect 16948 7964 17000 8016
rect 17408 7964 17460 8016
rect 16672 7896 16724 7948
rect 16856 7896 16908 7948
rect 17960 7896 18012 7948
rect 18512 7964 18564 8016
rect 18880 8032 18932 8084
rect 22468 8032 22520 8084
rect 26240 8075 26292 8084
rect 26240 8041 26249 8075
rect 26249 8041 26283 8075
rect 26283 8041 26292 8075
rect 26240 8032 26292 8041
rect 33968 8032 34020 8084
rect 20260 7964 20312 8016
rect 4620 7760 4672 7812
rect 5724 7760 5776 7812
rect 2780 7692 2832 7744
rect 9680 7803 9732 7812
rect 9680 7769 9689 7803
rect 9689 7769 9723 7803
rect 9723 7769 9732 7803
rect 9680 7760 9732 7769
rect 10140 7760 10192 7812
rect 10968 7760 11020 7812
rect 6000 7692 6052 7744
rect 8760 7692 8812 7744
rect 9220 7692 9272 7744
rect 11888 7692 11940 7744
rect 12900 7760 12952 7812
rect 13268 7760 13320 7812
rect 13636 7803 13688 7812
rect 13636 7769 13645 7803
rect 13645 7769 13679 7803
rect 13679 7769 13688 7803
rect 13636 7760 13688 7769
rect 13912 7828 13964 7880
rect 17500 7828 17552 7880
rect 14648 7760 14700 7812
rect 13176 7692 13228 7744
rect 13820 7692 13872 7744
rect 14740 7692 14792 7744
rect 14832 7692 14884 7744
rect 16304 7692 16356 7744
rect 16672 7803 16724 7812
rect 16672 7769 16681 7803
rect 16681 7769 16715 7803
rect 16715 7769 16724 7803
rect 19892 7896 19944 7948
rect 20720 7964 20772 8016
rect 21180 7896 21232 7948
rect 16672 7760 16724 7769
rect 17776 7692 17828 7744
rect 19616 7760 19668 7812
rect 21088 7828 21140 7880
rect 24216 7964 24268 8016
rect 21548 7828 21600 7880
rect 26424 7964 26476 8016
rect 24676 7896 24728 7948
rect 22008 7871 22060 7880
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 22100 7828 22152 7880
rect 23204 7828 23256 7880
rect 23388 7828 23440 7880
rect 26148 7871 26200 7880
rect 26148 7837 26157 7871
rect 26157 7837 26191 7871
rect 26191 7837 26200 7871
rect 26148 7828 26200 7837
rect 38292 7871 38344 7880
rect 38292 7837 38301 7871
rect 38301 7837 38335 7871
rect 38335 7837 38344 7871
rect 38292 7828 38344 7837
rect 21180 7760 21232 7812
rect 23572 7760 23624 7812
rect 19984 7692 20036 7744
rect 20996 7692 21048 7744
rect 25596 7760 25648 7812
rect 24952 7692 25004 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5724 7488 5776 7540
rect 4528 7420 4580 7472
rect 5172 7420 5224 7472
rect 6368 7420 6420 7472
rect 6552 7420 6604 7472
rect 7380 7420 7432 7472
rect 7932 7463 7984 7472
rect 7932 7429 7941 7463
rect 7941 7429 7975 7463
rect 7975 7429 7984 7463
rect 7932 7420 7984 7429
rect 9864 7420 9916 7472
rect 10232 7488 10284 7540
rect 12072 7488 12124 7540
rect 10876 7420 10928 7472
rect 11244 7420 11296 7472
rect 11336 7420 11388 7472
rect 13544 7420 13596 7472
rect 15200 7488 15252 7540
rect 16488 7488 16540 7540
rect 16856 7488 16908 7540
rect 16948 7488 17000 7540
rect 18512 7488 18564 7540
rect 18788 7488 18840 7540
rect 23112 7488 23164 7540
rect 24492 7531 24544 7540
rect 24492 7497 24501 7531
rect 24501 7497 24535 7531
rect 24535 7497 24544 7531
rect 24492 7488 24544 7497
rect 24860 7531 24912 7540
rect 24860 7497 24869 7531
rect 24869 7497 24903 7531
rect 24903 7497 24912 7531
rect 24860 7488 24912 7497
rect 37464 7488 37516 7540
rect 17868 7420 17920 7472
rect 18144 7420 18196 7472
rect 4804 7352 4856 7404
rect 1676 7284 1728 7336
rect 3332 7284 3384 7336
rect 4160 7284 4212 7336
rect 5264 7284 5316 7336
rect 5540 7284 5592 7336
rect 6276 7284 6328 7336
rect 6000 7216 6052 7268
rect 9220 7352 9272 7404
rect 7104 7284 7156 7336
rect 9312 7284 9364 7336
rect 10508 7352 10560 7404
rect 11152 7352 11204 7404
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 15476 7352 15528 7404
rect 15844 7352 15896 7404
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 10508 7216 10560 7268
rect 11612 7216 11664 7268
rect 14188 7327 14240 7336
rect 13452 7259 13504 7268
rect 13452 7225 13461 7259
rect 13461 7225 13495 7259
rect 13495 7225 13504 7259
rect 13452 7216 13504 7225
rect 4528 7148 4580 7200
rect 11060 7148 11112 7200
rect 11796 7148 11848 7200
rect 12348 7148 12400 7200
rect 12532 7148 12584 7200
rect 13912 7148 13964 7200
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 17040 7284 17092 7336
rect 18512 7352 18564 7404
rect 18604 7352 18656 7404
rect 19064 7352 19116 7404
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18236 7284 18288 7336
rect 16212 7148 16264 7200
rect 18144 7216 18196 7268
rect 18512 7216 18564 7268
rect 20812 7420 20864 7472
rect 21548 7420 21600 7472
rect 22836 7420 22888 7472
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 21640 7352 21692 7404
rect 23204 7352 23256 7404
rect 25964 7420 26016 7472
rect 26608 7352 26660 7404
rect 38108 7395 38160 7404
rect 38108 7361 38117 7395
rect 38117 7361 38151 7395
rect 38151 7361 38160 7395
rect 38108 7352 38160 7361
rect 17868 7148 17920 7200
rect 18788 7148 18840 7200
rect 18880 7148 18932 7200
rect 20628 7216 20680 7268
rect 21088 7216 21140 7268
rect 21364 7259 21416 7268
rect 21364 7225 21373 7259
rect 21373 7225 21407 7259
rect 21407 7225 21416 7259
rect 21364 7216 21416 7225
rect 24584 7284 24636 7336
rect 24492 7216 24544 7268
rect 19984 7148 20036 7200
rect 22008 7148 22060 7200
rect 22744 7191 22796 7200
rect 22744 7157 22753 7191
rect 22753 7157 22787 7191
rect 22787 7157 22796 7191
rect 22744 7148 22796 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3516 6944 3568 6996
rect 4620 6944 4672 6996
rect 9036 6944 9088 6996
rect 6368 6876 6420 6928
rect 8116 6876 8168 6928
rect 9128 6876 9180 6928
rect 1584 6808 1636 6860
rect 3240 6808 3292 6860
rect 4528 6851 4580 6860
rect 4528 6817 4537 6851
rect 4537 6817 4571 6851
rect 4571 6817 4580 6851
rect 4528 6808 4580 6817
rect 5448 6808 5500 6860
rect 6276 6740 6328 6792
rect 7104 6808 7156 6860
rect 12072 6944 12124 6996
rect 10692 6808 10744 6860
rect 12624 6876 12676 6928
rect 13268 6876 13320 6928
rect 14004 6876 14056 6928
rect 15844 6944 15896 6996
rect 17040 6944 17092 6996
rect 17132 6944 17184 6996
rect 17868 6944 17920 6996
rect 19064 6944 19116 6996
rect 18144 6876 18196 6928
rect 20076 6944 20128 6996
rect 22744 6944 22796 6996
rect 4068 6672 4120 6724
rect 4804 6715 4856 6724
rect 4804 6681 4813 6715
rect 4813 6681 4847 6715
rect 4847 6681 4856 6715
rect 4804 6672 4856 6681
rect 6644 6672 6696 6724
rect 7012 6715 7064 6724
rect 7012 6681 7021 6715
rect 7021 6681 7055 6715
rect 7055 6681 7064 6715
rect 7012 6672 7064 6681
rect 7472 6672 7524 6724
rect 1860 6604 1912 6656
rect 4160 6604 4212 6656
rect 9312 6740 9364 6792
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 10416 6783 10468 6792
rect 9680 6740 9732 6749
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 9128 6672 9180 6724
rect 10692 6715 10744 6724
rect 10692 6681 10701 6715
rect 10701 6681 10735 6715
rect 10735 6681 10744 6715
rect 10692 6672 10744 6681
rect 12808 6740 12860 6792
rect 14280 6740 14332 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 15108 6783 15160 6792
rect 14556 6740 14608 6749
rect 12624 6672 12676 6724
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 17132 6808 17184 6860
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 18052 6808 18104 6860
rect 19248 6808 19300 6860
rect 20168 6851 20220 6860
rect 15660 6740 15712 6792
rect 15844 6740 15896 6792
rect 16212 6740 16264 6792
rect 18604 6740 18656 6792
rect 18880 6740 18932 6792
rect 19616 6740 19668 6792
rect 20168 6817 20177 6851
rect 20177 6817 20211 6851
rect 20211 6817 20220 6851
rect 20168 6808 20220 6817
rect 21180 6808 21232 6860
rect 9220 6604 9272 6656
rect 9956 6604 10008 6656
rect 10600 6604 10652 6656
rect 11060 6604 11112 6656
rect 11612 6604 11664 6656
rect 12532 6604 12584 6656
rect 12808 6604 12860 6656
rect 14188 6604 14240 6656
rect 14280 6604 14332 6656
rect 16120 6604 16172 6656
rect 19064 6672 19116 6724
rect 20720 6783 20772 6792
rect 20720 6749 20729 6783
rect 20729 6749 20763 6783
rect 20763 6749 20772 6783
rect 20720 6740 20772 6749
rect 20996 6740 21048 6792
rect 22284 6876 22336 6928
rect 23388 6851 23440 6860
rect 23388 6817 23397 6851
rect 23397 6817 23431 6851
rect 23431 6817 23440 6851
rect 23388 6808 23440 6817
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 27252 6808 27304 6860
rect 31024 6808 31076 6860
rect 22100 6740 22152 6792
rect 20812 6672 20864 6724
rect 23756 6740 23808 6792
rect 25872 6783 25924 6792
rect 25872 6749 25881 6783
rect 25881 6749 25915 6783
rect 25915 6749 25924 6783
rect 25872 6740 25924 6749
rect 30380 6740 30432 6792
rect 35716 6740 35768 6792
rect 19432 6604 19484 6656
rect 20536 6604 20588 6656
rect 22100 6647 22152 6656
rect 22100 6613 22109 6647
rect 22109 6613 22143 6647
rect 22143 6613 22152 6647
rect 22744 6647 22796 6656
rect 22100 6604 22152 6613
rect 22744 6613 22753 6647
rect 22753 6613 22787 6647
rect 22787 6613 22796 6647
rect 22744 6604 22796 6613
rect 23296 6604 23348 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4528 6400 4580 6452
rect 7472 6400 7524 6452
rect 8208 6400 8260 6452
rect 10048 6400 10100 6452
rect 2320 6375 2372 6384
rect 2320 6341 2329 6375
rect 2329 6341 2363 6375
rect 2363 6341 2372 6375
rect 2320 6332 2372 6341
rect 4160 6332 4212 6384
rect 5724 6332 5776 6384
rect 7104 6332 7156 6384
rect 3976 6264 4028 6316
rect 8668 6332 8720 6384
rect 9680 6332 9732 6384
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 10876 6400 10928 6452
rect 10968 6332 11020 6384
rect 12164 6400 12216 6452
rect 18880 6400 18932 6452
rect 19248 6400 19300 6452
rect 19708 6400 19760 6452
rect 13728 6332 13780 6384
rect 14188 6375 14240 6384
rect 14188 6341 14197 6375
rect 14197 6341 14231 6375
rect 14231 6341 14240 6375
rect 14188 6332 14240 6341
rect 15384 6332 15436 6384
rect 16580 6332 16632 6384
rect 17132 6332 17184 6384
rect 21180 6400 21232 6452
rect 22284 6443 22336 6452
rect 22284 6409 22293 6443
rect 22293 6409 22327 6443
rect 22327 6409 22336 6443
rect 22284 6400 22336 6409
rect 23572 6443 23624 6452
rect 23572 6409 23581 6443
rect 23581 6409 23615 6443
rect 23615 6409 23624 6443
rect 23572 6400 23624 6409
rect 24400 6400 24452 6452
rect 20076 6375 20128 6384
rect 20076 6341 20085 6375
rect 20085 6341 20119 6375
rect 20119 6341 20128 6375
rect 20076 6332 20128 6341
rect 20168 6332 20220 6384
rect 20720 6332 20772 6384
rect 20904 6332 20956 6384
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 9496 6264 9548 6316
rect 10508 6264 10560 6316
rect 11612 6264 11664 6316
rect 16488 6264 16540 6316
rect 17592 6307 17644 6316
rect 17592 6273 17601 6307
rect 17601 6273 17635 6307
rect 17635 6273 17644 6307
rect 17592 6264 17644 6273
rect 17776 6264 17828 6316
rect 18144 6264 18196 6316
rect 18604 6264 18656 6316
rect 19064 6264 19116 6316
rect 19616 6264 19668 6316
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 3700 6128 3752 6180
rect 4988 6128 5040 6180
rect 5448 6128 5500 6180
rect 8116 6128 8168 6180
rect 3424 6060 3476 6112
rect 7840 6060 7892 6112
rect 10692 6196 10744 6248
rect 10876 6196 10928 6248
rect 10968 6128 11020 6180
rect 13268 6196 13320 6248
rect 15108 6196 15160 6248
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 20260 6264 20312 6316
rect 20444 6264 20496 6316
rect 21180 6264 21232 6316
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 22468 6332 22520 6384
rect 9680 6060 9732 6112
rect 22560 6196 22612 6248
rect 14648 6060 14700 6112
rect 16856 6060 16908 6112
rect 20996 6128 21048 6180
rect 21364 6171 21416 6180
rect 21364 6137 21373 6171
rect 21373 6137 21407 6171
rect 21407 6137 21416 6171
rect 21364 6128 21416 6137
rect 35808 6264 35860 6316
rect 17500 6060 17552 6112
rect 19248 6060 19300 6112
rect 20168 6060 20220 6112
rect 20444 6060 20496 6112
rect 38016 6128 38068 6180
rect 22928 6060 22980 6112
rect 23112 6103 23164 6112
rect 23112 6069 23121 6103
rect 23121 6069 23155 6103
rect 23155 6069 23164 6103
rect 23112 6060 23164 6069
rect 24952 6060 25004 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3056 5856 3108 5908
rect 3424 5856 3476 5908
rect 3976 5856 4028 5908
rect 6736 5856 6788 5908
rect 7012 5856 7064 5908
rect 5356 5788 5408 5840
rect 5724 5831 5776 5840
rect 5724 5797 5733 5831
rect 5733 5797 5767 5831
rect 5767 5797 5776 5831
rect 5724 5788 5776 5797
rect 8484 5856 8536 5908
rect 9036 5856 9088 5908
rect 9404 5856 9456 5908
rect 10324 5856 10376 5908
rect 16856 5856 16908 5908
rect 17040 5856 17092 5908
rect 17868 5856 17920 5908
rect 18696 5856 18748 5908
rect 18880 5856 18932 5908
rect 19984 5856 20036 5908
rect 20352 5856 20404 5908
rect 20720 5856 20772 5908
rect 21732 5856 21784 5908
rect 23848 5856 23900 5908
rect 37556 5856 37608 5908
rect 12348 5831 12400 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 4988 5720 5040 5772
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 11244 5720 11296 5772
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 7840 5652 7892 5704
rect 8668 5652 8720 5704
rect 9128 5695 9180 5704
rect 9128 5661 9137 5695
rect 9137 5661 9171 5695
rect 9171 5661 9180 5695
rect 9956 5695 10008 5704
rect 9128 5652 9180 5661
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 10048 5652 10100 5704
rect 6828 5584 6880 5636
rect 10324 5584 10376 5636
rect 10784 5652 10836 5704
rect 12348 5797 12357 5831
rect 12357 5797 12391 5831
rect 12391 5797 12400 5831
rect 12348 5788 12400 5797
rect 12532 5788 12584 5840
rect 14004 5788 14056 5840
rect 14372 5831 14424 5840
rect 14372 5797 14381 5831
rect 14381 5797 14415 5831
rect 14415 5797 14424 5831
rect 14372 5788 14424 5797
rect 14648 5788 14700 5840
rect 23112 5788 23164 5840
rect 12624 5720 12676 5772
rect 14188 5720 14240 5772
rect 11796 5652 11848 5704
rect 12808 5652 12860 5704
rect 14280 5695 14332 5704
rect 10876 5516 10928 5568
rect 11244 5584 11296 5636
rect 12348 5584 12400 5636
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 16120 5652 16172 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17868 5720 17920 5772
rect 19800 5720 19852 5772
rect 19892 5720 19944 5772
rect 21180 5720 21232 5772
rect 21916 5720 21968 5772
rect 11612 5516 11664 5568
rect 11888 5516 11940 5568
rect 12624 5516 12676 5568
rect 14004 5584 14056 5636
rect 15016 5627 15068 5636
rect 15016 5593 15025 5627
rect 15025 5593 15059 5627
rect 15059 5593 15068 5627
rect 15016 5584 15068 5593
rect 15108 5627 15160 5636
rect 15108 5593 15117 5627
rect 15117 5593 15151 5627
rect 15151 5593 15160 5627
rect 15108 5584 15160 5593
rect 15844 5584 15896 5636
rect 17868 5584 17920 5636
rect 18236 5652 18288 5704
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 18788 5652 18840 5704
rect 20076 5652 20128 5704
rect 20812 5695 20864 5704
rect 20812 5661 20821 5695
rect 20821 5661 20855 5695
rect 20855 5661 20864 5695
rect 20812 5652 20864 5661
rect 20996 5652 21048 5704
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 37740 5652 37792 5704
rect 16856 5516 16908 5568
rect 20076 5516 20128 5568
rect 22008 5559 22060 5568
rect 22008 5525 22017 5559
rect 22017 5525 22051 5559
rect 22051 5525 22060 5559
rect 22008 5516 22060 5525
rect 23388 5559 23440 5568
rect 23388 5525 23397 5559
rect 23397 5525 23431 5559
rect 23431 5525 23440 5559
rect 23388 5516 23440 5525
rect 37556 5516 37608 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 2228 5244 2280 5296
rect 5908 5312 5960 5364
rect 6552 5312 6604 5364
rect 6092 5244 6144 5296
rect 6276 5244 6328 5296
rect 6460 5244 6512 5296
rect 6920 5312 6972 5364
rect 7104 5312 7156 5364
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 9404 5312 9456 5364
rect 9588 5312 9640 5364
rect 10048 5312 10100 5364
rect 11060 5355 11112 5364
rect 1584 5176 1636 5228
rect 8484 5176 8536 5228
rect 9220 5176 9272 5228
rect 2872 5108 2924 5160
rect 4068 5108 4120 5160
rect 4160 5108 4212 5160
rect 3884 4972 3936 5024
rect 4988 5108 5040 5160
rect 6541 5151 6593 5160
rect 6541 5117 6561 5151
rect 6561 5117 6593 5151
rect 6541 5108 6593 5117
rect 6920 5108 6972 5160
rect 9588 5176 9640 5228
rect 9956 5244 10008 5296
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11796 5312 11848 5364
rect 11888 5312 11940 5364
rect 10048 5176 10100 5228
rect 10692 5176 10744 5228
rect 10784 5176 10836 5228
rect 12532 5312 12584 5364
rect 13176 5244 13228 5296
rect 4620 4972 4672 5024
rect 4988 4972 5040 5024
rect 6368 5040 6420 5092
rect 5724 4972 5776 5024
rect 11244 5040 11296 5092
rect 8392 4972 8444 5024
rect 9680 4972 9732 5024
rect 10692 4972 10744 5024
rect 12624 5108 12676 5160
rect 14096 5312 14148 5364
rect 14372 5312 14424 5364
rect 15200 5312 15252 5364
rect 14464 5244 14516 5296
rect 15752 5312 15804 5364
rect 16488 5312 16540 5364
rect 17408 5312 17460 5364
rect 18144 5312 18196 5364
rect 14280 5176 14332 5228
rect 15752 5176 15804 5228
rect 16120 5219 16172 5228
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 16304 5176 16356 5228
rect 17776 5176 17828 5228
rect 18144 5219 18196 5228
rect 18144 5185 18153 5219
rect 18153 5185 18187 5219
rect 18187 5185 18196 5219
rect 19156 5244 19208 5296
rect 24124 5312 24176 5364
rect 18144 5176 18196 5185
rect 13176 5108 13228 5160
rect 11612 5040 11664 5092
rect 11704 4972 11756 5024
rect 12164 4972 12216 5024
rect 13452 4972 13504 5024
rect 17500 5151 17552 5160
rect 17500 5117 17509 5151
rect 17509 5117 17543 5151
rect 17543 5117 17552 5151
rect 17500 5108 17552 5117
rect 18604 5108 18656 5160
rect 20260 5176 20312 5228
rect 21824 5219 21876 5228
rect 17868 5040 17920 5092
rect 18236 5040 18288 5092
rect 13912 4972 13964 5024
rect 19432 5108 19484 5160
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 22284 5176 22336 5228
rect 22928 5176 22980 5228
rect 32404 5176 32456 5228
rect 20812 5108 20864 5160
rect 18788 5040 18840 5092
rect 19248 5040 19300 5092
rect 18972 4972 19024 5024
rect 20536 5040 20588 5092
rect 19524 4972 19576 5024
rect 19984 4972 20036 5024
rect 20444 4972 20496 5024
rect 22284 5015 22336 5024
rect 22284 4981 22293 5015
rect 22293 4981 22327 5015
rect 22327 4981 22336 5015
rect 22284 4972 22336 4981
rect 38200 5015 38252 5024
rect 38200 4981 38209 5015
rect 38209 4981 38243 5015
rect 38243 4981 38252 5015
rect 38200 4972 38252 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2504 4768 2556 4820
rect 3332 4700 3384 4752
rect 3792 4700 3844 4752
rect 7288 4743 7340 4752
rect 7288 4709 7297 4743
rect 7297 4709 7331 4743
rect 7331 4709 7340 4743
rect 7288 4700 7340 4709
rect 7656 4768 7708 4820
rect 8208 4768 8260 4820
rect 8300 4700 8352 4752
rect 8760 4768 8812 4820
rect 8944 4768 8996 4820
rect 9404 4768 9456 4820
rect 10600 4768 10652 4820
rect 1584 4632 1636 4684
rect 2044 4632 2096 4684
rect 2964 4632 3016 4684
rect 10968 4700 11020 4752
rect 4436 4564 4488 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5356 4564 5408 4616
rect 7196 4564 7248 4616
rect 7656 4564 7708 4616
rect 8208 4564 8260 4616
rect 8944 4564 8996 4616
rect 9956 4564 10008 4616
rect 10692 4632 10744 4684
rect 11520 4768 11572 4820
rect 11796 4768 11848 4820
rect 12440 4768 12492 4820
rect 12808 4768 12860 4820
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 11428 4700 11480 4752
rect 10876 4564 10928 4616
rect 11796 4564 11848 4616
rect 12256 4607 12308 4616
rect 12256 4573 12265 4607
rect 12265 4573 12299 4607
rect 12299 4573 12308 4607
rect 12256 4564 12308 4573
rect 5724 4496 5776 4548
rect 3976 4471 4028 4480
rect 3976 4437 3985 4471
rect 3985 4437 4019 4471
rect 4019 4437 4028 4471
rect 3976 4428 4028 4437
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 4804 4428 4856 4480
rect 9680 4496 9732 4548
rect 9772 4496 9824 4548
rect 8392 4428 8444 4480
rect 8944 4428 8996 4480
rect 11612 4428 11664 4480
rect 12072 4496 12124 4548
rect 12532 4564 12584 4616
rect 12992 4564 13044 4616
rect 12716 4496 12768 4548
rect 13176 4632 13228 4684
rect 13452 4632 13504 4684
rect 14464 4700 14516 4752
rect 14188 4632 14240 4684
rect 14648 4632 14700 4684
rect 13912 4564 13964 4616
rect 14004 4564 14056 4616
rect 16488 4768 16540 4820
rect 16672 4768 16724 4820
rect 15016 4700 15068 4752
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 15016 4564 15068 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 13176 4496 13228 4548
rect 13728 4496 13780 4548
rect 16764 4700 16816 4752
rect 17040 4700 17092 4752
rect 17408 4700 17460 4752
rect 17776 4700 17828 4752
rect 16672 4632 16724 4684
rect 22100 4811 22152 4820
rect 22100 4777 22109 4811
rect 22109 4777 22143 4811
rect 22143 4777 22152 4811
rect 22100 4768 22152 4777
rect 22376 4700 22428 4752
rect 16396 4564 16448 4616
rect 17776 4607 17828 4616
rect 17776 4573 17785 4607
rect 17785 4573 17819 4607
rect 17819 4573 17828 4607
rect 17776 4564 17828 4573
rect 18328 4564 18380 4616
rect 19340 4564 19392 4616
rect 19616 4564 19668 4616
rect 19524 4539 19576 4548
rect 19524 4505 19533 4539
rect 19533 4505 19567 4539
rect 19567 4505 19576 4539
rect 19524 4496 19576 4505
rect 20168 4539 20220 4548
rect 20168 4505 20177 4539
rect 20177 4505 20211 4539
rect 20211 4505 20220 4539
rect 20168 4496 20220 4505
rect 20812 4564 20864 4616
rect 21180 4564 21232 4616
rect 21824 4564 21876 4616
rect 23480 4632 23532 4684
rect 31300 4607 31352 4616
rect 21088 4496 21140 4548
rect 21364 4496 21416 4548
rect 31300 4573 31309 4607
rect 31309 4573 31343 4607
rect 31343 4573 31352 4607
rect 31300 4564 31352 4573
rect 15200 4428 15252 4480
rect 15752 4428 15804 4480
rect 17500 4428 17552 4480
rect 17592 4428 17644 4480
rect 19432 4428 19484 4480
rect 19984 4428 20036 4480
rect 20628 4428 20680 4480
rect 20720 4428 20772 4480
rect 24124 4428 24176 4480
rect 38200 4471 38252 4480
rect 38200 4437 38209 4471
rect 38209 4437 38243 4471
rect 38243 4437 38252 4471
rect 38200 4428 38252 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2780 4224 2832 4276
rect 3148 4224 3200 4276
rect 3884 4224 3936 4276
rect 1676 4199 1728 4208
rect 1676 4165 1685 4199
rect 1685 4165 1719 4199
rect 1719 4165 1728 4199
rect 1676 4156 1728 4165
rect 3240 4156 3292 4208
rect 3700 4156 3752 4208
rect 8208 4156 8260 4208
rect 9312 4224 9364 4276
rect 9588 4224 9640 4276
rect 8944 4156 8996 4208
rect 9956 4156 10008 4208
rect 848 4088 900 4140
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 10508 4088 10560 4140
rect 11428 4156 11480 4208
rect 12164 4224 12216 4276
rect 14372 4224 14424 4276
rect 14648 4224 14700 4276
rect 17040 4224 17092 4276
rect 17224 4224 17276 4276
rect 12532 4156 12584 4208
rect 12716 4156 12768 4208
rect 17776 4156 17828 4208
rect 18236 4156 18288 4208
rect 19432 4224 19484 4276
rect 31300 4224 31352 4276
rect 11980 4088 12032 4140
rect 12440 4088 12492 4140
rect 12808 4088 12860 4140
rect 13360 4088 13412 4140
rect 13728 4088 13780 4140
rect 13912 4088 13964 4140
rect 14096 4088 14148 4140
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14464 4088 14516 4140
rect 2964 3952 3016 4004
rect 15108 4020 15160 4072
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 15844 4088 15896 4140
rect 16672 4088 16724 4140
rect 17500 4131 17552 4140
rect 17500 4097 17509 4131
rect 17509 4097 17543 4131
rect 17543 4097 17552 4131
rect 17500 4088 17552 4097
rect 17868 4088 17920 4140
rect 18420 4088 18472 4140
rect 20720 4156 20772 4208
rect 23112 4156 23164 4208
rect 19432 4131 19484 4140
rect 19432 4097 19441 4131
rect 19441 4097 19475 4131
rect 19475 4097 19484 4131
rect 19432 4088 19484 4097
rect 19524 4131 19576 4140
rect 19524 4097 19533 4131
rect 19533 4097 19567 4131
rect 19567 4097 19576 4131
rect 19524 4088 19576 4097
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 21456 4088 21508 4140
rect 22468 4088 22520 4140
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 38016 4131 38068 4140
rect 38016 4097 38025 4131
rect 38025 4097 38059 4131
rect 38059 4097 38068 4131
rect 38016 4088 38068 4097
rect 5172 3952 5224 4004
rect 6460 3952 6512 4004
rect 8852 3952 8904 4004
rect 3700 3884 3752 3936
rect 5356 3884 5408 3936
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 10140 3952 10192 4004
rect 12072 3952 12124 4004
rect 12348 3995 12400 4004
rect 12348 3961 12357 3995
rect 12357 3961 12391 3995
rect 12391 3961 12400 3995
rect 12348 3952 12400 3961
rect 12992 3952 13044 4004
rect 14464 3952 14516 4004
rect 14556 3952 14608 4004
rect 15200 3952 15252 4004
rect 9220 3884 9272 3936
rect 9404 3884 9456 3936
rect 10232 3884 10284 3936
rect 10324 3884 10376 3936
rect 12164 3884 12216 3936
rect 12440 3884 12492 3936
rect 13084 3884 13136 3936
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 13728 3884 13780 3936
rect 14740 3884 14792 3936
rect 15108 3884 15160 3936
rect 15568 3952 15620 4004
rect 17316 3952 17368 4004
rect 17684 3952 17736 4004
rect 15936 3884 15988 3936
rect 17776 3884 17828 3936
rect 18144 3884 18196 3936
rect 18328 3884 18380 3936
rect 18420 3884 18472 3936
rect 19984 3952 20036 4004
rect 19156 3884 19208 3936
rect 23020 3952 23072 4004
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 20996 3884 21048 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 37188 3884 37240 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3976 3680 4028 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 9496 3680 9548 3732
rect 10600 3680 10652 3732
rect 12164 3680 12216 3732
rect 9680 3612 9732 3664
rect 11336 3612 11388 3664
rect 11796 3612 11848 3664
rect 12624 3680 12676 3732
rect 12992 3680 13044 3732
rect 13176 3680 13228 3732
rect 16580 3680 16632 3732
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 18512 3680 18564 3732
rect 19156 3680 19208 3732
rect 19892 3680 19944 3732
rect 14188 3612 14240 3664
rect 18236 3612 18288 3664
rect 1584 3544 1636 3596
rect 3516 3544 3568 3596
rect 4620 3544 4672 3596
rect 4712 3544 4764 3596
rect 7196 3544 7248 3596
rect 9404 3544 9456 3596
rect 10784 3544 10836 3596
rect 4160 3476 4212 3528
rect 6000 3476 6052 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 8300 3476 8352 3528
rect 9128 3476 9180 3528
rect 10232 3476 10284 3528
rect 664 3340 716 3392
rect 3332 3340 3384 3392
rect 4712 3408 4764 3460
rect 7380 3340 7432 3392
rect 9772 3408 9824 3460
rect 10048 3408 10100 3460
rect 10508 3476 10560 3528
rect 11888 3476 11940 3528
rect 12624 3544 12676 3596
rect 16856 3544 16908 3596
rect 16948 3544 17000 3596
rect 17776 3544 17828 3596
rect 20628 3680 20680 3732
rect 24584 3723 24636 3732
rect 24584 3689 24593 3723
rect 24593 3689 24627 3723
rect 24627 3689 24636 3723
rect 24584 3680 24636 3689
rect 35808 3680 35860 3732
rect 21916 3612 21968 3664
rect 10600 3408 10652 3460
rect 10876 3408 10928 3460
rect 12440 3408 12492 3460
rect 12992 3476 13044 3528
rect 13084 3476 13136 3528
rect 14464 3476 14516 3528
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15200 3476 15252 3528
rect 15476 3476 15528 3528
rect 16580 3476 16632 3528
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 18052 3476 18104 3528
rect 18420 3476 18472 3528
rect 22192 3544 22244 3596
rect 35716 3612 35768 3664
rect 19248 3476 19300 3528
rect 7748 3340 7800 3392
rect 12624 3340 12676 3392
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 15660 3408 15712 3460
rect 16856 3408 16908 3460
rect 20628 3476 20680 3528
rect 21180 3476 21232 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 22008 3519 22060 3528
rect 22008 3485 22017 3519
rect 22017 3485 22051 3519
rect 22051 3485 22060 3519
rect 22008 3476 22060 3485
rect 22284 3476 22336 3528
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 21088 3408 21140 3460
rect 37280 3476 37332 3528
rect 39304 3476 39356 3528
rect 38292 3408 38344 3460
rect 16580 3340 16632 3392
rect 17316 3340 17368 3392
rect 19248 3340 19300 3392
rect 19984 3340 20036 3392
rect 21456 3383 21508 3392
rect 21456 3349 21465 3383
rect 21465 3349 21499 3383
rect 21499 3349 21508 3383
rect 21456 3340 21508 3349
rect 21548 3340 21600 3392
rect 22284 3383 22336 3392
rect 22284 3349 22293 3383
rect 22293 3349 22327 3383
rect 22327 3349 22336 3383
rect 22284 3340 22336 3349
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 23940 3340 23992 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3148 3136 3200 3188
rect 3516 3136 3568 3188
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 2964 3000 3016 3052
rect 2596 2932 2648 2984
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 8208 3068 8260 3120
rect 11152 3136 11204 3188
rect 10692 3111 10744 3120
rect 10692 3077 10701 3111
rect 10701 3077 10735 3111
rect 10735 3077 10744 3111
rect 10692 3068 10744 3077
rect 3700 3000 3752 3052
rect 5356 3000 5408 3052
rect 6552 3043 6604 3052
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 4160 2932 4212 2984
rect 5908 2932 5960 2984
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 9404 3000 9456 3052
rect 9680 3000 9732 3052
rect 10324 3000 10376 3052
rect 1308 2796 1360 2848
rect 11152 2932 11204 2984
rect 12716 3136 12768 3188
rect 12900 3179 12952 3188
rect 12900 3145 12909 3179
rect 12909 3145 12943 3179
rect 12943 3145 12952 3179
rect 12900 3136 12952 3145
rect 13544 3179 13596 3188
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13544 3136 13596 3145
rect 13636 3136 13688 3188
rect 14740 3136 14792 3188
rect 15384 3136 15436 3188
rect 19524 3136 19576 3188
rect 20168 3136 20220 3188
rect 21548 3136 21600 3188
rect 22836 3136 22888 3188
rect 23296 3136 23348 3188
rect 25872 3136 25924 3188
rect 30380 3136 30432 3188
rect 34428 3136 34480 3188
rect 18236 3068 18288 3120
rect 11428 2932 11480 2984
rect 12348 3000 12400 3052
rect 12440 3000 12492 3052
rect 13360 3000 13412 3052
rect 13636 3000 13688 3052
rect 13728 3000 13780 3052
rect 14556 3000 14608 3052
rect 14740 3043 14792 3052
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 15844 3000 15896 3052
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 18052 3000 18104 3052
rect 18328 3043 18380 3052
rect 18328 3009 18337 3043
rect 18337 3009 18371 3043
rect 18371 3009 18380 3043
rect 18328 3000 18380 3009
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 19156 3000 19208 3052
rect 19984 3000 20036 3052
rect 20996 3043 21048 3052
rect 20996 3009 21005 3043
rect 21005 3009 21039 3043
rect 21039 3009 21048 3043
rect 20996 3000 21048 3009
rect 12624 2932 12676 2984
rect 21456 3068 21508 3120
rect 21916 3000 21968 3052
rect 28816 3068 28868 3120
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 26608 3043 26660 3052
rect 26608 3009 26617 3043
rect 26617 3009 26651 3043
rect 26651 3009 26660 3043
rect 26608 3000 26660 3009
rect 27712 3000 27764 3052
rect 32864 3000 32916 3052
rect 36912 3043 36964 3052
rect 36912 3009 36921 3043
rect 36921 3009 36955 3043
rect 36955 3009 36964 3043
rect 36912 3000 36964 3009
rect 37556 3000 37608 3052
rect 5540 2839 5592 2848
rect 5540 2805 5549 2839
rect 5549 2805 5583 2839
rect 5583 2805 5592 2839
rect 5540 2796 5592 2805
rect 8208 2839 8260 2848
rect 8208 2805 8217 2839
rect 8217 2805 8251 2839
rect 8251 2805 8260 2839
rect 8208 2796 8260 2805
rect 8392 2796 8444 2848
rect 11704 2864 11756 2916
rect 12716 2864 12768 2916
rect 16856 2864 16908 2916
rect 11612 2796 11664 2848
rect 11980 2796 12032 2848
rect 13636 2796 13688 2848
rect 13820 2796 13872 2848
rect 16764 2796 16816 2848
rect 17500 2796 17552 2848
rect 20904 2864 20956 2916
rect 22192 2864 22244 2916
rect 23204 2864 23256 2916
rect 28908 2864 28960 2916
rect 19064 2796 19116 2848
rect 23296 2839 23348 2848
rect 23296 2805 23305 2839
rect 23305 2805 23339 2839
rect 23339 2805 23348 2839
rect 23296 2796 23348 2805
rect 23848 2796 23900 2848
rect 25044 2839 25096 2848
rect 25044 2805 25053 2839
rect 25053 2805 25087 2839
rect 25087 2805 25096 2839
rect 25044 2796 25096 2805
rect 38016 2796 38068 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3148 2592 3200 2644
rect 4068 2592 4120 2644
rect 5724 2592 5776 2644
rect 4620 2567 4672 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 4620 2533 4629 2567
rect 4629 2533 4663 2567
rect 4663 2533 4672 2567
rect 4620 2524 4672 2533
rect 5264 2567 5316 2576
rect 5264 2533 5273 2567
rect 5273 2533 5307 2567
rect 5307 2533 5316 2567
rect 5264 2524 5316 2533
rect 5080 2363 5132 2372
rect 5080 2329 5089 2363
rect 5089 2329 5123 2363
rect 5123 2329 5132 2363
rect 5080 2320 5132 2329
rect 10876 2524 10928 2576
rect 10968 2456 11020 2508
rect 11796 2456 11848 2508
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 9680 2388 9732 2440
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 12716 2592 12768 2644
rect 12440 2524 12492 2576
rect 13728 2524 13780 2576
rect 12532 2456 12584 2508
rect 14464 2592 14516 2644
rect 19156 2592 19208 2644
rect 19248 2592 19300 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 26148 2592 26200 2644
rect 12440 2388 12492 2440
rect 12624 2388 12676 2440
rect 12808 2388 12860 2440
rect 18880 2524 18932 2576
rect 21088 2524 21140 2576
rect 24860 2524 24912 2576
rect 25136 2524 25188 2576
rect 19340 2456 19392 2508
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 22192 2456 22244 2508
rect 14832 2388 14884 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16856 2320 16908 2372
rect 17408 2388 17460 2440
rect 18696 2388 18748 2440
rect 19984 2388 20036 2440
rect 21548 2388 21600 2440
rect 23296 2431 23348 2440
rect 20444 2320 20496 2372
rect 21272 2320 21324 2372
rect 23296 2397 23305 2431
rect 23305 2397 23339 2431
rect 23339 2397 23348 2431
rect 23296 2388 23348 2397
rect 24492 2388 24544 2440
rect 24768 2456 24820 2508
rect 25780 2388 25832 2440
rect 34796 2592 34848 2644
rect 30196 2456 30248 2508
rect 28448 2431 28500 2440
rect 28448 2397 28457 2431
rect 28457 2397 28491 2431
rect 28491 2397 28500 2431
rect 29920 2431 29972 2440
rect 28448 2388 28500 2397
rect 29920 2397 29929 2431
rect 29929 2397 29963 2431
rect 29963 2397 29972 2431
rect 29920 2388 29972 2397
rect 33600 2431 33652 2440
rect 26424 2320 26476 2372
rect 28908 2320 28960 2372
rect 33600 2397 33609 2431
rect 33609 2397 33643 2431
rect 33643 2397 33652 2431
rect 33600 2388 33652 2397
rect 37648 2456 37700 2508
rect 37372 2388 37424 2440
rect 37740 2431 37792 2440
rect 37740 2397 37749 2431
rect 37749 2397 37783 2431
rect 37783 2397 37792 2431
rect 37740 2388 37792 2397
rect 34796 2320 34848 2372
rect 35440 2320 35492 2372
rect 3884 2252 3936 2304
rect 5816 2252 5868 2304
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 7104 2252 7156 2304
rect 8116 2295 8168 2304
rect 8116 2261 8125 2295
rect 8125 2261 8159 2295
rect 8159 2261 8168 2295
rect 8116 2252 8168 2261
rect 11152 2252 11204 2304
rect 12164 2252 12216 2304
rect 12256 2252 12308 2304
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 14372 2295 14424 2304
rect 14372 2261 14381 2295
rect 14381 2261 14415 2295
rect 14415 2261 14424 2295
rect 14372 2252 14424 2261
rect 14464 2252 14516 2304
rect 20812 2252 20864 2304
rect 23204 2252 23256 2304
rect 28356 2252 28408 2304
rect 29736 2295 29788 2304
rect 29736 2261 29745 2295
rect 29745 2261 29779 2295
rect 29779 2261 29788 2295
rect 29736 2252 29788 2261
rect 30380 2295 30432 2304
rect 30380 2261 30389 2295
rect 30389 2261 30423 2295
rect 30423 2261 30432 2295
rect 30380 2252 30432 2261
rect 30932 2252 30984 2304
rect 32220 2252 32272 2304
rect 33508 2252 33560 2304
rect 36728 2252 36780 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 6276 2048 6328 2100
rect 9956 2048 10008 2100
rect 10048 2048 10100 2100
rect 3424 1980 3476 2032
rect 12532 1980 12584 2032
rect 12716 2048 12768 2100
rect 20168 2048 20220 2100
rect 28448 2048 28500 2100
rect 30748 2048 30800 2100
rect 17776 1980 17828 2032
rect 19064 1980 19116 2032
rect 20076 1980 20128 2032
rect 28816 1980 28868 2032
rect 37740 1980 37792 2032
rect 3332 1912 3384 1964
rect 5356 1912 5408 1964
rect 17224 1912 17276 1964
rect 9128 1844 9180 1896
rect 22652 1844 22704 1896
rect 6000 1776 6052 1828
rect 22744 1776 22796 1828
rect 6644 1708 6696 1760
rect 22100 1708 22152 1760
rect 6552 1640 6604 1692
rect 9956 1640 10008 1692
rect 17132 1640 17184 1692
rect 13268 1572 13320 1624
rect 17224 1572 17276 1624
rect 23756 1572 23808 1624
rect 7564 1504 7616 1556
rect 13636 1504 13688 1556
rect 8024 1436 8076 1488
rect 15568 1504 15620 1556
rect 15200 1436 15252 1488
rect 26608 1436 26660 1488
rect 5908 1368 5960 1420
rect 14372 1368 14424 1420
rect 29000 1368 29052 1420
rect 29920 1368 29972 1420
rect 20 1300 72 1352
rect 8208 1300 8260 1352
rect 9036 1300 9088 1352
rect 20720 1300 20772 1352
rect 5540 1232 5592 1284
rect 17960 1232 18012 1284
rect 12900 1164 12952 1216
rect 17316 1164 17368 1216
rect 3516 756 3568 808
rect 8116 756 8168 808
<< metal2 >>
rect 18 39200 74 39800
rect 1306 39200 1362 39800
rect 1950 39200 2006 39800
rect 2594 39200 2650 39800
rect 3054 39536 3110 39545
rect 3054 39471 3110 39480
rect 32 36242 60 39200
rect 1320 36922 1348 39200
rect 1964 37262 1992 39200
rect 1952 37256 2004 37262
rect 2608 37244 2636 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 2884 37330 2912 38791
rect 2872 37324 2924 37330
rect 2872 37266 2924 37272
rect 2964 37256 3016 37262
rect 2608 37216 2820 37244
rect 1952 37198 2004 37204
rect 2792 37126 2820 37216
rect 2964 37198 3016 37204
rect 2780 37120 2832 37126
rect 2780 37062 2832 37068
rect 1308 36916 1360 36922
rect 1308 36858 1360 36864
rect 1766 36816 1822 36825
rect 1766 36751 1822 36760
rect 2320 36780 2372 36786
rect 1780 36378 1808 36751
rect 2320 36722 2372 36728
rect 2332 36378 2360 36722
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 2320 36372 2372 36378
rect 2320 36314 2372 36320
rect 20 36236 72 36242
rect 20 36178 72 36184
rect 2872 36100 2924 36106
rect 2872 36042 2924 36048
rect 1584 35624 1636 35630
rect 1584 35566 1636 35572
rect 2136 35624 2188 35630
rect 2136 35566 2188 35572
rect 1596 35465 1624 35566
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1780 34105 1808 34546
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 112 33516 164 33522
rect 112 33458 164 33464
rect 20 33448 72 33454
rect 20 33390 72 33396
rect 32 19825 60 33390
rect 124 23497 152 33458
rect 1124 33040 1176 33046
rect 1124 32982 1176 32988
rect 848 31816 900 31822
rect 848 31758 900 31764
rect 756 31408 808 31414
rect 756 31350 808 31356
rect 664 30728 716 30734
rect 664 30670 716 30676
rect 572 29300 624 29306
rect 572 29242 624 29248
rect 110 23488 166 23497
rect 110 23423 166 23432
rect 18 19816 74 19825
rect 18 19751 74 19760
rect 584 17270 612 29242
rect 572 17264 624 17270
rect 572 17206 624 17212
rect 676 15094 704 30670
rect 664 15088 716 15094
rect 664 15030 716 15036
rect 768 11898 796 31350
rect 756 11892 808 11898
rect 756 11834 808 11840
rect 860 4146 888 31758
rect 1032 31136 1084 31142
rect 1032 31078 1084 31084
rect 940 27056 992 27062
rect 940 26998 992 27004
rect 952 15706 980 26998
rect 1044 17542 1072 31078
rect 1136 21146 1164 32982
rect 1492 32972 1544 32978
rect 1492 32914 1544 32920
rect 1400 31340 1452 31346
rect 1400 31282 1452 31288
rect 1216 30796 1268 30802
rect 1216 30738 1268 30744
rect 1124 21140 1176 21146
rect 1124 21082 1176 21088
rect 1228 20602 1256 30738
rect 1412 30433 1440 31282
rect 1398 30424 1454 30433
rect 1398 30359 1454 30368
rect 1308 29028 1360 29034
rect 1308 28970 1360 28976
rect 1320 22710 1348 28970
rect 1504 25498 1532 32914
rect 1768 32768 1820 32774
rect 1766 32736 1768 32745
rect 1820 32736 1822 32745
rect 1766 32671 1822 32680
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1952 32224 2004 32230
rect 1952 32166 2004 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1860 31204 1912 31210
rect 1860 31146 1912 31152
rect 1766 30696 1822 30705
rect 1766 30631 1822 30640
rect 1780 30122 1808 30631
rect 1768 30116 1820 30122
rect 1768 30058 1820 30064
rect 1676 30048 1728 30054
rect 1676 29990 1728 29996
rect 1584 28960 1636 28966
rect 1584 28902 1636 28908
rect 1596 28082 1624 28902
rect 1584 28076 1636 28082
rect 1584 28018 1636 28024
rect 1584 26920 1636 26926
rect 1584 26862 1636 26868
rect 1492 25492 1544 25498
rect 1492 25434 1544 25440
rect 1596 24138 1624 26862
rect 1688 25106 1716 29990
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1780 29345 1808 29446
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1766 27976 1822 27985
rect 1766 27911 1768 27920
rect 1820 27911 1822 27920
rect 1768 27882 1820 27888
rect 1768 27328 1820 27334
rect 1766 27296 1768 27305
rect 1820 27296 1822 27305
rect 1766 27231 1822 27240
rect 1768 26240 1820 26246
rect 1768 26182 1820 26188
rect 1780 25265 1808 26182
rect 1766 25256 1822 25265
rect 1766 25191 1822 25200
rect 1688 25078 1808 25106
rect 1780 24886 1808 25078
rect 1768 24880 1820 24886
rect 1768 24822 1820 24828
rect 1872 24750 1900 31146
rect 1964 28558 1992 32166
rect 2148 30666 2176 35566
rect 2884 33114 2912 36042
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2228 32768 2280 32774
rect 2228 32710 2280 32716
rect 2240 32570 2268 32710
rect 2228 32564 2280 32570
rect 2228 32506 2280 32512
rect 2700 32230 2728 32846
rect 2688 32224 2740 32230
rect 2688 32166 2740 32172
rect 2976 32026 3004 37198
rect 3068 36786 3096 39471
rect 3882 39200 3938 39800
rect 4526 39200 4582 39800
rect 5814 39200 5870 39800
rect 6458 39200 6514 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 10966 39200 11022 39800
rect 11610 39200 11666 39800
rect 12898 39200 12954 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 15474 39200 15530 39800
rect 16118 39200 16174 39800
rect 16224 39222 16528 39250
rect 3146 37496 3202 37505
rect 3146 37431 3202 37440
rect 3160 36854 3188 37431
rect 3896 36854 3924 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37126 4660 37726
rect 5828 37262 5856 39200
rect 5724 37256 5776 37262
rect 5724 37198 5776 37204
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 3148 36848 3200 36854
rect 3148 36790 3200 36796
rect 3884 36848 3936 36854
rect 3884 36790 3936 36796
rect 3056 36780 3108 36786
rect 3056 36722 3108 36728
rect 5356 36644 5408 36650
rect 5356 36586 5408 36592
rect 3148 36576 3200 36582
rect 3148 36518 3200 36524
rect 3160 36242 3188 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3148 36236 3200 36242
rect 3148 36178 3200 36184
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 4080 34610 4108 35974
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34604 4120 34610
rect 4068 34546 4120 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 3424 33380 3476 33386
rect 3424 33322 3476 33328
rect 3056 32428 3108 32434
rect 3056 32370 3108 32376
rect 2964 32020 3016 32026
rect 2964 31962 3016 31968
rect 2136 30660 2188 30666
rect 2136 30602 2188 30608
rect 2044 30592 2096 30598
rect 2044 30534 2096 30540
rect 2056 30433 2084 30534
rect 2042 30424 2098 30433
rect 2042 30359 2098 30368
rect 2148 29238 2176 30602
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2596 29640 2648 29646
rect 2596 29582 2648 29588
rect 2136 29232 2188 29238
rect 2136 29174 2188 29180
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 1952 28552 2004 28558
rect 1952 28494 2004 28500
rect 2228 28416 2280 28422
rect 2228 28358 2280 28364
rect 2136 26988 2188 26994
rect 2136 26930 2188 26936
rect 2044 26784 2096 26790
rect 2044 26726 2096 26732
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1964 24954 1992 25230
rect 2056 25129 2084 26726
rect 2042 25120 2098 25129
rect 2042 25055 2098 25064
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 1860 24744 1912 24750
rect 1860 24686 1912 24692
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 1584 24132 1636 24138
rect 1584 24074 1636 24080
rect 1872 23662 1900 24210
rect 2148 24154 2176 26930
rect 2240 26042 2268 28358
rect 2424 27418 2452 29106
rect 2608 29073 2636 29582
rect 2594 29064 2650 29073
rect 2594 28999 2650 29008
rect 2596 28688 2648 28694
rect 2596 28630 2648 28636
rect 2424 27390 2544 27418
rect 2412 27328 2464 27334
rect 2412 27270 2464 27276
rect 2228 26036 2280 26042
rect 2228 25978 2280 25984
rect 2320 25968 2372 25974
rect 2318 25936 2320 25945
rect 2372 25936 2374 25945
rect 2318 25871 2374 25880
rect 2228 25832 2280 25838
rect 2228 25774 2280 25780
rect 1964 24126 2176 24154
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1872 23186 1900 23598
rect 1964 23186 1992 24126
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 2136 24064 2188 24070
rect 2136 24006 2188 24012
rect 1860 23180 1912 23186
rect 1860 23122 1912 23128
rect 1952 23180 2004 23186
rect 1952 23122 2004 23128
rect 1490 23080 1546 23089
rect 1490 23015 1546 23024
rect 1768 23044 1820 23050
rect 1308 22704 1360 22710
rect 1308 22646 1360 22652
rect 1216 20596 1268 20602
rect 1216 20538 1268 20544
rect 1032 17536 1084 17542
rect 1032 17478 1084 17484
rect 1504 17218 1532 23015
rect 1768 22986 1820 22992
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1688 22574 1716 22714
rect 1676 22568 1728 22574
rect 1582 22536 1638 22545
rect 1676 22510 1728 22516
rect 1582 22471 1638 22480
rect 1596 21554 1624 22471
rect 1688 22098 1716 22510
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1584 21548 1636 21554
rect 1584 21490 1636 21496
rect 1780 20262 1808 22986
rect 1872 21622 1900 23122
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 1964 22098 1992 22374
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 1860 21616 1912 21622
rect 1860 21558 1912 21564
rect 1950 21584 2006 21593
rect 1872 21010 1900 21558
rect 1950 21519 2006 21528
rect 1964 21486 1992 21519
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 1872 20466 1900 20946
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1872 19922 1900 20402
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1768 19372 1820 19378
rect 1872 19360 1900 19858
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1820 19332 1900 19360
rect 1768 19314 1820 19320
rect 1872 18834 1900 19332
rect 1860 18828 1912 18834
rect 1860 18770 1912 18776
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1766 18456 1822 18465
rect 1872 18426 1900 18634
rect 1766 18391 1822 18400
rect 1860 18420 1912 18426
rect 1780 17338 1808 18391
rect 1860 18362 1912 18368
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1504 17190 1900 17218
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 940 15700 992 15706
rect 940 15642 992 15648
rect 952 12918 980 15642
rect 1596 15570 1624 16594
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1688 15745 1716 16050
rect 1674 15736 1730 15745
rect 1674 15671 1730 15680
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1596 15026 1624 15506
rect 1584 15020 1636 15026
rect 1584 14962 1636 14968
rect 1596 14482 1624 14962
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1780 13818 1808 16390
rect 1872 13938 1900 17190
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1688 13790 1808 13818
rect 940 12912 992 12918
rect 940 12854 992 12860
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1596 11762 1624 12242
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 11218 1624 11698
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1596 10810 1624 11154
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1596 10674 1624 10746
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10130 1624 10610
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1400 9648 1452 9654
rect 1398 9616 1400 9625
rect 1452 9616 1454 9625
rect 1596 9586 1624 10066
rect 1398 9551 1454 9560
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1688 9178 1716 13790
rect 1768 13728 1820 13734
rect 1766 13696 1768 13705
rect 1820 13696 1822 13705
rect 1766 13631 1822 13640
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1872 9738 1900 12038
rect 1964 10742 1992 19450
rect 2056 18970 2084 24006
rect 2148 22574 2176 24006
rect 2240 23526 2268 25774
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2136 22568 2188 22574
rect 2136 22510 2188 22516
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2240 18358 2268 23258
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 2332 18222 2360 24822
rect 2424 23322 2452 27270
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2412 23180 2464 23186
rect 2412 23122 2464 23128
rect 2424 22234 2452 23122
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2516 22094 2544 27390
rect 2608 26994 2636 28630
rect 2700 28529 2728 30194
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2686 28520 2742 28529
rect 2686 28455 2742 28464
rect 2688 28416 2740 28422
rect 2688 28358 2740 28364
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2424 22066 2544 22094
rect 2424 21978 2452 22066
rect 2424 21950 2544 21978
rect 2410 21856 2466 21865
rect 2410 21791 2466 21800
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 17202 2360 17682
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 12850 2084 13330
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 12306 2084 12786
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1964 9874 1992 10678
rect 2148 10266 2176 15030
rect 2240 13161 2268 16934
rect 2332 16658 2360 17138
rect 2424 16998 2452 21791
rect 2516 21690 2544 21950
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2410 16688 2466 16697
rect 2320 16652 2372 16658
rect 2410 16623 2466 16632
rect 2320 16594 2372 16600
rect 2226 13152 2282 13161
rect 2226 13087 2282 13096
rect 2424 11830 2452 16623
rect 2516 16574 2544 21422
rect 2608 19786 2636 26726
rect 2596 19780 2648 19786
rect 2596 19722 2648 19728
rect 2700 19718 2728 28358
rect 2792 26314 2820 29038
rect 2884 28082 2912 29106
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2872 27396 2924 27402
rect 2872 27338 2924 27344
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2792 22658 2820 25978
rect 2884 23798 2912 27338
rect 2976 26450 3004 30534
rect 2964 26444 3016 26450
rect 2964 26386 3016 26392
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2976 25702 3004 26182
rect 3068 26081 3096 32370
rect 3436 30734 3464 33322
rect 3976 33312 4028 33318
rect 3976 33254 4028 33260
rect 3700 32428 3752 32434
rect 3700 32370 3752 32376
rect 3516 31340 3568 31346
rect 3516 31282 3568 31288
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3332 30048 3384 30054
rect 3332 29990 3384 29996
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3054 26072 3110 26081
rect 3054 26007 3110 26016
rect 2964 25696 3016 25702
rect 2964 25638 3016 25644
rect 3054 24848 3110 24857
rect 3054 24783 3110 24792
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 2872 23792 2924 23798
rect 2872 23734 2924 23740
rect 2792 22630 2912 22658
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2792 20806 2820 22510
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2884 19922 2912 22630
rect 2976 20058 3004 23802
rect 3068 22094 3096 24783
rect 3160 24138 3188 28970
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3344 27418 3372 29990
rect 3436 28082 3464 30670
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 3252 26994 3280 27406
rect 3344 27390 3464 27418
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3252 25378 3280 26930
rect 3344 26586 3372 27270
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3436 25974 3464 27390
rect 3424 25968 3476 25974
rect 3424 25910 3476 25916
rect 3332 25832 3384 25838
rect 3332 25774 3384 25780
rect 3344 25498 3372 25774
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3252 25350 3372 25378
rect 3240 25220 3292 25226
rect 3240 25162 3292 25168
rect 3252 24274 3280 25162
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3148 24132 3200 24138
rect 3148 24074 3200 24080
rect 3238 23760 3294 23769
rect 3238 23695 3294 23704
rect 3252 22506 3280 23695
rect 3344 22982 3372 25350
rect 3436 24886 3464 25910
rect 3424 24880 3476 24886
rect 3424 24822 3476 24828
rect 3424 24608 3476 24614
rect 3422 24576 3424 24585
rect 3476 24576 3478 24585
rect 3422 24511 3478 24520
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 3436 23662 3464 24210
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3240 22500 3292 22506
rect 3240 22442 3292 22448
rect 3068 22066 3280 22094
rect 3252 21978 3280 22066
rect 3160 21950 3280 21978
rect 3054 20904 3110 20913
rect 3054 20839 3110 20848
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2870 19408 2926 19417
rect 2870 19343 2926 19352
rect 2884 18698 2912 19343
rect 2872 18692 2924 18698
rect 2872 18634 2924 18640
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17338 2728 17478
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 3068 17218 3096 20839
rect 2884 17190 3096 17218
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2516 16546 2636 16574
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2516 13394 2544 13806
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2502 11928 2558 11937
rect 2502 11863 2558 11872
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1964 9846 2452 9874
rect 1872 9710 1992 9738
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8430 1624 8910
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 7886 1624 8366
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 7324 1624 7822
rect 1766 7576 1822 7585
rect 1766 7511 1768 7520
rect 1820 7511 1822 7520
rect 1768 7482 1820 7488
rect 1676 7336 1728 7342
rect 1596 7296 1676 7324
rect 1596 6866 1624 7296
rect 1676 7278 1728 7284
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 5778 1624 6802
rect 1872 6662 1900 8842
rect 1964 6914 1992 9710
rect 2136 9648 2188 9654
rect 2188 9596 2360 9602
rect 2136 9590 2360 9596
rect 2148 9574 2360 9590
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 1964 6886 2084 6914
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1596 5234 1624 5714
rect 1674 5536 1730 5545
rect 1674 5471 1730 5480
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1596 4690 1624 5170
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 1596 3602 1624 4626
rect 1688 4214 1716 5471
rect 2056 4690 2084 6886
rect 2240 5302 2268 9318
rect 2332 6497 2360 9574
rect 2318 6488 2374 6497
rect 2318 6423 2374 6432
rect 2320 6384 2372 6390
rect 2318 6352 2320 6361
rect 2372 6352 2374 6361
rect 2318 6287 2374 6296
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 2424 4321 2452 9846
rect 2516 9382 2544 11863
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2608 6914 2636 16546
rect 2700 16114 2728 16594
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 11778 2820 14214
rect 2884 12102 2912 17190
rect 3160 16402 3188 21950
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21690 3280 21830
rect 3344 21690 3372 22918
rect 3436 22094 3464 23598
rect 3528 22710 3556 31282
rect 3712 30025 3740 32370
rect 3792 31952 3844 31958
rect 3792 31894 3844 31900
rect 3698 30016 3754 30025
rect 3698 29951 3754 29960
rect 3804 29594 3832 31894
rect 3988 30258 4016 33254
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 5368 32502 5396 36586
rect 5540 36576 5592 36582
rect 5540 36518 5592 36524
rect 5552 36174 5580 36518
rect 5736 36378 5764 37198
rect 6472 36786 6500 39200
rect 7116 37262 7144 39200
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 6828 37188 6880 37194
rect 6828 37130 6880 37136
rect 6460 36780 6512 36786
rect 6460 36722 6512 36728
rect 5724 36372 5776 36378
rect 5724 36314 5776 36320
rect 5540 36168 5592 36174
rect 5540 36110 5592 36116
rect 5816 34740 5868 34746
rect 5816 34682 5868 34688
rect 5356 32496 5408 32502
rect 5356 32438 5408 32444
rect 4988 32360 5040 32366
rect 4988 32302 5040 32308
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5000 31482 5028 32302
rect 5632 31952 5684 31958
rect 5632 31894 5684 31900
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 5080 31748 5132 31754
rect 5080 31690 5132 31696
rect 4988 31476 5040 31482
rect 4988 31418 5040 31424
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4436 30592 4488 30598
rect 4436 30534 4488 30540
rect 4448 30433 4476 30534
rect 4434 30424 4490 30433
rect 4434 30359 4490 30368
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 4620 30184 4672 30190
rect 4620 30126 4672 30132
rect 4160 30048 4212 30054
rect 4080 30008 4160 30036
rect 4080 29646 4108 30008
rect 4160 29990 4212 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3608 29572 3660 29578
rect 3608 29514 3660 29520
rect 3712 29566 3832 29594
rect 4068 29640 4120 29646
rect 4068 29582 4120 29588
rect 3620 23050 3648 29514
rect 3712 24818 3740 29566
rect 3792 29504 3844 29510
rect 3792 29446 3844 29452
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3608 23044 3660 23050
rect 3608 22986 3660 22992
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3516 22094 3568 22098
rect 3436 22092 3568 22094
rect 3436 22066 3516 22092
rect 3712 22080 3740 24142
rect 3516 22034 3568 22040
rect 3620 22052 3740 22080
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3330 21312 3386 21321
rect 3330 21247 3386 21256
rect 3344 21078 3372 21247
rect 3332 21072 3384 21078
rect 3332 21014 3384 21020
rect 3344 20398 3372 21014
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3436 16590 3464 19858
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3240 16448 3292 16454
rect 3160 16396 3240 16402
rect 3160 16390 3292 16396
rect 3160 16374 3280 16390
rect 3160 14482 3188 16374
rect 3238 15736 3294 15745
rect 3238 15671 3294 15680
rect 3252 15366 3280 15671
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2976 12434 3004 13126
rect 2976 12406 3188 12434
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2792 11750 2912 11778
rect 2884 11694 2912 11750
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2870 10296 2926 10305
rect 2870 10231 2926 10240
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2516 6886 2636 6914
rect 2516 4826 2544 6886
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2410 4312 2466 4321
rect 2792 4282 2820 7686
rect 2884 5166 2912 10231
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 2962 8800 3018 8809
rect 2962 8735 3018 8744
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2976 4808 3004 8735
rect 3068 5914 3096 9046
rect 3160 8090 3188 12406
rect 3252 11898 3280 15302
rect 3528 13190 3556 20266
rect 3620 17218 3648 22052
rect 3698 21992 3754 22001
rect 3698 21927 3754 21936
rect 3712 20058 3740 21927
rect 3804 20874 3832 29446
rect 3884 29164 3936 29170
rect 4080 29152 4108 29582
rect 3936 29124 4108 29152
rect 3884 29106 3936 29112
rect 3976 29028 4028 29034
rect 3976 28970 4028 28976
rect 3884 28416 3936 28422
rect 3884 28358 3936 28364
rect 3896 28150 3924 28358
rect 3884 28144 3936 28150
rect 3884 28086 3936 28092
rect 3884 27940 3936 27946
rect 3884 27882 3936 27888
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3896 20534 3924 27882
rect 3988 22112 4016 28970
rect 4080 28558 4108 29124
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4632 28665 4660 30126
rect 4618 28656 4674 28665
rect 4618 28591 4674 28600
rect 4068 28552 4120 28558
rect 4068 28494 4120 28500
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4080 27713 4108 28358
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4066 27704 4122 27713
rect 4214 27707 4522 27716
rect 4066 27639 4122 27648
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4080 26353 4108 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4344 26512 4396 26518
rect 4344 26454 4396 26460
rect 4160 26444 4212 26450
rect 4160 26386 4212 26392
rect 4066 26344 4122 26353
rect 4172 26314 4200 26386
rect 4066 26279 4122 26288
rect 4160 26308 4212 26314
rect 4160 26250 4212 26256
rect 4068 25968 4120 25974
rect 4252 25968 4304 25974
rect 4120 25928 4252 25956
rect 4068 25910 4120 25916
rect 4252 25910 4304 25916
rect 4356 25838 4384 26454
rect 4344 25832 4396 25838
rect 4066 25800 4122 25809
rect 4344 25774 4396 25780
rect 4066 25735 4122 25744
rect 4080 24206 4108 25735
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4434 25256 4490 25265
rect 4172 24721 4200 25230
rect 4434 25191 4490 25200
rect 4448 24954 4476 25191
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 4436 24948 4488 24954
rect 4436 24890 4488 24896
rect 4158 24712 4214 24721
rect 4158 24647 4214 24656
rect 4540 24614 4568 25094
rect 4632 24886 4660 28358
rect 4724 26450 4752 31078
rect 5092 30734 5120 31690
rect 5080 30728 5132 30734
rect 5080 30670 5132 30676
rect 5172 30592 5224 30598
rect 5172 30534 5224 30540
rect 5184 30433 5212 30534
rect 5170 30424 5226 30433
rect 5170 30359 5226 30368
rect 5172 30320 5224 30326
rect 5172 30262 5224 30268
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4816 29102 4844 29582
rect 4988 29572 5040 29578
rect 4988 29514 5040 29520
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4816 28082 4844 29038
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4816 27674 4844 28018
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4816 27470 4844 27610
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 4804 27328 4856 27334
rect 4908 27316 4936 28494
rect 5000 27470 5028 29514
rect 5080 29164 5132 29170
rect 5080 29106 5132 29112
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4908 27288 5028 27316
rect 4804 27270 4856 27276
rect 4712 26444 4764 26450
rect 4712 26386 4764 26392
rect 4710 26072 4766 26081
rect 4710 26007 4766 26016
rect 4724 25294 4752 26007
rect 4816 25974 4844 27270
rect 4896 27124 4948 27130
rect 4896 27066 4948 27072
rect 4908 26518 4936 27066
rect 5000 27033 5028 27288
rect 5092 27169 5120 29106
rect 5184 28762 5212 30262
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5264 28416 5316 28422
rect 5264 28358 5316 28364
rect 5172 27328 5224 27334
rect 5172 27270 5224 27276
rect 5078 27160 5134 27169
rect 5078 27095 5134 27104
rect 4986 27024 5042 27033
rect 4986 26959 5042 26968
rect 4988 26852 5040 26858
rect 4988 26794 5040 26800
rect 4896 26512 4948 26518
rect 4896 26454 4948 26460
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4804 25968 4856 25974
rect 4804 25910 4856 25916
rect 4908 25820 4936 26318
rect 4816 25792 4936 25820
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4620 24880 4672 24886
rect 4620 24822 4672 24828
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24290 4660 24618
rect 4724 24410 4752 24890
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4632 24262 4752 24290
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4066 23896 4122 23905
rect 4632 23866 4660 24142
rect 4066 23831 4068 23840
rect 4120 23831 4122 23840
rect 4620 23860 4672 23866
rect 4068 23802 4120 23808
rect 4620 23802 4672 23808
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 23802
rect 4252 23180 4304 23186
rect 4172 23140 4252 23168
rect 4172 22778 4200 23140
rect 4252 23122 4304 23128
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4172 22642 4200 22714
rect 4528 22704 4580 22710
rect 4580 22664 4660 22692
rect 4528 22646 4580 22652
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 4172 22522 4200 22578
rect 4080 22494 4200 22522
rect 3976 22106 4028 22112
rect 3976 22048 4028 22054
rect 4080 22030 4108 22494
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22094 4660 22664
rect 4540 22066 4660 22094
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3974 21176 4030 21185
rect 3974 21111 4030 21120
rect 3988 20806 4016 21111
rect 4080 21010 4108 21966
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4448 21418 4476 21898
rect 4540 21486 4568 22066
rect 4618 21720 4674 21729
rect 4618 21655 4674 21664
rect 4528 21480 4580 21486
rect 4528 21422 4580 21428
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3884 20528 3936 20534
rect 4080 20505 4108 20538
rect 3884 20470 3936 20476
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3896 20262 3924 20334
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 20058 3924 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3698 19952 3754 19961
rect 3698 19887 3754 19896
rect 3712 17610 3740 19887
rect 4632 19786 4660 21655
rect 4724 21570 4752 24262
rect 4816 24138 4844 25792
rect 5000 25226 5028 26794
rect 5080 26784 5132 26790
rect 5080 26726 5132 26732
rect 5092 26518 5120 26726
rect 5080 26512 5132 26518
rect 5080 26454 5132 26460
rect 4988 25220 5040 25226
rect 4988 25162 5040 25168
rect 4986 24984 5042 24993
rect 4986 24919 5042 24928
rect 5000 24750 5028 24919
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 4804 24132 4856 24138
rect 4804 24074 4856 24080
rect 4816 22001 4844 24074
rect 4802 21992 4858 22001
rect 4802 21927 4858 21936
rect 4908 21729 4936 24346
rect 4894 21720 4950 21729
rect 4894 21655 4950 21664
rect 4724 21542 4844 21570
rect 4712 21480 4764 21486
rect 4712 21422 4764 21428
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4724 19718 4752 21422
rect 4816 20641 4844 21542
rect 4802 20632 4858 20641
rect 4802 20567 4858 20576
rect 5000 20534 5028 24686
rect 5078 24440 5134 24449
rect 5078 24375 5134 24384
rect 5092 23662 5120 24375
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 5078 23216 5134 23225
rect 5078 23151 5134 23160
rect 5092 21690 5120 23151
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5092 20874 5120 21626
rect 5184 21622 5212 27270
rect 5276 26042 5304 28358
rect 5368 26568 5396 29446
rect 5460 27334 5488 31826
rect 5644 31754 5672 31894
rect 5644 31726 5764 31754
rect 5540 30660 5592 30666
rect 5540 30602 5592 30608
rect 5552 30258 5580 30602
rect 5736 30274 5764 31726
rect 5828 30734 5856 34682
rect 6840 32910 6868 37130
rect 8404 37126 8432 39200
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8760 36916 8812 36922
rect 8760 36858 8812 36864
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 7196 32768 7248 32774
rect 7196 32710 7248 32716
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 6564 30938 6592 31282
rect 6552 30932 6604 30938
rect 6552 30874 6604 30880
rect 6656 30734 6684 32166
rect 6736 30796 6788 30802
rect 6736 30738 6788 30744
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 6460 30728 6512 30734
rect 6460 30670 6512 30676
rect 6644 30728 6696 30734
rect 6644 30670 6696 30676
rect 5540 30252 5592 30258
rect 5736 30246 6316 30274
rect 5540 30194 5592 30200
rect 5724 30184 5776 30190
rect 5724 30126 5776 30132
rect 5736 28014 5764 30126
rect 6184 29708 6236 29714
rect 6184 29650 6236 29656
rect 6092 29640 6144 29646
rect 6092 29582 6144 29588
rect 6104 28694 6132 29582
rect 6092 28688 6144 28694
rect 6092 28630 6144 28636
rect 6092 28416 6144 28422
rect 6092 28358 6144 28364
rect 5816 28144 5868 28150
rect 5816 28086 5868 28092
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5540 27940 5592 27946
rect 5540 27882 5592 27888
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5448 26920 5500 26926
rect 5448 26862 5500 26868
rect 5460 26761 5488 26862
rect 5446 26752 5502 26761
rect 5446 26687 5502 26696
rect 5368 26540 5488 26568
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5356 25764 5408 25770
rect 5356 25706 5408 25712
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5276 25362 5304 25638
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5276 24886 5304 25298
rect 5264 24880 5316 24886
rect 5264 24822 5316 24828
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5276 23662 5304 24550
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5262 23488 5318 23497
rect 5262 23423 5318 23432
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5172 21480 5224 21486
rect 5172 21422 5224 21428
rect 5184 21321 5212 21422
rect 5170 21312 5226 21321
rect 5170 21247 5226 21256
rect 5170 21176 5226 21185
rect 5170 21111 5226 21120
rect 5080 20868 5132 20874
rect 5080 20810 5132 20816
rect 5078 20768 5134 20777
rect 5078 20703 5134 20712
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 4894 19816 4950 19825
rect 4894 19751 4950 19760
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4802 19408 4858 19417
rect 4802 19343 4858 19352
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18834 4016 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4816 18834 4844 19343
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4710 18592 4766 18601
rect 4710 18527 4766 18536
rect 4160 18352 4212 18358
rect 4212 18312 4292 18340
rect 4160 18294 4212 18300
rect 4264 18222 4292 18312
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3896 17542 3924 18158
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3620 17190 4016 17218
rect 3882 16552 3938 16561
rect 3882 16487 3938 16496
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15366 3740 15846
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 3712 14822 3740 15030
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3712 12866 3740 14758
rect 3896 14346 3924 16487
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13025 3832 13670
rect 3790 13016 3846 13025
rect 3790 12951 3846 12960
rect 3712 12838 3832 12866
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3620 12170 3648 12718
rect 3698 12200 3754 12209
rect 3608 12164 3660 12170
rect 3698 12135 3754 12144
rect 3608 12106 3660 12112
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3424 11280 3476 11286
rect 3422 11248 3424 11257
rect 3476 11248 3478 11257
rect 3422 11183 3478 11192
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3238 10160 3294 10169
rect 3238 10095 3240 10104
rect 3292 10095 3294 10104
rect 3240 10066 3292 10072
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3252 6866 3280 10066
rect 3344 7954 3372 10406
rect 3528 8786 3556 11834
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3620 8956 3648 10678
rect 3712 9110 3740 12135
rect 3804 11898 3832 12838
rect 3896 12442 3924 13874
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 3896 11898 3924 12271
rect 3988 12073 4016 17190
rect 4080 16674 4108 17711
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4264 17241 4292 17546
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17270 4384 17478
rect 4344 17264 4396 17270
rect 4250 17232 4306 17241
rect 4344 17206 4396 17212
rect 4250 17167 4306 17176
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4080 16646 4292 16674
rect 4632 16658 4660 18022
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4080 16425 4108 16458
rect 4066 16416 4122 16425
rect 4066 16351 4122 16360
rect 4264 16114 4292 16646
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4356 16182 4384 16458
rect 4724 16454 4752 18527
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4080 15434 4108 15642
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4264 15026 4292 15574
rect 4620 15428 4672 15434
rect 4620 15370 4672 15376
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4526 14104 4582 14113
rect 4526 14039 4582 14048
rect 4540 14006 4568 14039
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4080 12714 4108 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4158 13016 4214 13025
rect 4448 12986 4476 13194
rect 4158 12951 4214 12960
rect 4436 12980 4488 12986
rect 4172 12918 4200 12951
rect 4436 12922 4488 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4540 12753 4568 12786
rect 4526 12744 4582 12753
rect 4068 12708 4120 12714
rect 4526 12679 4582 12688
rect 4068 12650 4120 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3974 12064 4030 12073
rect 3974 11999 4030 12008
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4080 11778 4108 12378
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11830 4200 12106
rect 3896 11750 4108 11778
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 9722 3832 11630
rect 3896 11121 3924 11750
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 11144 4028 11150
rect 3882 11112 3938 11121
rect 3976 11086 4028 11092
rect 3882 11047 3938 11056
rect 3882 10976 3938 10985
rect 3882 10911 3938 10920
rect 3896 10266 3924 10911
rect 3988 10810 4016 11086
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3988 10674 4016 10746
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3976 9648 4028 9654
rect 3974 9616 3976 9625
rect 4028 9616 4030 9625
rect 4080 9586 4108 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11082 4660 15370
rect 4724 13870 4752 15982
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4816 13530 4844 18770
rect 4908 17270 4936 19751
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4908 13410 4936 16934
rect 5000 16538 5028 17682
rect 5092 16998 5120 20703
rect 5184 17134 5212 21111
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5000 16510 5120 16538
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4816 13382 4936 13410
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10266 4660 10542
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4434 9888 4490 9897
rect 4434 9823 4490 9832
rect 3974 9551 4030 9560
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4448 9518 4476 9823
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4632 9364 4660 10066
rect 4724 9518 4752 12106
rect 4816 11218 4844 13382
rect 5000 13308 5028 16390
rect 5092 14958 5120 16510
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5184 16017 5212 16186
rect 5170 16008 5226 16017
rect 5170 15943 5226 15952
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5078 14784 5134 14793
rect 5078 14719 5134 14728
rect 4908 13280 5028 13308
rect 4908 12170 4936 13280
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 10985 4844 11018
rect 4802 10976 4858 10985
rect 4802 10911 4858 10920
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4632 9336 4752 9364
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 3620 8928 3832 8956
rect 3528 8758 3740 8786
rect 3712 8022 3740 8758
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2976 4780 3096 4808
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2976 4321 3004 4626
rect 2962 4312 3018 4321
rect 2410 4247 2466 4256
rect 2780 4276 2832 4282
rect 2962 4247 3018 4256
rect 2780 4218 2832 4224
rect 1676 4208 1728 4214
rect 1676 4150 1728 4156
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2976 3641 3004 3946
rect 2962 3632 3018 3641
rect 1584 3596 1636 3602
rect 2962 3567 3018 3576
rect 1584 3538 1636 3544
rect 664 3392 716 3398
rect 664 3334 716 3340
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 32 800 60 1294
rect 676 800 704 3334
rect 1596 3058 1624 3538
rect 2962 3360 3018 3369
rect 2962 3295 3018 3304
rect 2976 3058 3004 3295
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1320 800 1348 2790
rect 1596 2514 1624 2994
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2608 800 2636 2926
rect 3068 2774 3096 4780
rect 3344 4758 3372 7278
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3528 6474 3556 6938
rect 3436 6446 3556 6474
rect 3436 6118 3464 6446
rect 3698 6216 3754 6225
rect 3698 6151 3700 6160
rect 3752 6151 3754 6160
rect 3700 6122 3752 6128
rect 3424 6112 3476 6118
rect 3804 6066 3832 8928
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 3988 8401 4016 8842
rect 4172 8430 4200 8842
rect 4264 8498 4292 8978
rect 4342 8936 4398 8945
rect 4342 8871 4344 8880
rect 4396 8871 4398 8880
rect 4344 8842 4396 8848
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4160 8424 4212 8430
rect 3974 8392 4030 8401
rect 4160 8366 4212 8372
rect 3974 8327 4030 8336
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3884 8288 3936 8294
rect 3882 8256 3884 8265
rect 3936 8256 3938 8265
rect 3882 8191 3938 8200
rect 4080 7970 4108 8298
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 7948 3936 7954
rect 4080 7942 4200 7970
rect 4632 7954 4660 8502
rect 3884 7890 3936 7896
rect 3424 6054 3476 6060
rect 3436 5914 3464 6054
rect 3712 6038 3832 6066
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3332 4752 3384 4758
rect 3384 4700 3464 4706
rect 3332 4694 3464 4700
rect 3344 4678 3464 4694
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3160 3194 3188 4218
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3068 2746 3188 2774
rect 3160 2650 3188 2746
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3252 800 3280 4150
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3344 1970 3372 3334
rect 3436 2038 3464 4678
rect 3712 4214 3740 6038
rect 3896 5137 3924 7890
rect 4172 7342 4200 7942
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4160 7336 4212 7342
rect 4066 7304 4122 7313
rect 4160 7278 4212 7284
rect 4066 7239 4122 7248
rect 4080 6730 4108 7239
rect 4540 7206 4568 7414
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 7002 4660 7754
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6390 4200 6598
rect 4540 6458 4568 6802
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3988 5914 4016 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4724 5953 4752 9336
rect 4816 7886 4844 10911
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4816 6730 4844 7346
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4802 6080 4858 6089
rect 4802 6015 4858 6024
rect 4710 5944 4766 5953
rect 3976 5908 4028 5914
rect 4710 5879 4766 5888
rect 3976 5850 4028 5856
rect 3976 5704 4028 5710
rect 4028 5664 4200 5692
rect 3976 5646 4028 5652
rect 4172 5166 4200 5664
rect 4068 5160 4120 5166
rect 3882 5128 3938 5137
rect 4068 5102 4120 5108
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 3882 5063 3938 5072
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3942 3740 4014
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3528 3194 3556 3538
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3528 3097 3556 3130
rect 3514 3088 3570 3097
rect 3712 3058 3740 3878
rect 3804 3505 3832 4694
rect 3896 4282 3924 4966
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3988 4185 4016 4422
rect 3974 4176 4030 4185
rect 3974 4111 4030 4120
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 3514 3023 3570 3032
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3988 2825 4016 3674
rect 4080 3618 4108 5102
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4448 4486 4476 4558
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4080 3590 4292 3618
rect 4632 3602 4660 4966
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4724 4622 4752 4655
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4816 4486 4844 6015
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4908 4128 4936 11630
rect 5000 8294 5028 13126
rect 5092 12900 5120 14719
rect 5184 13172 5212 15943
rect 5276 15910 5304 23423
rect 5368 21690 5396 25706
rect 5460 23186 5488 26540
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5446 22944 5502 22953
rect 5446 22879 5502 22888
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5368 19922 5396 21082
rect 5460 20534 5488 22879
rect 5552 22642 5580 27882
rect 5828 27402 5856 28086
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 5816 27396 5868 27402
rect 5816 27338 5868 27344
rect 5644 25770 5672 27338
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 5736 26897 5764 26930
rect 5722 26888 5778 26897
rect 5722 26823 5778 26832
rect 5828 26466 5856 27338
rect 5736 26438 5856 26466
rect 5736 26314 5764 26438
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5632 25764 5684 25770
rect 5632 25706 5684 25712
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5354 19680 5410 19689
rect 5354 19615 5410 19624
rect 5368 19378 5396 19615
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5356 18760 5408 18766
rect 5354 18728 5356 18737
rect 5408 18728 5410 18737
rect 5354 18663 5410 18672
rect 5460 18154 5488 19722
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17678 5396 18022
rect 5552 17746 5580 22442
rect 5644 22166 5672 23462
rect 5736 23089 5764 25434
rect 5828 23474 5856 26318
rect 5920 26228 5948 27814
rect 6000 27532 6052 27538
rect 6000 27474 6052 27480
rect 6012 26353 6040 27474
rect 5998 26344 6054 26353
rect 5998 26279 6054 26288
rect 5920 26200 6040 26228
rect 5908 25832 5960 25838
rect 5908 25774 5960 25780
rect 5920 24993 5948 25774
rect 6012 25430 6040 26200
rect 6000 25424 6052 25430
rect 6000 25366 6052 25372
rect 5998 25120 6054 25129
rect 5998 25055 6054 25064
rect 5906 24984 5962 24993
rect 5906 24919 5962 24928
rect 6012 24886 6040 25055
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 5920 24410 5948 24686
rect 5908 24404 5960 24410
rect 5908 24346 5960 24352
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 5908 24064 5960 24070
rect 5906 24032 5908 24041
rect 5960 24032 5962 24041
rect 5906 23967 5962 23976
rect 5828 23446 5948 23474
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5722 23080 5778 23089
rect 5722 23015 5778 23024
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5632 22160 5684 22166
rect 5632 22102 5684 22108
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5644 21350 5672 21966
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5356 17672 5408 17678
rect 5644 17626 5672 21286
rect 5356 17614 5408 17620
rect 5552 17598 5672 17626
rect 5446 16688 5502 16697
rect 5356 16652 5408 16658
rect 5446 16623 5502 16632
rect 5356 16594 5408 16600
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5368 15502 5396 16594
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5368 15162 5396 15438
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 14550 5396 15098
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5368 13297 5396 14350
rect 5354 13288 5410 13297
rect 5354 13223 5410 13232
rect 5184 13144 5396 13172
rect 5092 12872 5212 12900
rect 5078 12472 5134 12481
rect 5078 12407 5134 12416
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 5000 7426 5028 7958
rect 5092 7546 5120 12407
rect 5184 12306 5212 12872
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7478 5212 11834
rect 5264 11620 5316 11626
rect 5264 11562 5316 11568
rect 5276 11286 5304 11562
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5172 7472 5224 7478
rect 5000 7398 5120 7426
rect 5172 7414 5224 7420
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 5000 5778 5028 6122
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 5092 5545 5120 7398
rect 5276 7342 5304 11086
rect 5368 8129 5396 13144
rect 5460 12889 5488 16623
rect 5552 14278 5580 17598
rect 5736 15570 5764 22714
rect 5828 21978 5856 23258
rect 5920 22098 5948 23446
rect 6012 22273 6040 24346
rect 5998 22264 6054 22273
rect 5998 22199 6054 22208
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 5998 21992 6054 22001
rect 5828 21950 5948 21978
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5828 19786 5856 21830
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5828 17320 5856 19178
rect 5920 19174 5948 21950
rect 5998 21927 6054 21936
rect 6012 20262 6040 21927
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 6012 18834 6040 19246
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 6104 18086 6132 28358
rect 6196 26858 6224 29650
rect 6184 26852 6236 26858
rect 6184 26794 6236 26800
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6196 24274 6224 26318
rect 6288 25498 6316 30246
rect 6368 29504 6420 29510
rect 6368 29446 6420 29452
rect 6276 25492 6328 25498
rect 6276 25434 6328 25440
rect 6274 25392 6330 25401
rect 6274 25327 6330 25336
rect 6288 25294 6316 25327
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5828 17292 6132 17320
rect 5998 17232 6054 17241
rect 5998 17167 6054 17176
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5828 15094 5856 16730
rect 5908 15428 5960 15434
rect 5908 15370 5960 15376
rect 5816 15088 5868 15094
rect 5816 15030 5868 15036
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5630 14104 5686 14113
rect 5630 14039 5686 14048
rect 5446 12880 5502 12889
rect 5446 12815 5502 12824
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5446 11520 5502 11529
rect 5446 11455 5502 11464
rect 5460 8945 5488 11455
rect 5552 9110 5580 12718
rect 5644 12322 5672 14039
rect 5736 12442 5764 14758
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5828 13258 5856 13466
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5644 12294 5764 12322
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5644 11694 5672 12174
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5736 10180 5764 12294
rect 5828 12102 5856 12718
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11558 5856 12038
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11218 5856 11494
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10282 5856 11018
rect 5920 10441 5948 15370
rect 6012 14482 6040 17167
rect 6104 16794 6132 17292
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6104 14362 6132 16730
rect 6196 16454 6224 22170
rect 6288 22098 6316 23802
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 6276 21956 6328 21962
rect 6276 21898 6328 21904
rect 6288 19242 6316 21898
rect 6380 21010 6408 29446
rect 6472 28150 6500 30670
rect 6552 28484 6604 28490
rect 6552 28426 6604 28432
rect 6460 28144 6512 28150
rect 6460 28086 6512 28092
rect 6564 26330 6592 28426
rect 6748 27112 6776 30738
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 6932 29170 6960 30534
rect 7012 30048 7064 30054
rect 7012 29990 7064 29996
rect 7024 29209 7052 29990
rect 7010 29200 7066 29209
rect 6920 29164 6972 29170
rect 7010 29135 7066 29144
rect 6920 29106 6972 29112
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 6840 27538 6868 29038
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6932 28218 6960 28970
rect 7012 28484 7064 28490
rect 7012 28426 7064 28432
rect 6920 28212 6972 28218
rect 6920 28154 6972 28160
rect 7024 27713 7052 28426
rect 7116 28014 7144 30534
rect 7208 29238 7236 32710
rect 7288 31748 7340 31754
rect 7288 31690 7340 31696
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 7104 27872 7156 27878
rect 7104 27814 7156 27820
rect 7010 27704 7066 27713
rect 7010 27639 7066 27648
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 6748 27084 6868 27112
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6644 26908 6696 26914
rect 6642 26888 6644 26897
rect 6696 26888 6698 26897
rect 6642 26823 6698 26832
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6472 26302 6592 26330
rect 6472 22778 6500 26302
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 6564 23497 6592 26182
rect 6550 23488 6606 23497
rect 6550 23423 6606 23432
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6460 22772 6512 22778
rect 6460 22714 6512 22720
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6472 21010 6500 21626
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6564 20874 6592 22918
rect 6656 22710 6684 26726
rect 6748 25498 6776 26930
rect 6840 26081 6868 27084
rect 6826 26072 6882 26081
rect 6826 26007 6882 26016
rect 6932 25922 6960 27406
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 7024 26790 7052 27338
rect 7012 26784 7064 26790
rect 7012 26726 7064 26732
rect 7012 26308 7064 26314
rect 7012 26250 7064 26256
rect 6840 25894 6960 25922
rect 6840 25514 6868 25894
rect 6920 25832 6972 25838
rect 6918 25800 6920 25809
rect 6972 25800 6974 25809
rect 6918 25735 6974 25744
rect 6736 25492 6788 25498
rect 6840 25486 6960 25514
rect 6736 25434 6788 25440
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6734 24576 6790 24585
rect 6734 24511 6790 24520
rect 6748 24274 6776 24511
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 6748 23526 6776 24210
rect 6840 24206 6868 25094
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6734 23352 6790 23361
rect 6734 23287 6790 23296
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6656 21457 6684 21558
rect 6642 21448 6698 21457
rect 6642 21383 6698 21392
rect 6552 20868 6604 20874
rect 6552 20810 6604 20816
rect 6458 20224 6514 20233
rect 6458 20159 6514 20168
rect 6366 19544 6422 19553
rect 6366 19479 6422 19488
rect 6276 19236 6328 19242
rect 6276 19178 6328 19184
rect 6274 18864 6330 18873
rect 6274 18799 6330 18808
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 14822 6224 15846
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6012 14334 6132 14362
rect 6012 12850 6040 14334
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6104 13938 6132 14214
rect 6288 14056 6316 18799
rect 6380 17814 6408 19479
rect 6472 18290 6500 20159
rect 6642 20088 6698 20097
rect 6642 20023 6698 20032
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6368 17808 6420 17814
rect 6368 17750 6420 17756
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6472 17202 6500 17682
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6380 15366 6408 15506
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6472 15094 6500 17138
rect 6564 16658 6592 18702
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6564 16046 6592 16594
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6368 15088 6420 15094
rect 6366 15056 6368 15065
rect 6460 15088 6512 15094
rect 6420 15056 6422 15065
rect 6460 15030 6512 15036
rect 6366 14991 6422 15000
rect 6564 14482 6592 15982
rect 6656 15910 6684 20023
rect 6748 19446 6776 23287
rect 6840 23032 6868 24142
rect 6932 23905 6960 25486
rect 6918 23896 6974 23905
rect 6918 23831 6974 23840
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6932 23662 6960 23734
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6920 23044 6972 23050
rect 6840 23004 6920 23032
rect 6920 22986 6972 22992
rect 6932 21604 6960 22986
rect 7024 22098 7052 26250
rect 7116 24426 7144 27814
rect 7208 27062 7236 28970
rect 7196 27056 7248 27062
rect 7196 26998 7248 27004
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 7208 24682 7236 26726
rect 7300 25906 7328 31690
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8404 30326 8432 30534
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 8772 30122 8800 36858
rect 9048 36786 9076 39200
rect 10336 37330 10364 39200
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 9128 37256 9180 37262
rect 9128 37198 9180 37204
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 9140 36553 9168 37198
rect 9220 36712 9272 36718
rect 9220 36654 9272 36660
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9126 36544 9182 36553
rect 9126 36479 9182 36488
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 9036 30728 9088 30734
rect 9036 30670 9088 30676
rect 8944 30320 8996 30326
rect 8944 30262 8996 30268
rect 8852 30184 8904 30190
rect 8850 30152 8852 30161
rect 8904 30152 8906 30161
rect 8760 30116 8812 30122
rect 8850 30087 8906 30096
rect 8760 30058 8812 30064
rect 7748 30048 7800 30054
rect 7748 29990 7800 29996
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 7564 29844 7616 29850
rect 7564 29786 7616 29792
rect 7472 29504 7524 29510
rect 7472 29446 7524 29452
rect 7380 28144 7432 28150
rect 7380 28086 7432 28092
rect 7392 26994 7420 28086
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7392 26353 7420 26726
rect 7378 26344 7434 26353
rect 7378 26279 7434 26288
rect 7288 25900 7340 25906
rect 7288 25842 7340 25848
rect 7300 25809 7328 25842
rect 7286 25800 7342 25809
rect 7286 25735 7342 25744
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7300 24886 7328 25434
rect 7288 24880 7340 24886
rect 7288 24822 7340 24828
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 7116 24398 7236 24426
rect 7102 24168 7158 24177
rect 7102 24103 7104 24112
rect 7156 24103 7158 24112
rect 7104 24074 7156 24080
rect 7208 23526 7236 24398
rect 7300 23594 7328 24822
rect 7484 24070 7512 29446
rect 7576 29034 7604 29786
rect 7656 29232 7708 29238
rect 7656 29174 7708 29180
rect 7564 29028 7616 29034
rect 7564 28970 7616 28976
rect 7564 28552 7616 28558
rect 7564 28494 7616 28500
rect 7472 24064 7524 24070
rect 7576 24041 7604 28494
rect 7472 24006 7524 24012
rect 7562 24032 7618 24041
rect 7562 23967 7618 23976
rect 7668 23882 7696 29174
rect 7760 29073 7788 29990
rect 7840 29504 7892 29510
rect 7840 29446 7892 29452
rect 7932 29504 7984 29510
rect 7932 29446 7984 29452
rect 7746 29064 7802 29073
rect 7746 28999 7802 29008
rect 7748 27940 7800 27946
rect 7748 27882 7800 27888
rect 7760 25401 7788 27882
rect 7746 25392 7802 25401
rect 7746 25327 7802 25336
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7760 24410 7788 24754
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7746 24304 7802 24313
rect 7746 24239 7802 24248
rect 7392 23854 7696 23882
rect 7288 23588 7340 23594
rect 7288 23530 7340 23536
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 7012 21616 7064 21622
rect 6932 21576 7012 21604
rect 6828 21412 6880 21418
rect 6828 21354 6880 21360
rect 6840 21049 6868 21354
rect 6826 21040 6882 21049
rect 6826 20975 6882 20984
rect 6932 20466 6960 21576
rect 7012 21558 7064 21564
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6932 19922 6960 20402
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6748 17610 6776 19382
rect 6932 19378 6960 19858
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17746 6868 18158
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 17785 6960 18022
rect 6918 17776 6974 17785
rect 6828 17740 6880 17746
rect 6918 17711 6974 17720
rect 6828 17682 6880 17688
rect 6918 17640 6974 17649
rect 6736 17604 6788 17610
rect 6918 17575 6974 17584
rect 6736 17546 6788 17552
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6748 16153 6776 16458
rect 6734 16144 6790 16153
rect 6734 16079 6790 16088
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6288 14028 6408 14056
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5906 10432 5962 10441
rect 5906 10367 5962 10376
rect 5828 10254 6040 10282
rect 5736 10152 5856 10180
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9761 5672 9930
rect 5630 9752 5686 9761
rect 5630 9687 5686 9696
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5446 8936 5502 8945
rect 5446 8871 5502 8880
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8362 5672 8434
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5354 8120 5410 8129
rect 5354 8055 5410 8064
rect 5828 7993 5856 10152
rect 5906 10160 5962 10169
rect 5906 10095 5962 10104
rect 5814 7984 5870 7993
rect 5814 7919 5816 7928
rect 5868 7919 5870 7928
rect 5816 7890 5868 7896
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5460 6866 5488 7822
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7546 5764 7754
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5078 5536 5134 5545
rect 5078 5471 5134 5480
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 5030 5028 5102
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5368 4622 5396 5782
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4908 4100 5304 4128
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 2990 4200 3470
rect 4264 3233 4292 3590
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4724 3466 4752 3538
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4250 3224 4306 3233
rect 4250 3159 4306 3168
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 4080 2650 4108 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4620 2576 4672 2582
rect 4618 2544 4620 2553
rect 4672 2544 4674 2553
rect 4618 2479 4674 2488
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3516 808 3568 814
rect 18 200 74 800
rect 662 200 718 800
rect 1306 200 1362 800
rect 2594 200 2650 800
rect 3238 200 3294 800
rect 3514 776 3516 785
rect 3896 800 3924 2246
rect 5092 1306 5120 2314
rect 5184 1873 5212 3946
rect 5276 2774 5304 4100
rect 5368 3942 5396 4558
rect 5460 3942 5488 6122
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5354 3088 5410 3097
rect 5552 3040 5580 7278
rect 5736 6390 5764 7482
rect 5920 7154 5948 10095
rect 6012 8906 6040 10254
rect 6104 9382 6132 13194
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6012 8265 6040 8842
rect 5998 8256 6054 8265
rect 5998 8191 6054 8200
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6012 7274 6040 7686
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5920 7126 6040 7154
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5722 6216 5778 6225
rect 5722 6151 5778 6160
rect 5736 5846 5764 6151
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5736 5114 5764 5782
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5736 5086 5856 5114
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4554 5764 4966
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5354 3023 5356 3032
rect 5408 3023 5410 3032
rect 5356 2994 5408 3000
rect 5460 3012 5580 3040
rect 5276 2746 5396 2774
rect 5262 2680 5318 2689
rect 5262 2615 5318 2624
rect 5276 2582 5304 2615
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5368 1970 5396 2746
rect 5460 2666 5488 3012
rect 5538 2952 5594 2961
rect 5538 2887 5594 2896
rect 5552 2854 5580 2887
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5828 2774 5856 5086
rect 5920 4026 5948 5306
rect 6012 4185 6040 7126
rect 6090 5400 6146 5409
rect 6090 5335 6146 5344
rect 6104 5302 6132 5335
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 5998 4176 6054 4185
rect 5998 4111 6054 4120
rect 5920 3998 6132 4026
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 5736 2746 5856 2774
rect 5460 2638 5580 2666
rect 5736 2650 5764 2746
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 5170 1864 5226 1873
rect 5170 1799 5226 1808
rect 5092 1278 5212 1306
rect 5552 1290 5580 2638
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5184 800 5212 1278
rect 5540 1284 5592 1290
rect 5540 1226 5592 1232
rect 5828 800 5856 2246
rect 5920 1426 5948 2926
rect 6012 1834 6040 3470
rect 6104 2281 6132 3998
rect 6196 2774 6224 11630
rect 6288 11218 6316 13874
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6288 9489 6316 9522
rect 6274 9480 6330 9489
rect 6274 9415 6330 9424
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6288 7342 6316 7890
rect 6380 7478 6408 14028
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6564 13326 6592 13738
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6564 12782 6592 13262
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6656 12434 6684 15302
rect 6932 14890 6960 17575
rect 7024 16114 7052 20810
rect 7116 19281 7144 23462
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7300 22438 7328 22578
rect 7392 22574 7420 23854
rect 7470 23760 7526 23769
rect 7760 23746 7788 24239
rect 7470 23695 7526 23704
rect 7576 23718 7788 23746
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7286 21992 7342 22001
rect 7286 21927 7342 21936
rect 7196 21888 7248 21894
rect 7196 21830 7248 21836
rect 7208 21554 7236 21830
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7208 20534 7236 21490
rect 7196 20528 7248 20534
rect 7196 20470 7248 20476
rect 7300 20398 7328 21927
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7102 19272 7158 19281
rect 7102 19207 7158 19216
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 16250 7144 18022
rect 7194 17912 7250 17921
rect 7194 17847 7250 17856
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7208 15552 7236 17847
rect 7024 15524 7236 15552
rect 7288 15564 7340 15570
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6826 14376 6882 14385
rect 6826 14311 6828 14320
rect 6880 14311 6882 14320
rect 6828 14282 6880 14288
rect 6826 14240 6882 14249
rect 6826 14175 6882 14184
rect 6734 13560 6790 13569
rect 6734 13495 6790 13504
rect 6748 13258 6776 13495
rect 6840 13258 6868 14175
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6564 12406 6684 12434
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 7472 6420 7478
rect 6472 7449 6500 11698
rect 6564 7478 6592 12406
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 11762 6776 12242
rect 6840 11898 6868 13194
rect 6932 13025 6960 13670
rect 6918 13016 6974 13025
rect 6918 12951 6974 12960
rect 6932 12918 6960 12951
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 7024 12209 7052 15524
rect 7288 15506 7340 15512
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7116 12434 7144 13194
rect 7116 12406 7236 12434
rect 7010 12200 7066 12209
rect 7010 12135 7066 12144
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6734 11248 6790 11257
rect 6734 11183 6790 11192
rect 6828 11212 6880 11218
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10713 6684 10746
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 10130 6684 10542
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6748 9874 6776 11183
rect 6828 11154 6880 11160
rect 6656 9846 6776 9874
rect 6552 7472 6604 7478
rect 6368 7414 6420 7420
rect 6458 7440 6514 7449
rect 6552 7414 6604 7420
rect 6458 7375 6514 7384
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 5778 6316 6734
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5302 6316 5714
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6380 5098 6408 6870
rect 6656 6848 6684 9846
rect 6840 9353 6868 11154
rect 6920 11144 6972 11150
rect 6972 11104 7052 11132
rect 6920 11086 6972 11092
rect 6826 9344 6882 9353
rect 6826 9279 6882 9288
rect 6828 9104 6880 9110
rect 6826 9072 6828 9081
rect 6880 9072 6882 9081
rect 6826 9007 6882 9016
rect 6828 8968 6880 8974
rect 6880 8928 6960 8956
rect 6828 8910 6880 8916
rect 6932 8430 6960 8928
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6472 6820 6684 6848
rect 6472 5681 6500 6820
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6458 5672 6514 5681
rect 6458 5607 6514 5616
rect 6564 5370 6592 5714
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6472 5148 6500 5238
rect 6541 5160 6593 5166
rect 6472 5120 6541 5148
rect 6541 5102 6593 5108
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6380 2825 6408 5034
rect 6550 4040 6606 4049
rect 6460 4004 6512 4010
rect 6550 3975 6606 3984
rect 6460 3946 6512 3952
rect 6366 2816 6422 2825
rect 6196 2746 6316 2774
rect 6366 2751 6422 2760
rect 6090 2272 6146 2281
rect 6090 2207 6146 2216
rect 6288 2106 6316 2746
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6000 1828 6052 1834
rect 6000 1770 6052 1776
rect 6472 1465 6500 3946
rect 6564 3534 6592 3975
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6564 2961 6592 2994
rect 6550 2952 6606 2961
rect 6550 2887 6606 2896
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 1698 6592 2246
rect 6656 1766 6684 6666
rect 6840 6497 6868 8230
rect 6932 8022 6960 8366
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 7024 7800 7052 11104
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7116 10130 7144 10202
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7208 8673 7236 12406
rect 7300 12102 7328 15506
rect 7392 14482 7420 22510
rect 7484 22506 7512 23695
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7576 22137 7604 23718
rect 7656 23588 7708 23594
rect 7656 23530 7708 23536
rect 7562 22128 7618 22137
rect 7562 22063 7618 22072
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7470 21720 7526 21729
rect 7470 21655 7526 21664
rect 7484 21486 7512 21655
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7470 21312 7526 21321
rect 7470 21247 7526 21256
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7378 12064 7434 12073
rect 7378 11999 7434 12008
rect 7392 11082 7420 11999
rect 7484 11218 7512 21247
rect 7576 20874 7604 21966
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7562 20496 7618 20505
rect 7562 20431 7618 20440
rect 7576 16658 7604 20431
rect 7668 19938 7696 23530
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7760 20856 7788 23462
rect 7852 21729 7880 29446
rect 7944 26314 7972 29446
rect 7932 26308 7984 26314
rect 7932 26250 7984 26256
rect 8024 26308 8076 26314
rect 8024 26250 8076 26256
rect 8036 25974 8064 26250
rect 8024 25968 8076 25974
rect 8024 25910 8076 25916
rect 8128 25820 8156 29990
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 8220 29170 8248 29786
rect 8772 29646 8800 30058
rect 8668 29640 8720 29646
rect 8668 29582 8720 29588
rect 8760 29640 8812 29646
rect 8760 29582 8812 29588
rect 8680 29345 8708 29582
rect 8298 29336 8354 29345
rect 8298 29271 8354 29280
rect 8666 29336 8722 29345
rect 8666 29271 8722 29280
rect 8850 29336 8906 29345
rect 8956 29306 8984 30262
rect 8850 29271 8906 29280
rect 8944 29300 8996 29306
rect 8312 29170 8340 29271
rect 8208 29164 8260 29170
rect 8208 29106 8260 29112
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8300 28484 8352 28490
rect 8300 28426 8352 28432
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8220 26926 8248 27474
rect 8208 26920 8260 26926
rect 8206 26888 8208 26897
rect 8260 26888 8262 26897
rect 8206 26823 8262 26832
rect 8312 25974 8340 28426
rect 8760 28416 8812 28422
rect 8760 28358 8812 28364
rect 8482 28112 8538 28121
rect 8482 28047 8484 28056
rect 8536 28047 8538 28056
rect 8484 28018 8536 28024
rect 8484 27940 8536 27946
rect 8484 27882 8536 27888
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8404 27441 8432 27814
rect 8390 27432 8446 27441
rect 8390 27367 8446 27376
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 8404 25838 8432 27270
rect 8036 25792 8156 25820
rect 8392 25832 8444 25838
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7838 21720 7894 21729
rect 7838 21655 7894 21664
rect 7760 20828 7880 20856
rect 7668 19910 7788 19938
rect 7760 19446 7788 19910
rect 7852 19786 7880 20828
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7748 19440 7800 19446
rect 7654 19408 7710 19417
rect 7748 19382 7800 19388
rect 7654 19343 7710 19352
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7668 16266 7696 19343
rect 7748 19304 7800 19310
rect 7746 19272 7748 19281
rect 7800 19272 7802 19281
rect 7746 19207 7802 19216
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7852 18057 7880 18158
rect 7838 18048 7894 18057
rect 7838 17983 7894 17992
rect 7944 17218 7972 23666
rect 8036 23186 8064 25792
rect 8392 25774 8444 25780
rect 8116 25424 8168 25430
rect 8116 25366 8168 25372
rect 8128 25265 8156 25366
rect 8114 25256 8170 25265
rect 8114 25191 8170 25200
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8128 24449 8156 25094
rect 8220 24954 8248 25094
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8300 24948 8352 24954
rect 8300 24890 8352 24896
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8114 24440 8170 24449
rect 8114 24375 8170 24384
rect 8128 23594 8156 24375
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8114 23488 8170 23497
rect 8114 23423 8170 23432
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8036 22273 8064 22510
rect 8022 22264 8078 22273
rect 8022 22199 8078 22208
rect 8022 22128 8078 22137
rect 8022 22063 8078 22072
rect 8036 18714 8064 22063
rect 8128 20806 8156 23423
rect 8220 22080 8248 24550
rect 8312 23662 8340 24890
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8404 24274 8432 24686
rect 8496 24313 8524 27882
rect 8668 27872 8720 27878
rect 8668 27814 8720 27820
rect 8576 25968 8628 25974
rect 8576 25910 8628 25916
rect 8482 24304 8538 24313
rect 8392 24268 8444 24274
rect 8482 24239 8538 24248
rect 8392 24210 8444 24216
rect 8404 23662 8432 24210
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8404 23186 8432 23598
rect 8588 23254 8616 25910
rect 8680 25226 8708 27814
rect 8772 27713 8800 28358
rect 8758 27704 8814 27713
rect 8758 27639 8814 27648
rect 8760 27464 8812 27470
rect 8758 27432 8760 27441
rect 8812 27432 8814 27441
rect 8758 27367 8814 27376
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 8680 24410 8708 25162
rect 8668 24404 8720 24410
rect 8668 24346 8720 24352
rect 8772 24290 8800 27367
rect 8864 25974 8892 29271
rect 8944 29242 8996 29248
rect 9048 28218 9076 30670
rect 9140 29594 9168 31214
rect 9232 30326 9260 36654
rect 9220 30320 9272 30326
rect 9220 30262 9272 30268
rect 9232 30190 9260 30262
rect 9220 30184 9272 30190
rect 9220 30126 9272 30132
rect 9312 30184 9364 30190
rect 9312 30126 9364 30132
rect 9140 29566 9260 29594
rect 9128 29504 9180 29510
rect 9128 29446 9180 29452
rect 9036 28212 9088 28218
rect 9036 28154 9088 28160
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8852 25968 8904 25974
rect 8852 25910 8904 25916
rect 8850 25800 8906 25809
rect 8850 25735 8906 25744
rect 8680 24262 8800 24290
rect 8680 23254 8708 24262
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 8576 23248 8628 23254
rect 8496 23208 8576 23236
rect 8392 23180 8444 23186
rect 8392 23122 8444 23128
rect 8392 23044 8444 23050
rect 8392 22986 8444 22992
rect 8220 22052 8340 22080
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8220 21185 8248 21898
rect 8206 21176 8262 21185
rect 8206 21111 8262 21120
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8116 20800 8168 20806
rect 8220 20777 8248 20946
rect 8116 20742 8168 20748
rect 8206 20768 8262 20777
rect 8206 20703 8262 20712
rect 8312 20618 8340 22052
rect 8404 21486 8432 22986
rect 8496 21706 8524 23208
rect 8576 23190 8628 23196
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8588 21865 8616 22510
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8680 22001 8708 22034
rect 8666 21992 8722 22001
rect 8666 21927 8722 21936
rect 8668 21888 8720 21894
rect 8574 21856 8630 21865
rect 8668 21830 8720 21836
rect 8574 21791 8630 21800
rect 8496 21678 8616 21706
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8220 20590 8340 20618
rect 8220 20346 8248 20590
rect 8128 20318 8248 20346
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8128 18902 8156 20318
rect 8312 19258 8340 20334
rect 8404 19854 8432 21082
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8312 19230 8432 19258
rect 8300 19168 8352 19174
rect 8206 19136 8262 19145
rect 8300 19110 8352 19116
rect 8206 19071 8262 19080
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8036 18686 8156 18714
rect 7576 16238 7696 16266
rect 7760 17190 7972 17218
rect 7576 14793 7604 16238
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7668 15434 7696 16118
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7562 14784 7618 14793
rect 7562 14719 7618 14728
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7576 13410 7604 14554
rect 7576 13382 7696 13410
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7194 8664 7250 8673
rect 7194 8599 7250 8608
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 6932 7772 7052 7800
rect 6826 6488 6882 6497
rect 6826 6423 6882 6432
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6748 2774 6776 5850
rect 6932 5794 6960 7772
rect 7116 7342 7144 7958
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7116 6866 7144 7278
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7024 5914 7052 6666
rect 7116 6390 7144 6802
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6932 5766 7052 5794
rect 6918 5672 6974 5681
rect 6828 5636 6880 5642
rect 6918 5607 6974 5616
rect 6828 5578 6880 5584
rect 6840 5114 6868 5578
rect 6932 5370 6960 5607
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6920 5160 6972 5166
rect 6840 5108 6920 5114
rect 6840 5102 6972 5108
rect 6840 5086 6960 5102
rect 7024 4457 7052 5766
rect 7102 5400 7158 5409
rect 7102 5335 7104 5344
rect 7156 5335 7158 5344
rect 7104 5306 7156 5312
rect 7208 4622 7236 8502
rect 7300 5273 7328 10950
rect 7392 10033 7420 11018
rect 7378 10024 7434 10033
rect 7378 9959 7434 9968
rect 7472 9988 7524 9994
rect 7392 7954 7420 9959
rect 7472 9930 7524 9936
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7286 5264 7342 5273
rect 7286 5199 7342 5208
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7196 4616 7248 4622
rect 7300 4593 7328 4694
rect 7196 4558 7248 4564
rect 7286 4584 7342 4593
rect 7286 4519 7342 4528
rect 7010 4448 7066 4457
rect 7010 4383 7066 4392
rect 7300 4128 7328 4519
rect 7208 4100 7328 4128
rect 7208 3602 7236 4100
rect 7286 4040 7342 4049
rect 7286 3975 7342 3984
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7300 3058 7328 3975
rect 7392 3398 7420 7414
rect 7484 7041 7512 9930
rect 7562 9208 7618 9217
rect 7562 9143 7618 9152
rect 7576 9042 7604 9143
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7470 7032 7526 7041
rect 7470 6967 7526 6976
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7484 6458 7512 6666
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6748 2746 6868 2774
rect 6840 2553 6868 2746
rect 6826 2544 6882 2553
rect 6826 2479 6882 2488
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 6644 1760 6696 1766
rect 6644 1702 6696 1708
rect 6552 1692 6604 1698
rect 6552 1634 6604 1640
rect 6458 1456 6514 1465
rect 5908 1420 5960 1426
rect 6458 1391 6514 1400
rect 5908 1362 5960 1368
rect 7116 800 7144 2246
rect 7576 1562 7604 8842
rect 7668 4826 7696 13382
rect 7760 11937 7788 17190
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7944 15473 7972 15506
rect 7930 15464 7986 15473
rect 8128 15434 8156 18686
rect 8220 18290 8248 19071
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8312 17882 8340 19110
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8220 16833 8248 17546
rect 8404 17082 8432 19230
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8496 18630 8524 19110
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8496 17678 8524 18566
rect 8588 18222 8616 21678
rect 8680 20942 8708 21830
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8666 20360 8722 20369
rect 8666 20295 8722 20304
rect 8680 19718 8708 20295
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8772 18698 8800 24006
rect 8864 23662 8892 25735
rect 8956 23905 8984 28018
rect 9036 26376 9088 26382
rect 9140 26364 9168 29446
rect 9232 28994 9260 29566
rect 9324 29238 9352 30126
rect 9312 29232 9364 29238
rect 9312 29174 9364 29180
rect 9416 29170 9444 36654
rect 10324 36644 10376 36650
rect 10324 36586 10376 36592
rect 10232 31136 10284 31142
rect 10232 31078 10284 31084
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 9232 28966 9352 28994
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 9232 27130 9260 27338
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 9324 27010 9352 28966
rect 9416 28694 9444 29106
rect 9404 28688 9456 28694
rect 9404 28630 9456 28636
rect 9404 28552 9456 28558
rect 9402 28520 9404 28529
rect 9456 28520 9458 28529
rect 9402 28455 9458 28464
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9088 26336 9168 26364
rect 9232 26982 9352 27010
rect 9036 26318 9088 26324
rect 9036 26240 9088 26246
rect 9036 26182 9088 26188
rect 9048 25820 9076 26182
rect 9128 25832 9180 25838
rect 9048 25792 9128 25820
rect 8942 23896 8998 23905
rect 8942 23831 8998 23840
rect 8944 23792 8996 23798
rect 8944 23734 8996 23740
rect 8956 23662 8984 23734
rect 8852 23656 8904 23662
rect 8852 23598 8904 23604
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 8864 23497 8892 23598
rect 8850 23488 8906 23497
rect 8850 23423 8906 23432
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 8850 21992 8906 22001
rect 8850 21927 8906 21936
rect 8864 21622 8892 21927
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8666 18456 8722 18465
rect 8666 18391 8722 18400
rect 8576 18216 8628 18222
rect 8574 18184 8576 18193
rect 8628 18184 8630 18193
rect 8574 18119 8630 18128
rect 8574 18048 8630 18057
rect 8574 17983 8630 17992
rect 8588 17746 8616 17983
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8574 17368 8630 17377
rect 8574 17303 8630 17312
rect 8404 17054 8524 17082
rect 8588 17066 8616 17303
rect 8206 16824 8262 16833
rect 8206 16759 8262 16768
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 7930 15399 7986 15408
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 7838 15192 7894 15201
rect 7838 15127 7840 15136
rect 7892 15127 7894 15136
rect 7840 15098 7892 15104
rect 7852 13852 7880 15098
rect 8022 14920 8078 14929
rect 8022 14855 8078 14864
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7944 14006 7972 14486
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 7852 13824 7972 13852
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7746 11928 7802 11937
rect 7746 11863 7802 11872
rect 7746 11792 7802 11801
rect 7746 11727 7802 11736
rect 7760 8294 7788 11727
rect 7852 9518 7880 12310
rect 7944 12073 7972 13824
rect 7930 12064 7986 12073
rect 7930 11999 7986 12008
rect 8036 11234 8064 14855
rect 8220 14793 8248 16458
rect 8206 14784 8262 14793
rect 8206 14719 8262 14728
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 12617 8156 14282
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8114 12608 8170 12617
rect 8114 12543 8170 12552
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8128 11370 8156 12106
rect 8220 11529 8248 12854
rect 8312 12442 8340 16662
rect 8496 15450 8524 17054
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8574 16688 8630 16697
rect 8574 16623 8630 16632
rect 8588 16590 8616 16623
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8404 15434 8524 15450
rect 8392 15428 8524 15434
rect 8444 15422 8524 15428
rect 8392 15370 8444 15376
rect 8392 13864 8444 13870
rect 8588 13852 8616 16526
rect 8680 16522 8708 18391
rect 8772 17814 8800 18634
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8772 16998 8800 17206
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8772 16425 8800 16594
rect 8864 16454 8892 20810
rect 8852 16448 8904 16454
rect 8758 16416 8814 16425
rect 8852 16390 8904 16396
rect 8758 16351 8814 16360
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8680 15570 8708 15982
rect 8850 15872 8906 15881
rect 8850 15807 8906 15816
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8444 13824 8616 13852
rect 8392 13806 8444 13812
rect 8588 13433 8616 13824
rect 8574 13424 8630 13433
rect 8574 13359 8630 13368
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8404 12322 8432 13194
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8496 12714 8524 12922
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8312 12294 8432 12322
rect 8312 12238 8340 12294
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8390 12200 8446 12209
rect 8390 12135 8392 12144
rect 8444 12135 8446 12144
rect 8392 12106 8444 12112
rect 8404 11665 8432 12106
rect 8390 11656 8446 11665
rect 8390 11591 8446 11600
rect 8206 11520 8262 11529
rect 8206 11455 8262 11464
rect 8128 11342 8248 11370
rect 7932 11212 7984 11218
rect 8036 11206 8156 11234
rect 7932 11154 7984 11160
rect 7944 11121 7972 11154
rect 7930 11112 7986 11121
rect 7930 11047 7986 11056
rect 7944 9994 7972 11047
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7838 8664 7894 8673
rect 7838 8599 7894 8608
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7954 7788 8230
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7746 7440 7802 7449
rect 7746 7375 7802 7384
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4729 7788 7375
rect 7852 7290 7880 8599
rect 7932 7472 7984 7478
rect 7930 7440 7932 7449
rect 7984 7440 7986 7449
rect 7930 7375 7986 7384
rect 7852 7262 7972 7290
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5710 7880 6054
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7746 4720 7802 4729
rect 7746 4655 7802 4664
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 4162 7696 4558
rect 7668 4134 7788 4162
rect 7760 3913 7788 4134
rect 7746 3904 7802 3913
rect 7746 3839 7802 3848
rect 7944 3777 7972 7262
rect 7930 3768 7986 3777
rect 7930 3703 7986 3712
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7564 1556 7616 1562
rect 7564 1498 7616 1504
rect 7760 800 7788 3334
rect 8036 1494 8064 10610
rect 8128 9994 8156 11206
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 7018 8156 8774
rect 8220 7721 8248 11342
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8298 10704 8354 10713
rect 8298 10639 8300 10648
rect 8352 10639 8354 10648
rect 8300 10610 8352 10616
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 9178 8340 9318
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8206 7712 8262 7721
rect 8206 7647 8262 7656
rect 8128 6990 8248 7018
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8128 6322 8156 6870
rect 8220 6458 8248 6990
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8128 5681 8156 6122
rect 8114 5672 8170 5681
rect 8114 5607 8170 5616
rect 8404 5534 8432 11018
rect 8496 9654 8524 12378
rect 8574 12336 8630 12345
rect 8574 12271 8630 12280
rect 8588 12238 8616 12271
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8588 9897 8616 11999
rect 8680 11898 8708 15370
rect 8772 14414 8800 15438
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8680 10985 8708 11018
rect 8666 10976 8722 10985
rect 8666 10911 8722 10920
rect 8772 10198 8800 14350
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8574 9888 8630 9897
rect 8574 9823 8630 9832
rect 8758 9752 8814 9761
rect 8758 9687 8814 9696
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8482 9480 8538 9489
rect 8482 9415 8538 9424
rect 8496 5914 8524 9415
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8588 8838 8616 9318
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8220 5506 8432 5534
rect 8220 4826 8248 5506
rect 8482 5400 8538 5409
rect 8482 5335 8538 5344
rect 8496 5234 8524 5335
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8298 4856 8354 4865
rect 8208 4820 8260 4826
rect 8298 4791 8354 4800
rect 8208 4762 8260 4768
rect 8220 4622 8248 4762
rect 8312 4758 8340 4791
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8404 4486 8432 4966
rect 8588 4672 8616 8502
rect 8680 8090 8708 9318
rect 8772 8673 8800 9687
rect 8758 8664 8814 8673
rect 8758 8599 8814 8608
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8666 7848 8722 7857
rect 8666 7783 8722 7792
rect 8680 6474 8708 7783
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7585 8800 7686
rect 8758 7576 8814 7585
rect 8758 7511 8814 7520
rect 8680 6446 8800 6474
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8680 5817 8708 6326
rect 8666 5808 8722 5817
rect 8666 5743 8722 5752
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8680 5409 8708 5646
rect 8666 5400 8722 5409
rect 8666 5335 8722 5344
rect 8772 4826 8800 6446
rect 8864 5370 8892 15807
rect 8956 13326 8984 23190
rect 9048 20874 9076 25792
rect 9128 25774 9180 25780
rect 9128 25356 9180 25362
rect 9128 25298 9180 25304
rect 9140 24993 9168 25298
rect 9126 24984 9182 24993
rect 9126 24919 9182 24928
rect 9128 24744 9180 24750
rect 9126 24712 9128 24721
rect 9180 24712 9182 24721
rect 9126 24647 9182 24656
rect 9232 24410 9260 26982
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9324 26314 9352 26522
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9312 25424 9364 25430
rect 9312 25366 9364 25372
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9232 22574 9260 24346
rect 9324 23361 9352 25366
rect 9310 23352 9366 23361
rect 9310 23287 9366 23296
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22642 9352 23054
rect 9312 22636 9364 22642
rect 9312 22578 9364 22584
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22234 9168 22442
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 9220 22228 9272 22234
rect 9220 22170 9272 22176
rect 9232 21690 9260 22170
rect 9416 21962 9444 27474
rect 9508 27062 9536 30534
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 9862 30016 9918 30025
rect 9862 29951 9918 29960
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 9784 29617 9812 29650
rect 9770 29608 9826 29617
rect 9876 29578 9904 29951
rect 9968 29753 9996 30262
rect 10140 30252 10192 30258
rect 10060 30212 10140 30240
rect 9954 29744 10010 29753
rect 9954 29679 10010 29688
rect 9770 29543 9826 29552
rect 9864 29572 9916 29578
rect 9864 29514 9916 29520
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9784 28966 9812 29446
rect 10060 28994 10088 30212
rect 10140 30194 10192 30200
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10152 29481 10180 29582
rect 10138 29472 10194 29481
rect 10138 29407 10194 29416
rect 10244 29238 10272 31078
rect 10232 29232 10284 29238
rect 10232 29174 10284 29180
rect 10060 28966 10180 28994
rect 9772 28960 9824 28966
rect 9772 28902 9824 28908
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 9588 28484 9640 28490
rect 9588 28426 9640 28432
rect 9600 28121 9628 28426
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9678 28248 9734 28257
rect 9678 28183 9734 28192
rect 9692 28150 9720 28183
rect 9784 28150 9812 28358
rect 9680 28144 9732 28150
rect 9586 28112 9642 28121
rect 9680 28086 9732 28092
rect 9772 28144 9824 28150
rect 9772 28086 9824 28092
rect 9586 28047 9642 28056
rect 9586 27704 9642 27713
rect 9642 27662 9720 27690
rect 9876 27674 9904 28494
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9968 27713 9996 28018
rect 9954 27704 10010 27713
rect 9586 27639 9642 27648
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 9496 27056 9548 27062
rect 9496 26998 9548 27004
rect 9494 26616 9550 26625
rect 9494 26551 9550 26560
rect 9508 26246 9536 26551
rect 9496 26240 9548 26246
rect 9496 26182 9548 26188
rect 9600 25838 9628 27474
rect 9692 27402 9720 27662
rect 9772 27668 9824 27674
rect 9772 27610 9824 27616
rect 9864 27668 9916 27674
rect 9954 27639 10010 27648
rect 9864 27610 9916 27616
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9784 26217 9812 27610
rect 10060 27606 10088 28358
rect 10152 28082 10180 28966
rect 10336 28558 10364 36586
rect 10508 34400 10560 34406
rect 10508 34342 10560 34348
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10428 28778 10456 30670
rect 10520 29714 10548 34342
rect 10612 31754 10640 37198
rect 10784 37188 10836 37194
rect 10784 37130 10836 37136
rect 10692 36576 10744 36582
rect 10692 36518 10744 36524
rect 10704 35086 10732 36518
rect 10692 35080 10744 35086
rect 10692 35022 10744 35028
rect 10796 34610 10824 37130
rect 10980 36938 11008 39200
rect 11624 37126 11652 39200
rect 12912 37126 12940 39200
rect 13556 37262 13584 39200
rect 14844 37330 14872 39200
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 12992 37256 13044 37262
rect 12992 37198 13044 37204
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 11612 37120 11664 37126
rect 11612 37062 11664 37068
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 10980 36922 11100 36938
rect 10980 36916 11112 36922
rect 10980 36910 11060 36916
rect 11060 36858 11112 36864
rect 11704 36780 11756 36786
rect 11704 36722 11756 36728
rect 10968 36712 11020 36718
rect 10968 36654 11020 36660
rect 10980 36242 11008 36654
rect 10968 36236 11020 36242
rect 10968 36178 11020 36184
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 10612 31726 10732 31754
rect 10704 30394 10732 31726
rect 10980 30734 11008 36178
rect 11716 35222 11744 36722
rect 12256 36168 12308 36174
rect 12256 36110 12308 36116
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11704 35216 11756 35222
rect 11704 35158 11756 35164
rect 11152 34672 11204 34678
rect 11152 34614 11204 34620
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10784 30388 10836 30394
rect 10784 30330 10836 30336
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10612 30025 10640 30194
rect 10598 30016 10654 30025
rect 10598 29951 10654 29960
rect 10598 29880 10654 29889
rect 10598 29815 10654 29824
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10612 29578 10640 29815
rect 10600 29572 10652 29578
rect 10600 29514 10652 29520
rect 10704 29458 10732 30330
rect 10796 29889 10824 30330
rect 10782 29880 10838 29889
rect 10782 29815 10838 29824
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 10782 29608 10838 29617
rect 10782 29543 10784 29552
rect 10836 29543 10838 29552
rect 10784 29514 10836 29520
rect 10612 29430 10732 29458
rect 10506 28792 10562 28801
rect 10428 28750 10506 28778
rect 10506 28727 10562 28736
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10048 27600 10100 27606
rect 10048 27542 10100 27548
rect 10152 27418 10180 28018
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 9968 27390 10180 27418
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9876 26382 9904 26794
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9770 26208 9826 26217
rect 9770 26143 9826 26152
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9508 25294 9536 25434
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 9586 25120 9642 25129
rect 9508 24410 9536 25094
rect 9586 25055 9642 25064
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9126 21448 9182 21457
rect 9126 21383 9182 21392
rect 9140 21078 9168 21383
rect 9310 21312 9366 21321
rect 9310 21247 9366 21256
rect 9128 21072 9180 21078
rect 9128 21014 9180 21020
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9232 20641 9260 20810
rect 9034 20632 9090 20641
rect 9218 20632 9274 20641
rect 9090 20590 9168 20618
rect 9034 20567 9090 20576
rect 9140 19904 9168 20590
rect 9218 20567 9274 20576
rect 9232 20466 9260 20567
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9220 19916 9272 19922
rect 9140 19876 9220 19904
rect 9220 19858 9272 19864
rect 9036 19780 9088 19786
rect 9324 19768 9352 21247
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9416 19786 9444 20470
rect 9508 19825 9536 23462
rect 9600 22710 9628 25055
rect 9862 24984 9918 24993
rect 9862 24919 9918 24928
rect 9678 24032 9734 24041
rect 9678 23967 9734 23976
rect 9588 22704 9640 22710
rect 9588 22646 9640 22652
rect 9692 22098 9720 23967
rect 9770 23080 9826 23089
rect 9770 23015 9826 23024
rect 9784 22982 9812 23015
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9784 21468 9812 22646
rect 9646 21440 9812 21468
rect 9646 21400 9674 21440
rect 9600 21372 9674 21400
rect 9600 19961 9628 21372
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9678 20360 9734 20369
rect 9678 20295 9734 20304
rect 9586 19952 9642 19961
rect 9586 19887 9642 19896
rect 9494 19816 9550 19825
rect 9088 19740 9352 19768
rect 9404 19780 9456 19786
rect 9036 19722 9088 19728
rect 9494 19751 9550 19760
rect 9404 19722 9456 19728
rect 9048 19417 9076 19722
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 19446 9536 19654
rect 9496 19440 9548 19446
rect 9034 19408 9090 19417
rect 9496 19382 9548 19388
rect 9034 19343 9090 19352
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 9048 17921 9076 19246
rect 9508 19009 9536 19382
rect 9692 19310 9720 20295
rect 9680 19304 9732 19310
rect 9586 19272 9642 19281
rect 9680 19246 9732 19252
rect 9586 19207 9642 19216
rect 9494 19000 9550 19009
rect 9494 18935 9550 18944
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9232 18601 9260 18702
rect 9218 18592 9274 18601
rect 9218 18527 9274 18536
rect 9600 18272 9628 19207
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9508 18244 9628 18272
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9317 18193 9444 18204
rect 9317 18184 9458 18193
rect 9317 18176 9402 18184
rect 9034 17912 9090 17921
rect 9034 17847 9090 17856
rect 9232 17762 9260 18158
rect 9317 17954 9345 18176
rect 9402 18119 9458 18128
rect 9317 17926 9444 17954
rect 9416 17814 9444 17926
rect 9404 17808 9456 17814
rect 9048 17734 9352 17762
rect 9404 17750 9456 17756
rect 9048 17270 9076 17734
rect 9324 17660 9352 17734
rect 9404 17672 9456 17678
rect 9324 17632 9404 17660
rect 9404 17614 9456 17620
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9140 16697 9168 17206
rect 9126 16688 9182 16697
rect 9126 16623 9182 16632
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12850 8984 13262
rect 9048 13258 9076 16458
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9232 13705 9260 15574
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9218 13696 9274 13705
rect 9218 13631 9274 13640
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9218 13288 9274 13297
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8956 10169 8984 12786
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9048 12374 9076 12650
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 8942 10160 8998 10169
rect 8942 10095 8998 10104
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8850 4992 8906 5001
rect 8850 4927 8906 4936
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8864 4706 8892 4927
rect 8956 4826 8984 9687
rect 9048 7585 9076 11766
rect 9140 11694 9168 13262
rect 9218 13223 9274 13232
rect 9232 12238 9260 13223
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9324 11898 9352 13806
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11218 9168 11630
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9140 10606 9168 11154
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9324 10742 9352 10950
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9140 10130 9168 10542
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9140 9586 9168 10066
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9310 9480 9366 9489
rect 9128 9444 9180 9450
rect 9310 9415 9366 9424
rect 9128 9386 9180 9392
rect 9140 8498 9168 9386
rect 9324 8906 9352 9415
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9140 7886 9168 8434
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9034 7576 9090 7585
rect 9034 7511 9090 7520
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9048 6769 9076 6938
rect 9140 6934 9168 7822
rect 9232 7750 9260 8570
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9128 6928 9180 6934
rect 9128 6870 9180 6876
rect 9034 6760 9090 6769
rect 9140 6730 9168 6870
rect 9034 6695 9090 6704
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9232 6662 9260 7346
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6798 9352 7278
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9220 6656 9272 6662
rect 9126 6624 9182 6633
rect 9220 6598 9272 6604
rect 9126 6559 9182 6568
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8864 4678 8984 4706
rect 8588 4644 8708 4672
rect 8680 4570 8708 4644
rect 8956 4622 8984 4678
rect 8944 4616 8996 4622
rect 8680 4542 8892 4570
rect 8944 4558 8996 4564
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8206 4312 8262 4321
rect 8206 4247 8262 4256
rect 8220 4214 8248 4247
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8206 3224 8262 3233
rect 8206 3159 8262 3168
rect 8220 3126 8248 3159
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8024 1488 8076 1494
rect 8024 1430 8076 1436
rect 8128 814 8156 2246
rect 8220 1358 8248 2790
rect 8312 1737 8340 3470
rect 8404 2854 8432 4422
rect 8482 4040 8538 4049
rect 8864 4010 8892 4542
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4214 8984 4422
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 9048 4049 9076 5850
rect 9140 5794 9168 6559
rect 9324 6361 9352 6734
rect 9310 6352 9366 6361
rect 9310 6287 9366 6296
rect 9416 5914 9444 17206
rect 9508 16289 9536 18244
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17377 9628 18022
rect 9586 17368 9642 17377
rect 9586 17303 9642 17312
rect 9494 16280 9550 16289
rect 9494 16215 9550 16224
rect 9600 16182 9628 17303
rect 9692 16658 9720 18702
rect 9784 18340 9812 20742
rect 9876 19310 9904 24919
rect 9968 23769 9996 27390
rect 10230 26888 10286 26897
rect 10230 26823 10286 26832
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 10060 24138 10088 26522
rect 10140 26444 10192 26450
rect 10140 26386 10192 26392
rect 10152 25974 10180 26386
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 10046 23896 10102 23905
rect 10046 23831 10102 23840
rect 9954 23760 10010 23769
rect 9954 23695 10010 23704
rect 10060 22710 10088 23831
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9968 21622 9996 22578
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10060 21729 10088 22034
rect 10046 21720 10102 21729
rect 10046 21655 10102 21664
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9968 20806 9996 21422
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9968 19417 9996 20334
rect 9954 19408 10010 19417
rect 9954 19343 10010 19352
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9876 18601 9904 18838
rect 9862 18592 9918 18601
rect 9968 18578 9996 19178
rect 10060 18698 10088 20742
rect 10152 19446 10180 25638
rect 10244 25362 10272 26823
rect 10336 25838 10364 27542
rect 10324 25832 10376 25838
rect 10324 25774 10376 25780
rect 10232 25356 10284 25362
rect 10232 25298 10284 25304
rect 10244 24041 10272 25298
rect 10230 24032 10286 24041
rect 10230 23967 10286 23976
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10244 22642 10272 23802
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10244 21554 10272 22578
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10336 21010 10364 25774
rect 10428 21078 10456 28358
rect 10520 22166 10548 28727
rect 10612 24818 10640 29430
rect 10784 29096 10836 29102
rect 10784 29038 10836 29044
rect 10796 28529 10824 29038
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10782 28520 10838 28529
rect 10782 28455 10838 28464
rect 10692 27872 10744 27878
rect 10692 27814 10744 27820
rect 10704 27713 10732 27814
rect 10690 27704 10746 27713
rect 10690 27639 10746 27648
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10704 26314 10732 26726
rect 10796 26450 10824 28455
rect 10888 27062 10916 28562
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 10980 27878 11008 28154
rect 10968 27872 11020 27878
rect 10968 27814 11020 27820
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 10980 27402 11008 27542
rect 11072 27538 11100 29650
rect 11164 28150 11192 34614
rect 11900 34202 11928 35634
rect 11888 34196 11940 34202
rect 11888 34138 11940 34144
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11716 30802 11744 31622
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 11072 27334 11100 27474
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11256 27130 11284 30534
rect 12084 30433 12112 31282
rect 12268 30938 12296 36110
rect 13004 35834 13032 37198
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 12992 35828 13044 35834
rect 12992 35770 13044 35776
rect 13360 34944 13412 34950
rect 13360 34886 13412 34892
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12256 30932 12308 30938
rect 12256 30874 12308 30880
rect 12070 30424 12126 30433
rect 12070 30359 12126 30368
rect 11886 30288 11942 30297
rect 11886 30223 11888 30232
rect 11940 30223 11942 30232
rect 12256 30252 12308 30258
rect 11888 30194 11940 30200
rect 12256 30194 12308 30200
rect 12268 30161 12296 30194
rect 12254 30152 12310 30161
rect 12254 30087 12310 30096
rect 11704 30048 11756 30054
rect 11704 29990 11756 29996
rect 11716 29782 11744 29990
rect 11704 29776 11756 29782
rect 11704 29718 11756 29724
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11808 29306 11836 29718
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 12162 29200 12218 29209
rect 12268 29186 12296 30087
rect 12452 29714 12480 31214
rect 12544 30666 12572 33934
rect 12716 30864 12768 30870
rect 12716 30806 12768 30812
rect 12532 30660 12584 30666
rect 12532 30602 12584 30608
rect 12624 30388 12676 30394
rect 12624 30330 12676 30336
rect 12636 30054 12664 30330
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12440 29708 12492 29714
rect 12440 29650 12492 29656
rect 12544 29560 12572 29990
rect 12624 29572 12676 29578
rect 12544 29532 12624 29560
rect 12624 29514 12676 29520
rect 12218 29158 12296 29186
rect 12162 29135 12218 29144
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11244 27124 11296 27130
rect 11296 27084 11376 27112
rect 11244 27066 11296 27072
rect 10876 27056 10928 27062
rect 10876 26998 10928 27004
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 10980 26489 11008 26930
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 10966 26480 11022 26489
rect 10784 26444 10836 26450
rect 10966 26415 11022 26424
rect 10784 26386 10836 26392
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 10508 22160 10560 22166
rect 10508 22102 10560 22108
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10520 21865 10548 21966
rect 10506 21856 10562 21865
rect 10506 21791 10562 21800
rect 10520 21593 10548 21791
rect 10704 21593 10732 23734
rect 10782 23352 10838 23361
rect 10782 23287 10838 23296
rect 10506 21584 10562 21593
rect 10690 21584 10746 21593
rect 10506 21519 10562 21528
rect 10600 21548 10652 21554
rect 10690 21519 10746 21528
rect 10600 21490 10652 21496
rect 10508 21412 10560 21418
rect 10508 21354 10560 21360
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10324 20868 10376 20874
rect 10324 20810 10376 20816
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10244 19922 10272 20538
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10230 19816 10286 19825
rect 10230 19751 10286 19760
rect 10244 19446 10272 19751
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10138 18864 10194 18873
rect 10138 18799 10194 18808
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9968 18550 10088 18578
rect 9862 18527 9918 18536
rect 9784 18312 9996 18340
rect 9968 18136 9996 18312
rect 9777 18108 9996 18136
rect 9777 18068 9805 18108
rect 10060 18068 10088 18550
rect 10152 18358 10180 18799
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 9771 18040 9805 18068
rect 9968 18040 10088 18068
rect 9771 17954 9799 18040
rect 9771 17926 9812 17954
rect 9784 17610 9812 17926
rect 9968 17746 9996 18040
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9508 15434 9536 16050
rect 9692 15570 9720 16594
rect 9784 16522 9812 17546
rect 9862 17096 9918 17105
rect 9862 17031 9918 17040
rect 9876 16794 9904 17031
rect 10140 16992 10192 16998
rect 9968 16952 10140 16980
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9968 15586 9996 16952
rect 10140 16934 10192 16940
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10152 16114 10180 16458
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9784 15558 9996 15586
rect 10060 15570 10088 16050
rect 10048 15564 10100 15570
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9680 15360 9732 15366
rect 9678 15328 9680 15337
rect 9732 15328 9734 15337
rect 9678 15263 9734 15272
rect 9586 15192 9642 15201
rect 9586 15127 9642 15136
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 9508 13297 9536 15030
rect 9600 14346 9628 15127
rect 9784 14770 9812 15558
rect 10048 15506 10100 15512
rect 10048 15428 10100 15434
rect 10048 15370 10100 15376
rect 10060 15337 10088 15370
rect 10046 15328 10102 15337
rect 10046 15263 10102 15272
rect 9862 15192 9918 15201
rect 9862 15127 9918 15136
rect 9876 14958 9904 15127
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9692 14742 9812 14770
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9494 13288 9550 13297
rect 9494 13223 9550 13232
rect 9496 12912 9548 12918
rect 9494 12880 9496 12889
rect 9548 12880 9550 12889
rect 9494 12815 9550 12824
rect 9692 12434 9720 14742
rect 9968 14482 9996 14758
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 12434 9904 14010
rect 10046 13968 10102 13977
rect 10046 13903 10102 13912
rect 10060 13870 10088 13903
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9692 12406 9812 12434
rect 9876 12406 9996 12434
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 9042 9536 10950
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9508 6633 9536 8842
rect 9494 6624 9550 6633
rect 9494 6559 9550 6568
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9140 5766 9352 5794
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9034 4040 9090 4049
rect 8482 3975 8538 3984
rect 8852 4004 8904 4010
rect 8496 3738 8524 3975
rect 9034 3975 9090 3984
rect 8852 3946 8904 3952
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 9034 3632 9090 3641
rect 9034 3567 9090 3576
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8390 2000 8446 2009
rect 8390 1935 8446 1944
rect 8298 1728 8354 1737
rect 8298 1663 8354 1672
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8116 808 8168 814
rect 3568 776 3570 785
rect 3514 711 3570 720
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 5814 200 5870 800
rect 7102 200 7158 800
rect 7746 200 7802 800
rect 8404 800 8432 1935
rect 9048 1358 9076 3567
rect 9140 3534 9168 5646
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9232 3942 9260 5170
rect 9324 4282 9352 5766
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 4826 9444 5306
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9218 3632 9274 3641
rect 9416 3602 9444 3878
rect 9508 3738 9536 6258
rect 9600 5370 9628 12174
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11354 9720 12106
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9692 11150 9720 11290
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 10577 9720 10678
rect 9678 10568 9734 10577
rect 9678 10503 9734 10512
rect 9678 8120 9734 8129
rect 9678 8055 9734 8064
rect 9692 7818 9720 8055
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7177 9720 7754
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9680 6792 9732 6798
rect 9784 6780 9812 12406
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 8129 9904 8230
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 9732 6752 9812 6780
rect 9680 6734 9732 6740
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9692 6118 9720 6326
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4282 9628 5170
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9770 4992 9826 5001
rect 9692 4865 9720 4966
rect 9770 4927 9826 4936
rect 9678 4856 9734 4865
rect 9678 4791 9734 4800
rect 9784 4554 9812 4927
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9692 3670 9720 4490
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9218 3567 9274 3576
rect 9404 3596 9456 3602
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9232 2446 9260 3567
rect 9404 3538 9456 3544
rect 9416 3058 9444 3538
rect 9678 3496 9734 3505
rect 9772 3460 9824 3466
rect 9734 3440 9772 3448
rect 9678 3431 9772 3440
rect 9692 3420 9772 3431
rect 9692 3058 9720 3420
rect 9772 3402 9824 3408
rect 9876 3194 9904 7414
rect 9968 6662 9996 12406
rect 10152 12170 10180 16050
rect 10336 14278 10364 20810
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10324 14272 10376 14278
rect 10244 14220 10324 14226
rect 10244 14214 10376 14220
rect 10244 14198 10364 14214
rect 10244 12238 10272 14198
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10138 11656 10194 11665
rect 10138 11591 10194 11600
rect 10152 11286 10180 11591
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10060 9489 10088 10542
rect 10244 9518 10272 12038
rect 10140 9512 10192 9518
rect 10046 9480 10102 9489
rect 10140 9454 10192 9460
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10046 9415 10102 9424
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9956 6656 10008 6662
rect 10060 6633 10088 8502
rect 10152 8294 10180 9454
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 9956 6598 10008 6604
rect 10046 6624 10102 6633
rect 10046 6559 10102 6568
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 5710 10088 6394
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9968 5302 9996 5646
rect 10046 5400 10102 5409
rect 10046 5335 10048 5344
rect 10100 5335 10102 5344
rect 10048 5306 10100 5312
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9968 4214 9996 4558
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 10060 3466 10088 5170
rect 10152 4010 10180 7754
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10244 3942 10272 7482
rect 10336 5914 10364 13738
rect 10428 11014 10456 19246
rect 10520 17610 10548 21354
rect 10612 20942 10640 21490
rect 10690 21448 10746 21457
rect 10690 21383 10746 21392
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10598 19952 10654 19961
rect 10598 19887 10654 19896
rect 10612 19854 10640 19887
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10600 19440 10652 19446
rect 10600 19382 10652 19388
rect 10612 17762 10640 19382
rect 10704 19224 10732 21383
rect 10796 20534 10824 23287
rect 10888 21457 10916 25162
rect 11072 24721 11100 26726
rect 11242 26072 11298 26081
rect 11242 26007 11298 26016
rect 11150 25528 11206 25537
rect 11150 25463 11206 25472
rect 11058 24712 11114 24721
rect 11058 24647 11114 24656
rect 11058 24576 11114 24585
rect 11058 24511 11114 24520
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 10980 23662 11008 24210
rect 11072 24070 11100 24511
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10980 23118 11008 23598
rect 11072 23497 11100 23666
rect 11058 23488 11114 23497
rect 11058 23423 11114 23432
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 10980 22778 11008 23054
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10980 22574 11008 22714
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 22030 11008 22510
rect 11164 22234 11192 25463
rect 11256 24886 11284 26007
rect 11348 25974 11376 27084
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 11244 24880 11296 24886
rect 11244 24822 11296 24828
rect 11348 24750 11376 25230
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11348 24274 11376 24686
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11440 24154 11468 27950
rect 11348 24126 11468 24154
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11256 23361 11284 24006
rect 11242 23352 11298 23361
rect 11242 23287 11298 23296
rect 11256 23186 11284 23287
rect 11348 23186 11376 24126
rect 11532 23594 11560 28494
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11428 23588 11480 23594
rect 11428 23530 11480 23536
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 11256 22778 11284 22986
rect 11244 22772 11296 22778
rect 11244 22714 11296 22720
rect 11242 22536 11298 22545
rect 11242 22471 11298 22480
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 11058 21992 11114 22001
rect 10874 21448 10930 21457
rect 10874 21383 10930 21392
rect 10874 21040 10930 21049
rect 10874 20975 10930 20984
rect 10888 20806 10916 20975
rect 10980 20942 11008 21966
rect 11058 21927 11114 21936
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10784 20528 10836 20534
rect 10784 20470 10836 20476
rect 10980 20398 11008 20878
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 19916 10928 19922
rect 10980 19904 11008 20334
rect 10928 19876 11008 19904
rect 10876 19858 10928 19864
rect 10876 19780 10928 19786
rect 10928 19740 11008 19768
rect 10876 19722 10928 19728
rect 10874 19348 10930 19357
rect 10874 19283 10930 19292
rect 10784 19236 10836 19242
rect 10704 19196 10784 19224
rect 10784 19178 10836 19184
rect 10612 17734 10732 17762
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10612 17202 10640 17614
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10520 16250 10548 16458
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 14550 10548 14826
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10612 14482 10640 14894
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 14006 10548 14214
rect 10598 14104 10654 14113
rect 10598 14039 10654 14048
rect 10612 14006 10640 14039
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10506 13832 10562 13841
rect 10506 13767 10562 13776
rect 10520 12628 10548 13767
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10612 12782 10640 13398
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10520 12600 10640 12628
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10520 10713 10548 11698
rect 10506 10704 10562 10713
rect 10506 10639 10562 10648
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10428 7041 10456 9590
rect 10520 7410 10548 10134
rect 10612 8974 10640 12600
rect 10704 9042 10732 17734
rect 10796 17377 10824 19178
rect 10888 18222 10916 19283
rect 10876 18216 10928 18222
rect 10980 18193 11008 19740
rect 11072 19009 11100 21927
rect 11164 20874 11192 22170
rect 11256 21690 11284 22471
rect 11440 22409 11468 23530
rect 11624 22982 11652 25162
rect 11704 24880 11756 24886
rect 11704 24822 11756 24828
rect 11716 24449 11744 24822
rect 11702 24440 11758 24449
rect 11702 24375 11758 24384
rect 11704 24132 11756 24138
rect 11704 24074 11756 24080
rect 11716 23866 11744 24074
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11518 22672 11574 22681
rect 11518 22607 11574 22616
rect 11426 22400 11482 22409
rect 11426 22335 11482 22344
rect 11334 21992 11390 22001
rect 11334 21927 11390 21936
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11242 21448 11298 21457
rect 11242 21383 11298 21392
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 11256 19786 11284 21383
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11348 19553 11376 21927
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11334 19544 11390 19553
rect 11244 19508 11296 19514
rect 11334 19479 11390 19488
rect 11244 19450 11296 19456
rect 11256 19378 11284 19450
rect 11334 19408 11390 19417
rect 11244 19372 11296 19378
rect 11334 19343 11390 19352
rect 11244 19314 11296 19320
rect 11150 19272 11206 19281
rect 11150 19207 11206 19216
rect 11058 19000 11114 19009
rect 11058 18935 11114 18944
rect 11164 18834 11192 19207
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 10876 18158 10928 18164
rect 10966 18184 11022 18193
rect 10966 18119 11022 18128
rect 11256 18086 11284 19110
rect 11244 18080 11296 18086
rect 11164 18040 11244 18068
rect 10874 17912 10930 17921
rect 10874 17847 10930 17856
rect 10782 17368 10838 17377
rect 10782 17303 10838 17312
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10796 16522 10824 17070
rect 10888 16522 10916 17847
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 10796 16289 10824 16458
rect 10782 16280 10838 16289
rect 10782 16215 10838 16224
rect 10980 16182 11008 17138
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11072 16046 11100 16118
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10980 15201 11008 15914
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10966 15192 11022 15201
rect 11072 15162 11100 15506
rect 11164 15366 11192 18040
rect 11244 18022 11296 18028
rect 11242 17912 11298 17921
rect 11242 17847 11298 17856
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 10966 15127 11022 15136
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11256 15042 11284 17847
rect 11348 16182 11376 19343
rect 11440 18630 11468 20742
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11440 17134 11468 17274
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11532 16266 11560 22607
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11624 21962 11652 22034
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11624 21690 11652 21898
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11716 21026 11744 23802
rect 11808 21486 11836 26250
rect 11900 22001 11928 27406
rect 11978 26480 12034 26489
rect 11978 26415 11980 26424
rect 12032 26415 12034 26424
rect 11980 26386 12032 26392
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 12084 23798 12112 24074
rect 12176 23882 12204 29135
rect 12728 29102 12756 30806
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 12716 29096 12768 29102
rect 12544 29056 12716 29084
rect 12544 28914 12572 29056
rect 12716 29038 12768 29044
rect 12452 28886 12572 28914
rect 12348 28484 12400 28490
rect 12452 28472 12480 28886
rect 12530 28792 12586 28801
rect 12530 28727 12586 28736
rect 12400 28444 12480 28472
rect 12348 28426 12400 28432
rect 12544 28422 12572 28727
rect 12532 28416 12584 28422
rect 12532 28358 12584 28364
rect 12438 28112 12494 28121
rect 12438 28047 12440 28056
rect 12492 28047 12494 28056
rect 12624 28076 12676 28082
rect 12440 28018 12492 28024
rect 12624 28018 12676 28024
rect 12636 27962 12664 28018
rect 12452 27934 12664 27962
rect 12452 27146 12480 27934
rect 12820 27826 12848 30602
rect 12912 29714 12940 30670
rect 13372 30326 13400 34886
rect 15028 30734 15056 37062
rect 15212 36922 15240 37198
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15488 36854 15516 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 16500 37210 16528 39222
rect 17406 39200 17462 39800
rect 18050 39200 18106 39800
rect 19338 39200 19394 39800
rect 19982 39200 20038 39800
rect 20626 39200 20682 39800
rect 21914 39200 21970 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25134 39200 25190 39800
rect 26422 39200 26478 39800
rect 27066 39200 27122 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 31574 39200 31630 39800
rect 32218 39200 32274 39800
rect 33506 39200 33562 39800
rect 34150 39200 34206 39800
rect 35438 39200 35494 39800
rect 35544 39222 35848 39250
rect 16764 37460 16816 37466
rect 16764 37402 16816 37408
rect 16500 37194 16620 37210
rect 16120 37188 16172 37194
rect 16500 37188 16632 37194
rect 16500 37182 16580 37188
rect 16120 37130 16172 37136
rect 16580 37130 16632 37136
rect 15476 36848 15528 36854
rect 15476 36790 15528 36796
rect 15844 36644 15896 36650
rect 15844 36586 15896 36592
rect 15856 36378 15884 36586
rect 15844 36372 15896 36378
rect 15844 36314 15896 36320
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15384 30660 15436 30666
rect 15384 30602 15436 30608
rect 13360 30320 13412 30326
rect 13360 30262 13412 30268
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 14384 29850 14412 30126
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 13912 29776 13964 29782
rect 13912 29718 13964 29724
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 12544 27798 12848 27826
rect 12544 27402 12572 27798
rect 12716 27532 12768 27538
rect 12912 27520 12940 29650
rect 13082 29336 13138 29345
rect 13082 29271 13138 29280
rect 13096 29034 13124 29271
rect 13924 29102 13952 29718
rect 14752 29646 14780 29990
rect 14556 29640 14608 29646
rect 14384 29588 14556 29594
rect 14384 29582 14608 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14384 29566 14596 29582
rect 14292 29306 14320 29514
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14384 29170 14412 29566
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 13636 29096 13688 29102
rect 13464 29056 13636 29084
rect 13084 29028 13136 29034
rect 13084 28970 13136 28976
rect 13358 28520 13414 28529
rect 13358 28455 13360 28464
rect 13412 28455 13414 28464
rect 13360 28426 13412 28432
rect 13096 27934 13308 27962
rect 13096 27878 13124 27934
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 13176 27872 13228 27878
rect 13176 27814 13228 27820
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 12716 27474 12768 27480
rect 12820 27492 12940 27520
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12452 27118 12572 27146
rect 12728 27130 12756 27474
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 12452 26926 12480 26998
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12256 26852 12308 26858
rect 12256 26794 12308 26800
rect 12268 24138 12296 26794
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12452 26314 12480 26454
rect 12544 26314 12572 27118
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12820 26489 12848 27492
rect 13096 27441 13124 27542
rect 13082 27432 13138 27441
rect 12992 27396 13044 27402
rect 13082 27367 13138 27376
rect 12992 27338 13044 27344
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12806 26480 12862 26489
rect 12806 26415 12862 26424
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12452 25158 12480 25978
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12176 23854 12296 23882
rect 12072 23792 12124 23798
rect 12072 23734 12124 23740
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12176 23497 12204 23598
rect 12162 23488 12218 23497
rect 12162 23423 12218 23432
rect 12268 23338 12296 23854
rect 12176 23310 12296 23338
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 11886 21992 11942 22001
rect 11886 21927 11942 21936
rect 11992 21622 12020 23122
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11886 21448 11942 21457
rect 11886 21383 11942 21392
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11624 20998 11744 21026
rect 11624 20330 11652 20998
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11716 20058 11744 20810
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11808 19938 11836 21286
rect 11716 19910 11836 19938
rect 11610 19544 11666 19553
rect 11610 19479 11666 19488
rect 11624 19446 11652 19479
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11440 16238 11560 16266
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15570 11376 15982
rect 11440 15706 11468 16238
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11426 15600 11482 15609
rect 11336 15564 11388 15570
rect 11532 15570 11560 16050
rect 11426 15535 11482 15544
rect 11520 15564 11572 15570
rect 11336 15506 11388 15512
rect 11072 15014 11284 15042
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10796 14521 10824 14554
rect 10782 14512 10838 14521
rect 10782 14447 10838 14456
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10796 12481 10824 12854
rect 10782 12472 10838 12481
rect 10782 12407 10838 12416
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 12102 10824 12310
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10782 11928 10838 11937
rect 10782 11863 10838 11872
rect 10796 11762 10824 11863
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10796 10985 10824 11562
rect 10782 10976 10838 10985
rect 10782 10911 10838 10920
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10796 10577 10824 10610
rect 10782 10568 10838 10577
rect 10782 10503 10838 10512
rect 10888 9738 10916 13194
rect 11072 12889 11100 15014
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 11164 14226 11192 14826
rect 11440 14618 11468 15535
rect 11520 15506 11572 15512
rect 11532 15026 11560 15506
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11532 14482 11560 14962
rect 11624 14890 11652 18226
rect 11716 17921 11744 19910
rect 11900 19836 11928 21383
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 11992 20369 12020 20470
rect 12084 20398 12112 23122
rect 12072 20392 12124 20398
rect 11978 20360 12034 20369
rect 12072 20334 12124 20340
rect 11978 20295 12034 20304
rect 11808 19808 11928 19836
rect 11702 17912 11758 17921
rect 11702 17847 11758 17856
rect 11808 17660 11836 19808
rect 12176 19768 12204 23310
rect 12254 23080 12310 23089
rect 12254 23015 12256 23024
rect 12308 23015 12310 23024
rect 12256 22986 12308 22992
rect 12438 22808 12494 22817
rect 12438 22743 12440 22752
rect 12492 22743 12494 22752
rect 12440 22714 12492 22720
rect 12256 22704 12308 22710
rect 12254 22672 12256 22681
rect 12308 22672 12310 22681
rect 12544 22658 12572 25094
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12636 23497 12664 23598
rect 12622 23488 12678 23497
rect 12622 23423 12678 23432
rect 12254 22607 12310 22616
rect 12452 22630 12572 22658
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12254 22400 12310 22409
rect 12254 22335 12310 22344
rect 12268 21622 12296 22335
rect 12452 21894 12480 22630
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12452 21350 12480 21830
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12346 20904 12402 20913
rect 12346 20839 12402 20848
rect 12360 20448 12388 20839
rect 12452 20788 12480 21082
rect 12544 21049 12572 21286
rect 12530 21040 12586 21049
rect 12530 20975 12586 20984
rect 12532 20936 12584 20942
rect 12530 20904 12532 20913
rect 12584 20904 12586 20913
rect 12530 20839 12586 20848
rect 12532 20800 12584 20806
rect 12452 20760 12532 20788
rect 12532 20742 12584 20748
rect 11900 19740 12204 19768
rect 12268 20420 12388 20448
rect 11900 19334 11928 19740
rect 12268 19446 12296 20420
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12544 20074 12572 20334
rect 12360 20046 12572 20074
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 11900 19306 12204 19334
rect 11886 19136 11942 19145
rect 11886 19071 11942 19080
rect 11900 18873 11928 19071
rect 11980 18896 12032 18902
rect 11886 18864 11942 18873
rect 11980 18838 12032 18844
rect 12070 18864 12126 18873
rect 11886 18799 11942 18808
rect 11888 18692 11940 18698
rect 11888 18634 11940 18640
rect 11900 18601 11928 18634
rect 11886 18592 11942 18601
rect 11886 18527 11942 18536
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11900 17814 11928 18158
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11808 17632 11928 17660
rect 11796 17536 11848 17542
rect 11702 17504 11758 17513
rect 11796 17478 11848 17484
rect 11702 17439 11758 17448
rect 11716 17338 11744 17439
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11808 17241 11836 17478
rect 11794 17232 11850 17241
rect 11794 17167 11850 17176
rect 11794 15736 11850 15745
rect 11794 15671 11850 15680
rect 11808 15434 11836 15671
rect 11900 15434 11928 17632
rect 11992 17270 12020 18838
rect 12070 18799 12126 18808
rect 12084 18465 12112 18799
rect 12070 18456 12126 18465
rect 12070 18391 12126 18400
rect 12176 18204 12204 19306
rect 12360 18986 12388 20046
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12452 19700 12480 19926
rect 12544 19825 12572 19926
rect 12530 19816 12586 19825
rect 12530 19751 12586 19760
rect 12532 19712 12584 19718
rect 12452 19672 12532 19700
rect 12532 19654 12584 19660
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 19310 12480 19382
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12268 18958 12388 18986
rect 12268 18902 12296 18958
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12544 18834 12572 19178
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12346 18456 12402 18465
rect 12346 18391 12348 18400
rect 12400 18391 12402 18400
rect 12348 18362 12400 18368
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12176 18176 12296 18204
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 12084 17513 12112 18090
rect 12268 17898 12296 18176
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17921 12480 18022
rect 12438 17912 12494 17921
rect 12268 17870 12388 17898
rect 12162 17640 12218 17649
rect 12162 17575 12164 17584
rect 12216 17575 12218 17584
rect 12164 17546 12216 17552
rect 12256 17536 12308 17542
rect 12070 17504 12126 17513
rect 12256 17478 12308 17484
rect 12070 17439 12126 17448
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 12072 16992 12124 16998
rect 12268 16969 12296 17478
rect 12072 16934 12124 16940
rect 12254 16960 12310 16969
rect 11992 16726 12020 16934
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 12084 16425 12112 16934
rect 12254 16895 12310 16904
rect 12162 16688 12218 16697
rect 12162 16623 12218 16632
rect 12176 16522 12204 16623
rect 12360 16590 12388 17870
rect 12438 17847 12494 17856
rect 12544 17678 12572 18294
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12636 17592 12664 22646
rect 12728 22273 12756 26318
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12820 22778 12848 25774
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12806 22400 12862 22409
rect 12806 22335 12862 22344
rect 12714 22264 12770 22273
rect 12714 22199 12770 22208
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12728 20874 12756 21966
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 19786 12756 19858
rect 12716 19780 12768 19786
rect 12716 19722 12768 19728
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12728 17660 12756 18158
rect 12820 17954 12848 22335
rect 12912 21486 12940 26862
rect 13004 24857 13032 27338
rect 13188 27316 13216 27814
rect 13096 27288 13216 27316
rect 12990 24848 13046 24857
rect 12990 24783 13046 24792
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13004 21486 13032 24550
rect 13096 21876 13124 27288
rect 13176 27056 13228 27062
rect 13176 26998 13228 27004
rect 13188 22574 13216 26998
rect 13280 26926 13308 27934
rect 13464 27033 13492 29056
rect 13636 29038 13688 29044
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 13820 28960 13872 28966
rect 13820 28902 13872 28908
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 13450 27024 13506 27033
rect 13372 26994 13450 27010
rect 13360 26988 13450 26994
rect 13412 26982 13450 26988
rect 13450 26959 13506 26968
rect 13544 26988 13596 26994
rect 13360 26930 13412 26936
rect 13268 26920 13320 26926
rect 13464 26899 13492 26959
rect 13544 26930 13596 26936
rect 13268 26862 13320 26868
rect 13452 26784 13504 26790
rect 13556 26761 13584 26930
rect 13648 26897 13676 27950
rect 13634 26888 13690 26897
rect 13634 26823 13690 26832
rect 13740 26772 13768 28426
rect 13832 28150 13860 28902
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13924 27996 13952 29038
rect 14188 28076 14240 28082
rect 13452 26726 13504 26732
rect 13542 26752 13598 26761
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 13280 26314 13308 26386
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 13360 25696 13412 25702
rect 13360 25638 13412 25644
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 13280 24410 13308 24618
rect 13268 24404 13320 24410
rect 13268 24346 13320 24352
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13280 23186 13308 24074
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13266 23080 13322 23089
rect 13266 23015 13322 23024
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13174 22128 13230 22137
rect 13174 22063 13176 22072
rect 13228 22063 13230 22072
rect 13176 22034 13228 22040
rect 13176 21888 13228 21894
rect 13096 21848 13176 21876
rect 13176 21830 13228 21836
rect 13082 21584 13138 21593
rect 13082 21519 13138 21528
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 12912 20602 12940 21422
rect 12990 21312 13046 21321
rect 12990 21247 13046 21256
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12912 19825 12940 19994
rect 12898 19816 12954 19825
rect 12898 19751 12954 19760
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18873 12940 19110
rect 12898 18864 12954 18873
rect 12898 18799 12954 18808
rect 13004 18222 13032 21247
rect 13096 20806 13124 21519
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13082 19952 13138 19961
rect 13082 19887 13138 19896
rect 13096 19378 13124 19887
rect 13188 19514 13216 21830
rect 13280 19938 13308 23015
rect 13372 20534 13400 25638
rect 13464 23798 13492 26726
rect 13542 26687 13598 26696
rect 13648 26744 13768 26772
rect 13832 27968 13952 27996
rect 14016 28036 14188 28064
rect 13648 25770 13676 26744
rect 13832 26314 13860 27968
rect 14016 27946 14044 28036
rect 14188 28018 14240 28024
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 14016 26518 14044 27474
rect 14280 27396 14332 27402
rect 14280 27338 14332 27344
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14292 27282 14320 27338
rect 14004 26512 14056 26518
rect 14004 26454 14056 26460
rect 13820 26308 13872 26314
rect 13820 26250 13872 26256
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13636 25764 13688 25770
rect 13636 25706 13688 25712
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13464 20534 13492 23530
rect 13556 23361 13584 25230
rect 13636 25152 13688 25158
rect 13636 25094 13688 25100
rect 13542 23352 13598 23361
rect 13542 23287 13598 23296
rect 13648 23050 13676 25094
rect 13740 24886 13768 25774
rect 13832 25158 13860 26250
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 13924 25906 13952 26182
rect 14016 25974 14044 26182
rect 14004 25968 14056 25974
rect 14004 25910 14056 25916
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 13912 25764 13964 25770
rect 13912 25706 13964 25712
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13728 24880 13780 24886
rect 13728 24822 13780 24828
rect 13728 24744 13780 24750
rect 13924 24732 13952 25706
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 13780 24704 13952 24732
rect 13728 24686 13780 24692
rect 13740 23633 13768 24686
rect 13910 24440 13966 24449
rect 13910 24375 13966 24384
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13832 23905 13860 24210
rect 13924 24070 13952 24375
rect 14016 24138 14044 25298
rect 14108 24886 14136 27270
rect 14292 27254 14412 27282
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13818 23896 13874 23905
rect 14200 23866 14228 26930
rect 13818 23831 13874 23840
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 13820 23656 13872 23662
rect 13726 23624 13782 23633
rect 13820 23598 13872 23604
rect 13726 23559 13782 23568
rect 13636 23044 13688 23050
rect 13636 22986 13688 22992
rect 13544 22704 13596 22710
rect 13542 22672 13544 22681
rect 13596 22672 13598 22681
rect 13542 22607 13598 22616
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 13360 20528 13412 20534
rect 13360 20470 13412 20476
rect 13452 20528 13504 20534
rect 13556 20505 13584 22510
rect 13832 22030 13860 23598
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 13910 22672 13966 22681
rect 13910 22607 13966 22616
rect 13924 22574 13952 22607
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13832 21593 13860 21966
rect 13818 21584 13874 21593
rect 13818 21519 13874 21528
rect 13726 21448 13782 21457
rect 13726 21383 13782 21392
rect 13912 21412 13964 21418
rect 13740 21078 13768 21383
rect 13912 21354 13964 21360
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13452 20470 13504 20476
rect 13542 20496 13598 20505
rect 13542 20431 13598 20440
rect 13648 20058 13676 20946
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13740 20584 13768 20878
rect 13740 20556 13860 20584
rect 13726 20496 13782 20505
rect 13726 20431 13782 20440
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13280 19910 13584 19938
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13084 19372 13136 19378
rect 13136 19320 13216 19334
rect 13084 19314 13216 19320
rect 13096 19306 13216 19314
rect 13188 18698 13216 19306
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13280 18358 13308 19910
rect 13556 19854 13584 19910
rect 13740 19854 13768 20431
rect 13832 20398 13860 20556
rect 13924 20534 13952 21354
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13818 19952 13874 19961
rect 13818 19887 13874 19896
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13372 18873 13400 19722
rect 13464 19514 13492 19722
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13452 19304 13504 19310
rect 13452 19246 13504 19252
rect 13358 18864 13414 18873
rect 13464 18834 13492 19246
rect 13358 18799 13414 18808
rect 13452 18828 13504 18834
rect 13372 18601 13400 18799
rect 13452 18770 13504 18776
rect 13358 18592 13414 18601
rect 13358 18527 13414 18536
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12820 17926 13032 17954
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 12728 17632 12848 17660
rect 12636 17564 12756 17592
rect 12532 17536 12584 17542
rect 12452 17496 12532 17524
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12070 16416 12126 16425
rect 12070 16351 12126 16360
rect 12360 16266 12388 16526
rect 12452 16522 12480 17496
rect 12532 17478 12584 17484
rect 12728 17218 12756 17564
rect 12544 17190 12756 17218
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12268 16238 12388 16266
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11702 15328 11758 15337
rect 11702 15263 11758 15272
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11244 14340 11296 14346
rect 11624 14328 11652 14554
rect 11296 14300 11652 14328
rect 11244 14282 11296 14288
rect 11716 14260 11744 15263
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11794 14648 11850 14657
rect 11794 14583 11850 14592
rect 11532 14232 11744 14260
rect 11164 14198 11376 14226
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11058 12880 11114 12889
rect 11058 12815 11114 12824
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 10674 11008 12718
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11393 11100 11494
rect 11058 11384 11114 11393
rect 11058 11319 11114 11328
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 11072 10198 11100 11018
rect 11164 10713 11192 13466
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11256 12782 11284 12922
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11256 12306 11284 12718
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11256 11762 11284 12242
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11150 10704 11206 10713
rect 11150 10639 11206 10648
rect 11150 10568 11206 10577
rect 11150 10503 11206 10512
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9897 11100 9930
rect 11058 9888 11114 9897
rect 11058 9823 11114 9832
rect 10888 9710 11008 9738
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10874 9072 10930 9081
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10598 8664 10654 8673
rect 10598 8599 10654 8608
rect 10612 7936 10640 8599
rect 10612 7908 10732 7936
rect 10598 7848 10654 7857
rect 10598 7783 10654 7792
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10414 7032 10470 7041
rect 10414 6967 10470 6976
rect 10520 6916 10548 7210
rect 10428 6888 10548 6916
rect 10428 6798 10456 6888
rect 10416 6792 10468 6798
rect 10612 6746 10640 7783
rect 10704 6866 10732 7908
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10416 6734 10468 6740
rect 10520 6718 10640 6746
rect 10692 6724 10744 6730
rect 10414 6624 10470 6633
rect 10414 6559 10470 6568
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10324 5636 10376 5642
rect 10324 5578 10376 5584
rect 10336 5545 10364 5578
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10428 4740 10456 6559
rect 10520 6322 10548 6718
rect 10796 6712 10824 9046
rect 10874 9007 10930 9016
rect 10888 8673 10916 9007
rect 10874 8664 10930 8673
rect 10874 8599 10930 8608
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7478 10916 8230
rect 10980 7818 11008 9710
rect 11164 9704 11192 10503
rect 11072 9676 11192 9704
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 11072 7290 11100 9676
rect 11256 9602 11284 11562
rect 11348 10441 11376 14198
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 13297 11468 13330
rect 11426 13288 11482 13297
rect 11426 13223 11482 13232
rect 11334 10432 11390 10441
rect 11334 10367 11390 10376
rect 11334 10296 11390 10305
rect 11334 10231 11390 10240
rect 11164 9574 11284 9602
rect 11164 9382 11192 9574
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11242 9072 11298 9081
rect 11348 9058 11376 10231
rect 11440 9194 11468 13223
rect 11532 12306 11560 14232
rect 11808 13954 11836 14583
rect 11624 13926 11836 13954
rect 11624 13734 11652 13926
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11624 12889 11652 13359
rect 11716 13326 11744 13806
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11610 12880 11666 12889
rect 11610 12815 11666 12824
rect 11716 12782 11744 13262
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11532 10577 11560 11766
rect 11704 11688 11756 11694
rect 11702 11656 11704 11665
rect 11756 11656 11758 11665
rect 11702 11591 11758 11600
rect 11702 10840 11758 10849
rect 11702 10775 11758 10784
rect 11716 10742 11744 10775
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11518 10296 11574 10305
rect 11518 10231 11574 10240
rect 11532 10198 11560 10231
rect 11520 10192 11572 10198
rect 11716 10146 11744 10474
rect 11520 10134 11572 10140
rect 11624 10118 11744 10146
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9330 11560 9998
rect 11624 9994 11652 10118
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11716 9518 11744 9998
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11532 9302 11652 9330
rect 11440 9166 11560 9194
rect 11348 9030 11468 9058
rect 11242 9007 11244 9016
rect 11296 9007 11298 9016
rect 11244 8978 11296 8984
rect 11336 8492 11388 8498
rect 11164 8452 11336 8480
rect 11164 7410 11192 8452
rect 11336 8434 11388 8440
rect 11334 8392 11390 8401
rect 11334 8327 11390 8336
rect 11348 7954 11376 8327
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11072 7262 11192 7290
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 7041 11100 7142
rect 10874 7032 10930 7041
rect 10874 6967 10930 6976
rect 11058 7032 11114 7041
rect 11058 6967 11114 6976
rect 10744 6684 10824 6712
rect 10692 6666 10744 6672
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6440 10640 6598
rect 10692 6452 10744 6458
rect 10612 6412 10692 6440
rect 10692 6394 10744 6400
rect 10796 6361 10824 6684
rect 10888 6458 10916 6967
rect 11164 6746 11192 7262
rect 10980 6718 11192 6746
rect 10980 6474 11008 6718
rect 11060 6656 11112 6662
rect 11112 6616 11192 6644
rect 11060 6598 11112 6604
rect 10876 6452 10928 6458
rect 10980 6446 11100 6474
rect 10876 6394 10928 6400
rect 10968 6384 11020 6390
rect 10598 6352 10654 6361
rect 10508 6316 10560 6322
rect 10598 6287 10654 6296
rect 10782 6352 10838 6361
rect 10968 6326 11020 6332
rect 10782 6287 10838 6296
rect 10508 6258 10560 6264
rect 10612 4826 10640 6287
rect 10692 6248 10744 6254
rect 10876 6248 10928 6254
rect 10744 6196 10876 6202
rect 10692 6190 10928 6196
rect 10704 6174 10916 6190
rect 10980 6186 11008 6326
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10796 5234 10824 5646
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10704 5030 10732 5170
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10428 4712 10548 4740
rect 10520 4264 10548 4712
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10520 4236 10640 4264
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10232 3528 10284 3534
rect 10336 3505 10364 3878
rect 10520 3534 10548 4082
rect 10612 3738 10640 4236
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10704 3618 10732 4626
rect 10612 3590 10732 3618
rect 10796 3602 10824 5170
rect 10888 5114 10916 5510
rect 11072 5370 11100 6446
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10888 5086 11008 5114
rect 10980 4758 11008 5086
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10784 3596 10836 3602
rect 10508 3528 10560 3534
rect 10232 3470 10284 3476
rect 10322 3496 10378 3505
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 9140 1902 9168 2382
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9692 800 9720 2382
rect 10060 2106 10088 2382
rect 10244 2145 10272 3470
rect 10508 3470 10560 3476
rect 10612 3466 10640 3590
rect 10784 3538 10836 3544
rect 10690 3496 10746 3505
rect 10322 3431 10378 3440
rect 10600 3460 10652 3466
rect 10888 3466 10916 4558
rect 10690 3431 10746 3440
rect 10876 3460 10928 3466
rect 10600 3402 10652 3408
rect 10704 3126 10732 3431
rect 10876 3402 10928 3408
rect 11164 3194 11192 6616
rect 11256 5778 11284 7414
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11242 5672 11298 5681
rect 11242 5607 11244 5616
rect 11296 5607 11298 5616
rect 11244 5578 11296 5584
rect 11242 5264 11298 5273
rect 11242 5199 11298 5208
rect 11256 5098 11284 5199
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11348 3670 11376 7414
rect 11440 4758 11468 9030
rect 11532 8906 11560 9166
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11624 8786 11652 9302
rect 11716 9081 11744 9454
rect 11702 9072 11758 9081
rect 11702 9007 11758 9016
rect 11532 8758 11652 8786
rect 11532 4826 11560 8758
rect 11716 8430 11744 9007
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11716 8090 11744 8366
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11624 7274 11652 7958
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11716 7154 11744 8026
rect 11808 7206 11836 13670
rect 11900 13433 11928 15030
rect 11992 14006 12020 16118
rect 12162 15328 12218 15337
rect 12162 15263 12218 15272
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12084 14929 12112 15030
rect 12070 14920 12126 14929
rect 12070 14855 12126 14864
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11886 13424 11942 13433
rect 11886 13359 11942 13368
rect 12084 13258 12112 14855
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11900 12646 11928 12922
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11900 11218 11928 11698
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11900 10674 11928 11154
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11886 10568 11942 10577
rect 11886 10503 11888 10512
rect 11940 10503 11942 10512
rect 11888 10474 11940 10480
rect 12084 10112 12112 10678
rect 11900 10084 12112 10112
rect 11900 9081 11928 10084
rect 12176 10044 12204 15263
rect 12268 13841 12296 16238
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12452 15881 12480 16118
rect 12438 15872 12494 15881
rect 12438 15807 12494 15816
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12360 14396 12388 15642
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14521 12480 15030
rect 12438 14512 12494 14521
rect 12438 14447 12494 14456
rect 12360 14368 12480 14396
rect 12254 13832 12310 13841
rect 12254 13767 12310 13776
rect 12452 12646 12480 14368
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12544 12434 12572 17190
rect 12820 16674 12848 17632
rect 12912 17513 12940 17750
rect 12898 17504 12954 17513
rect 12898 17439 12954 17448
rect 12898 17368 12954 17377
rect 12898 17303 12954 17312
rect 12636 16646 12848 16674
rect 12636 13394 12664 16646
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12820 15881 12848 16458
rect 12806 15872 12862 15881
rect 12806 15807 12862 15816
rect 12820 15609 12848 15807
rect 12806 15600 12862 15609
rect 12806 15535 12862 15544
rect 12714 14784 12770 14793
rect 12714 14719 12770 14728
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12544 12406 12664 12434
rect 12438 12336 12494 12345
rect 12438 12271 12494 12280
rect 12452 11393 12480 12271
rect 12438 11384 12494 11393
rect 12438 11319 12494 11328
rect 12636 11286 12664 12406
rect 12728 12220 12756 14719
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 12481 12848 14350
rect 12806 12472 12862 12481
rect 12806 12407 12862 12416
rect 12912 12374 12940 17303
rect 13004 14482 13032 17926
rect 13358 17776 13414 17785
rect 13358 17711 13414 17720
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 16590 13124 17614
rect 13372 17134 13400 17711
rect 13360 17128 13412 17134
rect 13266 17096 13322 17105
rect 13360 17070 13412 17076
rect 13266 17031 13322 17040
rect 13280 16697 13308 17031
rect 13266 16688 13322 16697
rect 13266 16623 13322 16632
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13084 15632 13136 15638
rect 13188 15609 13216 15846
rect 13280 15745 13308 15846
rect 13266 15736 13322 15745
rect 13266 15671 13322 15680
rect 13084 15574 13136 15580
rect 13174 15600 13230 15609
rect 13096 15473 13124 15574
rect 13174 15535 13230 15544
rect 13082 15464 13138 15473
rect 13082 15399 13138 15408
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 13372 13954 13400 17070
rect 13464 14958 13492 18294
rect 13556 16250 13584 19382
rect 13648 16522 13676 19654
rect 13740 19417 13768 19654
rect 13832 19446 13860 19887
rect 13924 19786 13952 19994
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 13820 19440 13872 19446
rect 13726 19408 13782 19417
rect 13820 19382 13872 19388
rect 13726 19343 13782 19352
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 18630 13860 18770
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13910 18592 13966 18601
rect 13910 18527 13966 18536
rect 13726 17368 13782 17377
rect 13726 17303 13782 17312
rect 13740 17134 13768 17303
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13924 16697 13952 18527
rect 13910 16688 13966 16697
rect 13910 16623 13966 16632
rect 13924 16590 13952 16623
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13924 16114 13952 16526
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13648 15706 13676 15982
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13740 15201 13768 15982
rect 13726 15192 13782 15201
rect 13726 15127 13782 15136
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13372 13926 13492 13954
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13266 13560 13322 13569
rect 13266 13495 13322 13504
rect 13280 13462 13308 13495
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13176 13388 13228 13394
rect 13096 13348 13176 13376
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 12728 12192 12940 12220
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12268 10849 12296 11222
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12254 10840 12310 10849
rect 12254 10775 12310 10784
rect 12452 10130 12480 11086
rect 12544 11064 12572 11222
rect 12808 11076 12860 11082
rect 12544 11036 12756 11064
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12530 10160 12586 10169
rect 12440 10124 12492 10130
rect 12530 10095 12586 10104
rect 12440 10066 12492 10072
rect 11992 10016 12204 10044
rect 11992 9382 12020 10016
rect 12256 9988 12308 9994
rect 12176 9948 12256 9976
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11886 9072 11942 9081
rect 11886 9007 11942 9016
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 11886 8664 11942 8673
rect 11886 8599 11942 8608
rect 11900 8566 11928 8599
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7750 11928 7890
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 12084 7546 12112 8842
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11624 7126 11744 7154
rect 11796 7200 11848 7206
rect 12176 7154 12204 9948
rect 12256 9930 12308 9936
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12268 7460 12296 9590
rect 12544 9382 12572 10095
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12360 8344 12388 9318
rect 12636 9178 12664 10678
rect 12728 10130 12756 11036
rect 12808 11018 12860 11024
rect 12820 10169 12848 11018
rect 12912 10985 12940 12192
rect 12898 10976 12954 10985
rect 12898 10911 12954 10920
rect 12806 10160 12862 10169
rect 12716 10124 12768 10130
rect 12806 10095 12862 10104
rect 12716 10066 12768 10072
rect 12806 10024 12862 10033
rect 12806 9959 12862 9968
rect 12820 9178 12848 9959
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12544 8566 12572 8910
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 13004 8480 13032 13194
rect 13096 12714 13124 13348
rect 13176 13330 13228 13336
rect 13372 13138 13400 13806
rect 13280 13110 13400 13138
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13096 8974 13124 12310
rect 13188 10198 13216 12786
rect 13280 12345 13308 13110
rect 13464 13002 13492 13926
rect 13372 12974 13492 13002
rect 13372 12850 13400 12974
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13266 12336 13322 12345
rect 13266 12271 13322 12280
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13280 11150 13308 11562
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13280 8634 13308 8978
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8498 13400 12106
rect 13464 11830 13492 12854
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13556 11762 13584 14894
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 13569 13676 14282
rect 13634 13560 13690 13569
rect 13634 13495 13690 13504
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12782 13676 13330
rect 13740 12918 13768 15127
rect 13924 15026 13952 16050
rect 14016 15978 14044 22714
rect 14108 22438 14136 22986
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 21622 14136 22374
rect 14200 22098 14228 23666
rect 14292 22710 14320 27066
rect 14384 26314 14412 27254
rect 14476 26314 14504 29446
rect 14568 27577 14596 29566
rect 14648 29232 14700 29238
rect 14648 29174 14700 29180
rect 14554 27568 14610 27577
rect 14554 27503 14610 27512
rect 14660 27402 14688 29174
rect 14648 27396 14700 27402
rect 14648 27338 14700 27344
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14660 26450 14688 27066
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14752 26058 14780 29582
rect 14936 28490 14964 29990
rect 15396 29850 15424 30602
rect 16132 30394 16160 37130
rect 16120 30388 16172 30394
rect 16120 30330 16172 30336
rect 16304 30252 16356 30258
rect 16304 30194 16356 30200
rect 16316 30161 16344 30194
rect 16488 30184 16540 30190
rect 16302 30152 16358 30161
rect 16488 30126 16540 30132
rect 16302 30087 16358 30096
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 15292 29776 15344 29782
rect 15014 29744 15070 29753
rect 15292 29718 15344 29724
rect 15014 29679 15070 29688
rect 14924 28484 14976 28490
rect 14924 28426 14976 28432
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14476 26030 14780 26058
rect 14476 24800 14504 26030
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 14568 24993 14596 25842
rect 14844 25294 14872 25842
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14554 24984 14610 24993
rect 14554 24919 14610 24928
rect 14476 24772 14780 24800
rect 14646 24712 14702 24721
rect 14646 24647 14702 24656
rect 14660 24410 14688 24647
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 14384 23662 14412 23802
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14372 23248 14424 23254
rect 14372 23190 14424 23196
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14108 19786 14136 21422
rect 14186 21040 14242 21049
rect 14186 20975 14242 20984
rect 14200 20874 14228 20975
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14108 19553 14136 19722
rect 14094 19544 14150 19553
rect 14094 19479 14150 19488
rect 14094 19408 14150 19417
rect 14094 19343 14150 19352
rect 14108 18902 14136 19343
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14200 18222 14228 18634
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14278 18048 14334 18057
rect 14278 17983 14334 17992
rect 14094 17912 14150 17921
rect 14094 17847 14150 17856
rect 14108 17241 14136 17847
rect 14292 17626 14320 17983
rect 14384 17746 14412 23190
rect 14462 23080 14518 23089
rect 14462 23015 14464 23024
rect 14516 23015 14518 23024
rect 14464 22986 14516 22992
rect 14568 22574 14596 23598
rect 14648 22704 14700 22710
rect 14648 22646 14700 22652
rect 14556 22568 14608 22574
rect 14556 22510 14608 22516
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14476 22234 14504 22442
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14462 22128 14518 22137
rect 14462 22063 14518 22072
rect 14476 20874 14504 22063
rect 14464 20868 14516 20874
rect 14464 20810 14516 20816
rect 14462 20768 14518 20777
rect 14462 20703 14518 20712
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14292 17610 14412 17626
rect 14188 17604 14240 17610
rect 14292 17604 14424 17610
rect 14292 17598 14372 17604
rect 14188 17546 14240 17552
rect 14372 17546 14424 17552
rect 14094 17232 14150 17241
rect 14094 17167 14150 17176
rect 14200 16969 14228 17546
rect 14278 17368 14334 17377
rect 14278 17303 14334 17312
rect 14186 16960 14242 16969
rect 14186 16895 14242 16904
rect 14292 16640 14320 17303
rect 14370 17232 14426 17241
rect 14370 17167 14426 17176
rect 14384 16998 14412 17167
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14200 16612 14320 16640
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 14004 15428 14056 15434
rect 14004 15370 14056 15376
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13924 14414 13952 14962
rect 14016 14793 14044 15370
rect 14002 14784 14058 14793
rect 14002 14719 14058 14728
rect 14016 14550 14044 14719
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13818 13832 13874 13841
rect 13818 13767 13874 13776
rect 13832 13394 13860 13767
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 14108 13002 14136 16526
rect 13924 12974 14136 13002
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13740 12594 13768 12650
rect 13648 12566 13768 12594
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13542 11656 13598 11665
rect 13542 11591 13598 11600
rect 13556 11121 13584 11591
rect 13542 11112 13598 11121
rect 13542 11047 13598 11056
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13556 10810 13584 10950
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13450 10160 13506 10169
rect 13450 10095 13506 10104
rect 13544 10124 13596 10130
rect 13360 8492 13412 8498
rect 13004 8452 13124 8480
rect 12992 8356 13044 8362
rect 12360 8316 12992 8344
rect 12992 8298 13044 8304
rect 13096 8072 13124 8452
rect 13360 8434 13412 8440
rect 13372 8344 13400 8434
rect 13188 8316 13400 8344
rect 13188 8090 13216 8316
rect 13266 8256 13322 8265
rect 13266 8191 13322 8200
rect 13004 8044 13124 8072
rect 13176 8084 13228 8090
rect 12900 8016 12952 8022
rect 12898 7984 12900 7993
rect 12952 7984 12954 7993
rect 12898 7919 12954 7928
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 12260 7432 12296 7460
rect 12260 7392 12288 7432
rect 12260 7364 12296 7392
rect 11796 7142 11848 7148
rect 11992 7126 12204 7154
rect 11624 6662 11652 7126
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 6322 11652 6598
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11612 5568 11664 5574
rect 11610 5536 11612 5545
rect 11664 5536 11666 5545
rect 11610 5471 11666 5480
rect 11808 5370 11836 5646
rect 11900 5574 11928 6967
rect 11992 6474 12020 7126
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6644 12112 6938
rect 12084 6633 12204 6644
rect 12084 6624 12218 6633
rect 12084 6616 12162 6624
rect 12162 6559 12218 6568
rect 11992 6446 12112 6474
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11702 5128 11758 5137
rect 11612 5092 11664 5098
rect 11900 5114 11928 5306
rect 11758 5086 11928 5114
rect 11702 5063 11758 5072
rect 11612 5034 11664 5040
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11624 4486 11652 5034
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10230 2136 10286 2145
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10048 2100 10100 2106
rect 10230 2071 10286 2080
rect 10048 2042 10100 2048
rect 9968 1698 9996 2042
rect 9956 1692 10008 1698
rect 9956 1634 10008 1640
rect 10336 800 10364 2994
rect 11440 2990 11468 4150
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 10888 2582 10916 2615
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10980 2417 11008 2450
rect 10966 2408 11022 2417
rect 10966 2343 11022 2352
rect 11164 2310 11192 2926
rect 11716 2922 11744 4966
rect 11796 4820 11848 4826
rect 12084 4808 12112 6446
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12176 5030 12204 6394
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11796 4762 11848 4768
rect 11992 4780 12112 4808
rect 11808 4622 11836 4762
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11992 4146 12020 4780
rect 12070 4720 12126 4729
rect 12268 4706 12296 7364
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12360 5846 12388 7142
rect 12544 6662 12572 7142
rect 12624 6928 12676 6934
rect 12622 6896 12624 6905
rect 12676 6896 12678 6905
rect 12622 6831 12678 6840
rect 12806 6896 12862 6905
rect 12806 6831 12862 6840
rect 12820 6798 12848 6831
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12636 6304 12664 6666
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12452 6276 12664 6304
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12346 5672 12402 5681
rect 12346 5607 12348 5616
rect 12400 5607 12402 5616
rect 12348 5578 12400 5584
rect 12452 4826 12480 6276
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12544 5681 12572 5782
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12530 5672 12586 5681
rect 12636 5658 12664 5714
rect 12820 5710 12848 6598
rect 12808 5704 12860 5710
rect 12636 5630 12756 5658
rect 12808 5646 12860 5652
rect 12530 5607 12586 5616
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12530 5400 12586 5409
rect 12530 5335 12532 5344
rect 12584 5335 12586 5344
rect 12532 5306 12584 5312
rect 12636 5166 12664 5510
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12530 4856 12586 4865
rect 12440 4820 12492 4826
rect 12530 4791 12586 4800
rect 12440 4762 12492 4768
rect 12070 4655 12126 4664
rect 12176 4678 12296 4706
rect 12346 4720 12402 4729
rect 12084 4554 12112 4655
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 12176 4434 12204 4678
rect 12346 4655 12402 4664
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12084 4406 12204 4434
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12084 4010 12112 4406
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12176 4185 12204 4218
rect 12162 4176 12218 4185
rect 12162 4111 12218 4120
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12176 3738 12204 3878
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11624 800 11652 2790
rect 11808 2514 11836 3606
rect 11888 3528 11940 3534
rect 12268 3516 12296 4558
rect 12360 4010 12388 4655
rect 12544 4622 12572 4791
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12452 3942 12480 4082
rect 12544 4049 12572 4150
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12530 3768 12586 3777
rect 12636 3738 12664 5102
rect 12728 4554 12756 5630
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12716 4208 12768 4214
rect 12820 4185 12848 4762
rect 12716 4150 12768 4156
rect 12806 4176 12862 4185
rect 12530 3703 12586 3712
rect 12624 3732 12676 3738
rect 11940 3488 12296 3516
rect 11888 3470 11940 3476
rect 11992 2854 12020 3488
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12452 3058 12480 3402
rect 12544 3108 12572 3703
rect 12624 3674 12676 3680
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12636 3398 12664 3538
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12728 3194 12756 4150
rect 12806 4111 12808 4120
rect 12860 4111 12862 4120
rect 12808 4082 12860 4088
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12544 3080 12664 3108
rect 12636 3074 12664 3080
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12440 3052 12492 3058
rect 12636 3046 12756 3074
rect 12440 2994 12492 3000
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 12360 2564 12388 2994
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12440 2576 12492 2582
rect 12360 2536 12440 2564
rect 12440 2518 12492 2524
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12440 2440 12492 2446
rect 12176 2400 12440 2428
rect 12176 2310 12204 2400
rect 12440 2382 12492 2388
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 800 12296 2246
rect 12544 2038 12572 2450
rect 12636 2446 12664 2926
rect 12728 2922 12756 3046
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12728 2106 12756 2586
rect 12820 2446 12848 4082
rect 12912 3194 12940 7754
rect 13004 4826 13032 8044
rect 13176 8026 13228 8032
rect 13280 7993 13308 8191
rect 13464 8072 13492 10095
rect 13544 10066 13596 10072
rect 13372 8044 13492 8072
rect 13266 7984 13322 7993
rect 13266 7919 13322 7928
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13082 5808 13138 5817
rect 13082 5743 13138 5752
rect 13096 5545 13124 5743
rect 13082 5536 13138 5545
rect 13082 5471 13138 5480
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13004 4010 13032 4558
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 13096 3942 13124 5471
rect 13188 5302 13216 7686
rect 13280 6934 13308 7754
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 6644 13308 6870
rect 13372 6746 13400 8044
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7274 13492 7890
rect 13556 7562 13584 10066
rect 13648 9654 13676 12566
rect 13924 12458 13952 12974
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13740 12430 13952 12458
rect 13740 10996 13768 12430
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 12209 13860 12242
rect 13818 12200 13874 12209
rect 13818 12135 13874 12144
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 11393 13860 11698
rect 13924 11694 13952 12310
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13818 11384 13874 11393
rect 13818 11319 13874 11328
rect 13832 11150 13860 11319
rect 13924 11286 13952 11630
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14002 11112 14058 11121
rect 14002 11047 14004 11056
rect 14056 11047 14058 11056
rect 14004 11018 14056 11024
rect 13740 10968 13952 10996
rect 13726 10840 13782 10849
rect 13726 10775 13782 10784
rect 13740 10742 13768 10775
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13924 10198 13952 10968
rect 14002 10976 14058 10985
rect 14002 10911 14058 10920
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 14016 10044 14044 10911
rect 13818 10024 13874 10033
rect 13728 9988 13780 9994
rect 13818 9959 13874 9968
rect 13924 10016 14044 10044
rect 13728 9930 13780 9936
rect 13740 9722 13768 9930
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13648 8362 13676 9114
rect 13726 9072 13782 9081
rect 13726 9007 13782 9016
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13634 8256 13690 8265
rect 13634 8191 13690 8200
rect 13648 7818 13676 8191
rect 13740 8090 13768 9007
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13832 7834 13860 9959
rect 13924 9178 13952 10016
rect 14002 9888 14058 9897
rect 14002 9823 14058 9832
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13924 7886 13952 8978
rect 14016 8634 14044 9823
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14016 8265 14044 8434
rect 14002 8256 14058 8265
rect 14002 8191 14058 8200
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13740 7806 13860 7834
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13556 7534 13676 7562
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13372 6718 13492 6746
rect 13280 6616 13400 6644
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 5386 13308 6190
rect 13372 5817 13400 6616
rect 13358 5808 13414 5817
rect 13358 5743 13414 5752
rect 13280 5358 13318 5386
rect 13176 5296 13228 5302
rect 13290 5284 13318 5358
rect 13176 5238 13228 5244
rect 13280 5256 13318 5284
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13188 4690 13216 5102
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13004 3534 13032 3674
rect 13096 3534 13124 3878
rect 13188 3738 13216 4490
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13004 3233 13032 3334
rect 12990 3224 13046 3233
rect 12900 3188 12952 3194
rect 12990 3159 13046 3168
rect 12900 3130 12952 3136
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 13280 1630 13308 5256
rect 13464 5114 13492 6718
rect 13372 5086 13492 5114
rect 13372 4146 13400 5086
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13464 4865 13492 4966
rect 13450 4856 13506 4865
rect 13450 4791 13506 4800
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13360 3052 13412 3058
rect 13464 3040 13492 4626
rect 13556 3194 13584 7414
rect 13648 3942 13676 7534
rect 13740 6644 13768 7806
rect 13820 7744 13872 7750
rect 13818 7712 13820 7721
rect 13872 7712 13874 7721
rect 13818 7647 13874 7656
rect 13924 7410 13952 7822
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13924 7206 13952 7346
rect 13912 7200 13964 7206
rect 13818 7168 13874 7177
rect 13912 7142 13964 7148
rect 13818 7103 13874 7112
rect 13832 7018 13860 7103
rect 13832 6990 13952 7018
rect 13740 6616 13860 6644
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13740 4865 13768 6326
rect 13726 4856 13782 4865
rect 13726 4791 13782 4800
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13740 4457 13768 4490
rect 13726 4448 13782 4457
rect 13726 4383 13782 4392
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13740 3942 13768 4082
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13648 3058 13676 3130
rect 13412 3012 13492 3040
rect 13636 3052 13688 3058
rect 13360 2994 13412 3000
rect 13636 2994 13688 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13648 2854 13676 2994
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13740 2582 13768 2994
rect 13832 2854 13860 6616
rect 13924 5030 13952 6990
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 14016 6361 14044 6870
rect 14002 6352 14058 6361
rect 14002 6287 14058 6296
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14016 5642 14044 5782
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 14002 5536 14058 5545
rect 14002 5471 14058 5480
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14016 4622 14044 5471
rect 14108 5370 14136 12854
rect 14200 10577 14228 16612
rect 14476 16538 14504 20703
rect 14568 19446 14596 22510
rect 14660 22438 14688 22646
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14292 16510 14504 16538
rect 14292 14550 14320 16510
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14384 15881 14412 15982
rect 14370 15872 14426 15881
rect 14370 15807 14426 15816
rect 14280 14544 14332 14550
rect 14280 14486 14332 14492
rect 14476 14346 14504 16390
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14292 13190 14320 14282
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14384 12434 14412 14214
rect 14462 13424 14518 13433
rect 14462 13359 14518 13368
rect 14476 13258 14504 13359
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14292 12406 14412 12434
rect 14462 12472 14518 12481
rect 14462 12407 14518 12416
rect 14292 12170 14320 12406
rect 14476 12288 14504 12407
rect 14568 12374 14596 19382
rect 14660 17610 14688 20334
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14660 16590 14688 17546
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14660 15337 14688 15370
rect 14646 15328 14702 15337
rect 14646 15263 14702 15272
rect 14646 14512 14702 14521
rect 14646 14447 14702 14456
rect 14660 13870 14688 14447
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14384 12260 14504 12288
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 11354 14320 12106
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14186 10568 14242 10577
rect 14186 10503 14242 10512
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10305 14228 10406
rect 14186 10296 14242 10305
rect 14186 10231 14242 10240
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 14200 8401 14228 10134
rect 14292 8888 14320 11290
rect 14384 9994 14412 12260
rect 14554 12200 14610 12209
rect 14554 12135 14610 12144
rect 14568 11830 14596 12135
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14476 10985 14504 11630
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 11393 14596 11562
rect 14554 11384 14610 11393
rect 14554 11319 14610 11328
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14462 10976 14518 10985
rect 14462 10911 14518 10920
rect 14464 10736 14516 10742
rect 14462 10704 14464 10713
rect 14516 10704 14518 10713
rect 14462 10639 14518 10648
rect 14476 10441 14504 10639
rect 14462 10432 14518 10441
rect 14462 10367 14518 10376
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 9081 14412 9318
rect 14370 9072 14426 9081
rect 14370 9007 14426 9016
rect 14372 8900 14424 8906
rect 14292 8860 14372 8888
rect 14372 8842 14424 8848
rect 14476 8498 14504 9998
rect 14568 9500 14596 11018
rect 14660 9654 14688 12718
rect 14752 12481 14780 24772
rect 14844 23254 14872 25230
rect 14832 23248 14884 23254
rect 14832 23190 14884 23196
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 21486 14872 22374
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 20602 14872 20742
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 14936 19786 14964 26726
rect 15028 24750 15056 29679
rect 15304 29170 15332 29718
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 15200 28688 15252 28694
rect 15200 28630 15252 28636
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 15028 24410 15056 24686
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15120 24138 15148 27610
rect 15212 27402 15240 28630
rect 15304 27402 15332 29106
rect 15396 28490 15424 29786
rect 15384 28484 15436 28490
rect 15384 28426 15436 28432
rect 15200 27396 15252 27402
rect 15200 27338 15252 27344
rect 15292 27396 15344 27402
rect 15292 27338 15344 27344
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15212 26353 15240 26726
rect 15198 26344 15254 26353
rect 15198 26279 15254 26288
rect 15198 26208 15254 26217
rect 15198 26143 15254 26152
rect 15212 25906 15240 26143
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15200 25424 15252 25430
rect 15200 25366 15252 25372
rect 15212 24682 15240 25366
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15304 24562 15332 27338
rect 15396 25974 15424 28426
rect 15384 25968 15436 25974
rect 15384 25910 15436 25916
rect 15384 25696 15436 25702
rect 15488 25673 15516 29990
rect 15568 29844 15620 29850
rect 15568 29786 15620 29792
rect 15580 29238 15608 29786
rect 16500 29646 16528 30126
rect 16488 29640 16540 29646
rect 16488 29582 16540 29588
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15658 29200 15714 29209
rect 15658 29135 15660 29144
rect 15712 29135 15714 29144
rect 15660 29106 15712 29112
rect 15764 29073 15792 29446
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 15750 29064 15806 29073
rect 15750 28999 15806 29008
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15580 26858 15608 28018
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15568 26852 15620 26858
rect 15568 26794 15620 26800
rect 15672 26625 15700 26930
rect 15658 26616 15714 26625
rect 15658 26551 15714 26560
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15384 25638 15436 25644
rect 15474 25664 15530 25673
rect 15212 24534 15332 24562
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15016 24064 15068 24070
rect 15106 24032 15162 24041
rect 15068 24012 15106 24018
rect 15016 24006 15106 24012
rect 15028 23990 15106 24006
rect 15106 23967 15162 23976
rect 15016 23044 15068 23050
rect 15016 22986 15068 22992
rect 15028 22030 15056 22986
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15028 20913 15056 21490
rect 15014 20904 15070 20913
rect 15014 20839 15070 20848
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14830 19544 14886 19553
rect 14830 19479 14886 19488
rect 14924 19508 14976 19514
rect 14844 19446 14872 19479
rect 14924 19450 14976 19456
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 14936 18970 14964 19450
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14844 17542 14872 17818
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14738 12472 14794 12481
rect 14738 12407 14794 12416
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14568 9472 14688 9500
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14186 8392 14242 8401
rect 14186 8327 14242 8336
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 7342 14228 8230
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14186 7168 14242 7177
rect 14186 7103 14242 7112
rect 14200 6662 14228 7103
rect 14292 6798 14320 8434
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14188 6384 14240 6390
rect 14188 6326 14240 6332
rect 14200 5778 14228 6326
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14292 5710 14320 6598
rect 14384 5846 14412 8026
rect 14462 7712 14518 7721
rect 14462 7647 14518 7656
rect 14476 6798 14504 7647
rect 14568 6798 14596 9114
rect 14660 8090 14688 9472
rect 14752 9178 14780 12310
rect 14844 11642 14872 15914
rect 14936 12434 14964 18158
rect 15028 16454 15056 20839
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15028 15337 15056 16118
rect 15014 15328 15070 15337
rect 15014 15263 15070 15272
rect 15120 15094 15148 23967
rect 15212 23866 15240 24534
rect 15200 23860 15252 23866
rect 15200 23802 15252 23808
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15304 23497 15332 23802
rect 15290 23488 15346 23497
rect 15290 23423 15346 23432
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15212 22166 15240 22918
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15198 21720 15254 21729
rect 15304 21706 15332 22578
rect 15396 21962 15424 25638
rect 15474 25599 15530 25608
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15488 23254 15516 25434
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15580 22817 15608 25774
rect 15672 24750 15700 26386
rect 15764 24886 15792 28358
rect 15844 26512 15896 26518
rect 15844 26454 15896 26460
rect 15856 26042 15884 26454
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15948 25786 15976 29106
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 16120 27940 16172 27946
rect 16120 27882 16172 27888
rect 16132 27402 16160 27882
rect 16224 27606 16252 28494
rect 16396 28076 16448 28082
rect 16396 28018 16448 28024
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16212 27600 16264 27606
rect 16212 27542 16264 27548
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 16212 27396 16264 27402
rect 16212 27338 16264 27344
rect 16028 26988 16080 26994
rect 16028 26930 16080 26936
rect 16040 26330 16068 26930
rect 16132 26450 16160 27338
rect 16120 26444 16172 26450
rect 16120 26386 16172 26392
rect 16040 26302 16160 26330
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 15856 25758 15976 25786
rect 15856 25401 15884 25758
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15842 25392 15898 25401
rect 15842 25327 15898 25336
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15660 24744 15712 24750
rect 15660 24686 15712 24692
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15566 22808 15622 22817
rect 15566 22743 15622 22752
rect 15672 22522 15700 24346
rect 15764 22642 15792 24618
rect 15856 24313 15884 25230
rect 15948 25226 15976 25638
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 16040 25106 16068 25910
rect 15948 25078 16068 25106
rect 15842 24304 15898 24313
rect 15842 24239 15898 24248
rect 15948 22710 15976 25078
rect 16026 23760 16082 23769
rect 16026 23695 16082 23704
rect 16040 23594 16068 23695
rect 16028 23588 16080 23594
rect 16028 23530 16080 23536
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15672 22494 15792 22522
rect 15658 22400 15714 22409
rect 15658 22335 15714 22344
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15672 21894 15700 22335
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15254 21678 15332 21706
rect 15198 21655 15254 21664
rect 15304 20992 15332 21678
rect 15382 21720 15438 21729
rect 15382 21655 15384 21664
rect 15436 21655 15438 21664
rect 15384 21626 15436 21632
rect 15212 20964 15332 20992
rect 15212 20380 15240 20964
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15304 20602 15332 20810
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15292 20392 15344 20398
rect 15212 20352 15292 20380
rect 15396 20369 15424 20810
rect 15292 20334 15344 20340
rect 15382 20360 15438 20369
rect 15382 20295 15438 20304
rect 15198 19544 15254 19553
rect 15198 19479 15254 19488
rect 15212 17066 15240 19479
rect 15396 18698 15424 20295
rect 15488 18970 15516 20878
rect 15566 20768 15622 20777
rect 15566 20703 15622 20712
rect 15580 19786 15608 20703
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15580 19446 15608 19722
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15396 17954 15424 18634
rect 15488 18601 15516 18702
rect 15568 18692 15620 18698
rect 15568 18634 15620 18640
rect 15474 18592 15530 18601
rect 15474 18527 15530 18536
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15304 17926 15424 17954
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15212 16833 15240 17002
rect 15198 16824 15254 16833
rect 15198 16759 15254 16768
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15120 14618 15148 14826
rect 15212 14618 15240 16458
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15304 14498 15332 17926
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15396 16726 15424 17206
rect 15488 17066 15516 18158
rect 15580 17610 15608 18634
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15474 16824 15530 16833
rect 15474 16759 15530 16768
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15396 15881 15424 16118
rect 15382 15872 15438 15881
rect 15382 15807 15438 15816
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15212 14470 15332 14498
rect 15396 14482 15424 14894
rect 15384 14476 15436 14482
rect 15016 14000 15068 14006
rect 15120 13988 15148 14418
rect 15068 13960 15148 13988
rect 15016 13942 15068 13948
rect 15120 13240 15148 13960
rect 15212 13870 15240 14470
rect 15384 14418 15436 14424
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15120 13212 15332 13240
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 14936 12406 15148 12434
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14844 11614 14964 11642
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11082 14872 11494
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14830 10568 14886 10577
rect 14830 10503 14886 10512
rect 14844 10266 14872 10503
rect 14936 10266 14964 11614
rect 15028 11218 15056 12106
rect 15120 11558 15148 12406
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15120 10305 15148 11290
rect 15212 10742 15240 13087
rect 15304 12306 15332 13212
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15396 11830 15424 14418
rect 15488 13161 15516 16759
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 14958 15608 16594
rect 15672 15042 15700 18566
rect 15764 17746 15792 22494
rect 16028 22092 16080 22098
rect 16028 22034 16080 22040
rect 15936 21956 15988 21962
rect 15936 21898 15988 21904
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15856 21622 15884 21830
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 20262 15884 21422
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19786 15884 20198
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15764 15162 15792 17682
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15672 15014 15792 15042
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 13388 15620 13394
rect 15672 13376 15700 14214
rect 15620 13348 15700 13376
rect 15568 13330 15620 13336
rect 15474 13152 15530 13161
rect 15474 13087 15530 13096
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15384 11824 15436 11830
rect 15304 11784 15384 11812
rect 15304 11354 15332 11784
rect 15384 11766 15436 11772
rect 15488 11665 15516 12310
rect 15474 11656 15530 11665
rect 15384 11620 15436 11626
rect 15474 11591 15530 11600
rect 15384 11562 15436 11568
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15396 11234 15424 11562
rect 15304 11206 15424 11234
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15106 10296 15162 10305
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14924 10260 14976 10266
rect 15106 10231 15162 10240
rect 14924 10202 14976 10208
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14844 9602 14872 10066
rect 14936 9674 14964 10202
rect 15304 10062 15332 11206
rect 15580 11132 15608 13330
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15396 11104 15608 11132
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 14936 9646 15056 9674
rect 14844 9574 14964 9602
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14740 9036 14792 9042
rect 14740 8978 14792 8984
rect 14752 8906 14780 8978
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14844 8294 14872 8570
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14476 5386 14504 6734
rect 14660 6361 14688 7754
rect 14844 7750 14872 8230
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14646 6352 14702 6361
rect 14646 6287 14702 6296
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5846 14688 6054
rect 14648 5840 14700 5846
rect 14648 5782 14700 5788
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14372 5364 14424 5370
rect 14476 5358 14596 5386
rect 14372 5306 14424 5312
rect 14280 5228 14332 5234
rect 14108 5188 14280 5216
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13924 4146 13952 4558
rect 14108 4146 14136 5188
rect 14280 5170 14332 5176
rect 14186 4856 14242 4865
rect 14186 4791 14242 4800
rect 14200 4690 14228 4791
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 14384 4282 14412 5306
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14476 4758 14504 5238
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14476 4146 14504 4694
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14108 4049 14136 4082
rect 14292 4049 14320 4082
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 14462 4040 14518 4049
rect 14568 4010 14596 5358
rect 14646 4856 14702 4865
rect 14646 4791 14648 4800
rect 14700 4791 14702 4800
rect 14648 4762 14700 4768
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 4282 14688 4626
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14462 3975 14464 3984
rect 14108 3777 14136 3975
rect 14516 3975 14518 3984
rect 14556 4004 14608 4010
rect 14464 3946 14516 3952
rect 14556 3946 14608 3952
rect 14094 3768 14150 3777
rect 14094 3703 14150 3712
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13268 1624 13320 1630
rect 13268 1566 13320 1572
rect 13648 1562 13676 2246
rect 13636 1556 13688 1562
rect 13636 1498 13688 1504
rect 12900 1216 12952 1222
rect 12900 1158 12952 1164
rect 12912 800 12940 1158
rect 14200 800 14228 3606
rect 14476 3534 14504 3946
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14568 3058 14596 3946
rect 14752 3942 14780 7686
rect 14844 7177 14872 7686
rect 14830 7168 14886 7177
rect 14830 7103 14886 7112
rect 14936 6610 14964 9574
rect 15028 9432 15056 9646
rect 15108 9444 15160 9450
rect 15028 9404 15108 9432
rect 15108 9386 15160 9392
rect 15212 8616 15240 9930
rect 15304 9450 15332 9998
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 14844 6582 14964 6610
rect 15028 8588 15240 8616
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14844 3534 14872 6582
rect 15028 6474 15056 8588
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15198 8392 15254 8401
rect 15198 8327 15254 8336
rect 15212 7546 15240 8327
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15198 7168 15254 7177
rect 15198 7103 15254 7112
rect 15212 6905 15240 7103
rect 15198 6896 15254 6905
rect 15198 6831 15254 6840
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14936 6446 15056 6474
rect 14936 4604 14964 6446
rect 15120 6254 15148 6734
rect 15198 6624 15254 6633
rect 15198 6559 15254 6568
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15108 5636 15160 5642
rect 15108 5578 15160 5584
rect 15028 4758 15056 5578
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15016 4616 15068 4622
rect 14936 4576 15016 4604
rect 15016 4558 15068 4564
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14752 3058 14780 3130
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14476 2310 14504 2586
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14384 1426 14412 2246
rect 14372 1420 14424 1426
rect 14372 1362 14424 1368
rect 14844 800 14872 2382
rect 15028 2145 15056 4558
rect 15120 4457 15148 5578
rect 15212 5545 15240 6559
rect 15304 6236 15332 8502
rect 15396 6390 15424 11104
rect 15672 10792 15700 13194
rect 15764 12918 15792 15014
rect 15856 14657 15884 18906
rect 15842 14648 15898 14657
rect 15842 14583 15898 14592
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15764 11286 15792 12854
rect 15856 12850 15884 13874
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 11626 15884 12786
rect 15948 12594 15976 21898
rect 16040 21486 16068 22034
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16132 20942 16160 26302
rect 16224 25498 16252 27338
rect 16212 25492 16264 25498
rect 16212 25434 16264 25440
rect 16316 25226 16344 27814
rect 16408 27674 16436 28018
rect 16396 27668 16448 27674
rect 16396 27610 16448 27616
rect 16500 27554 16528 29582
rect 16776 28558 16804 37402
rect 17420 36854 17448 39200
rect 18064 37262 18092 39200
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 17408 36848 17460 36854
rect 17408 36790 17460 36796
rect 17972 31822 18000 37062
rect 19352 36922 19380 39200
rect 19996 37126 20024 39200
rect 20168 37392 20220 37398
rect 20168 37334 20220 37340
rect 20076 37256 20128 37262
rect 20076 37198 20128 37204
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 18696 36576 18748 36582
rect 18696 36518 18748 36524
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 18708 31346 18736 36518
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 17592 31272 17644 31278
rect 17592 31214 17644 31220
rect 17498 29472 17554 29481
rect 17498 29407 17554 29416
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16868 28762 16896 29106
rect 16856 28756 16908 28762
rect 16856 28698 16908 28704
rect 16580 28552 16632 28558
rect 16580 28494 16632 28500
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16592 27606 16620 28494
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16408 27526 16528 27554
rect 16580 27600 16632 27606
rect 16580 27542 16632 27548
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 16120 20936 16172 20942
rect 16026 20904 16082 20913
rect 16120 20878 16172 20884
rect 16026 20839 16082 20848
rect 16040 19961 16068 20839
rect 16118 20768 16174 20777
rect 16118 20703 16174 20712
rect 16132 20398 16160 20703
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16026 19952 16082 19961
rect 16026 19887 16082 19896
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16040 13190 16068 19450
rect 16118 18592 16174 18601
rect 16118 18527 16174 18536
rect 16132 17785 16160 18527
rect 16118 17776 16174 17785
rect 16118 17711 16174 17720
rect 16118 14648 16174 14657
rect 16118 14583 16174 14592
rect 16132 13297 16160 14583
rect 16224 14521 16252 22986
rect 16316 22438 16344 24686
rect 16408 23905 16436 27526
rect 16578 27024 16634 27033
rect 16578 26959 16634 26968
rect 16592 26450 16620 26959
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16500 25498 16528 25978
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16592 25158 16620 26250
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16394 23896 16450 23905
rect 16394 23831 16450 23840
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16316 21554 16344 22374
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16408 21400 16436 23462
rect 16488 22976 16540 22982
rect 16592 22964 16620 25094
rect 16684 23050 16712 27950
rect 16762 26480 16818 26489
rect 16762 26415 16818 26424
rect 16776 25412 16804 26415
rect 16868 25537 16896 28698
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17420 28393 17448 28494
rect 17406 28384 17462 28393
rect 17406 28319 17462 28328
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 16948 27872 17000 27878
rect 16948 27814 17000 27820
rect 16960 27713 16988 27814
rect 16946 27704 17002 27713
rect 16946 27639 17002 27648
rect 17052 27470 17080 28018
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16854 25528 16910 25537
rect 16854 25463 16910 25472
rect 16776 25384 16896 25412
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16776 23594 16804 24074
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 16672 23044 16724 23050
rect 16672 22986 16724 22992
rect 16540 22936 16620 22964
rect 16488 22918 16540 22924
rect 16500 22166 16528 22918
rect 16670 22808 16726 22817
rect 16670 22743 16726 22752
rect 16578 22672 16634 22681
rect 16684 22642 16712 22743
rect 16776 22642 16804 23530
rect 16868 23254 16896 25384
rect 16856 23248 16908 23254
rect 16856 23190 16908 23196
rect 16578 22607 16634 22616
rect 16672 22636 16724 22642
rect 16592 22438 16620 22607
rect 16672 22578 16724 22584
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16500 21729 16528 21898
rect 16486 21720 16542 21729
rect 16486 21655 16542 21664
rect 16408 21372 16528 21400
rect 16304 21140 16356 21146
rect 16356 21100 16436 21128
rect 16304 21082 16356 21088
rect 16408 20942 16436 21100
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 19553 16344 20334
rect 16394 19816 16450 19825
rect 16394 19751 16450 19760
rect 16302 19544 16358 19553
rect 16302 19479 16358 19488
rect 16408 18329 16436 19751
rect 16500 19514 16528 21372
rect 16592 21146 16620 21898
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16684 21026 16712 22578
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16776 21962 16804 22170
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16868 21842 16896 22442
rect 16960 21894 16988 26726
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 17052 24410 17080 24822
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 17040 24064 17092 24070
rect 17040 24006 17092 24012
rect 17052 22386 17080 24006
rect 17144 22506 17172 28154
rect 17512 28082 17540 29407
rect 17604 28558 17632 31214
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18512 30320 18564 30326
rect 18512 30262 18564 30268
rect 18328 29708 18380 29714
rect 18328 29650 18380 29656
rect 18340 29034 18368 29650
rect 18328 29028 18380 29034
rect 18380 28976 18460 28994
rect 18328 28970 18460 28976
rect 18340 28966 18460 28970
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 17500 28076 17552 28082
rect 17500 28018 17552 28024
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17420 27402 17448 27950
rect 17512 27878 17540 28018
rect 17500 27872 17552 27878
rect 17500 27814 17552 27820
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17408 27396 17460 27402
rect 17408 27338 17460 27344
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17328 26382 17356 26930
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17236 24342 17264 26182
rect 17420 24800 17448 27338
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17604 26897 17632 26930
rect 17590 26888 17646 26897
rect 17590 26823 17646 26832
rect 17592 26784 17644 26790
rect 17592 26726 17644 26732
rect 17500 25220 17552 25226
rect 17500 25162 17552 25168
rect 17512 24886 17540 25162
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17328 24772 17448 24800
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17224 23656 17276 23662
rect 17222 23624 17224 23633
rect 17276 23624 17278 23633
rect 17222 23559 17278 23568
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 17132 22500 17184 22506
rect 17132 22442 17184 22448
rect 17052 22358 17172 22386
rect 16592 20998 16712 21026
rect 16776 21814 16896 21842
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16592 20602 16620 20998
rect 16670 20768 16726 20777
rect 16670 20703 16726 20712
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16684 19417 16712 20703
rect 16776 20058 16804 21814
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16670 19408 16726 19417
rect 16670 19343 16726 19352
rect 16684 18408 16712 19343
rect 16868 18970 16896 20810
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16960 19922 16988 19994
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16946 19544 17002 19553
rect 16946 19479 17002 19488
rect 16960 19446 16988 19479
rect 16948 19440 17000 19446
rect 16948 19382 17000 19388
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16868 18698 16896 18906
rect 16856 18692 16908 18698
rect 16856 18634 16908 18640
rect 16684 18380 16804 18408
rect 16394 18320 16450 18329
rect 16394 18255 16450 18264
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 15638 16344 16390
rect 16408 16250 16436 18022
rect 16500 16538 16528 18158
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16592 17785 16620 17818
rect 16578 17776 16634 17785
rect 16578 17711 16634 17720
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16592 17338 16620 17478
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16592 16658 16620 17070
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16500 16510 16620 16538
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16500 15745 16528 16390
rect 16486 15736 16542 15745
rect 16486 15671 16542 15680
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16408 15366 16436 15574
rect 16592 15552 16620 16510
rect 16500 15524 16620 15552
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 14793 16344 14894
rect 16302 14784 16358 14793
rect 16302 14719 16358 14728
rect 16408 14634 16436 15098
rect 16500 14793 16528 15524
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16486 14784 16542 14793
rect 16486 14719 16542 14728
rect 16316 14606 16436 14634
rect 16210 14512 16266 14521
rect 16210 14447 16266 14456
rect 16316 14006 16344 14606
rect 16486 14512 16542 14521
rect 16396 14476 16448 14482
rect 16592 14482 16620 15370
rect 16684 15026 16712 18226
rect 16776 16182 16804 18380
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 16960 18154 16988 18294
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16762 15600 16818 15609
rect 16762 15535 16818 15544
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16670 14784 16726 14793
rect 16670 14719 16726 14728
rect 16486 14447 16542 14456
rect 16580 14476 16632 14482
rect 16396 14418 16448 14424
rect 16408 14249 16436 14418
rect 16394 14240 16450 14249
rect 16394 14175 16450 14184
rect 16304 14000 16356 14006
rect 16500 13977 16528 14447
rect 16580 14418 16632 14424
rect 16304 13942 16356 13948
rect 16486 13968 16542 13977
rect 16486 13903 16542 13912
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16118 13288 16174 13297
rect 16118 13223 16174 13232
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16224 12730 16252 13738
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16408 13394 16436 13631
rect 16684 13512 16712 14719
rect 16776 14482 16804 15535
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16868 14278 16896 17818
rect 17052 17746 17080 21830
rect 17144 21554 17172 22358
rect 17236 22166 17264 23122
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17144 21457 17172 21490
rect 17130 21448 17186 21457
rect 17130 21383 17186 21392
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17144 20874 17172 21014
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17144 19310 17172 20538
rect 17236 20398 17264 21966
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17328 19922 17356 24772
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 23662 17540 24550
rect 17604 24138 17632 26726
rect 17696 26353 17724 27270
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17682 26344 17738 26353
rect 17682 26279 17738 26288
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17696 25809 17724 25842
rect 17682 25800 17738 25809
rect 17682 25735 17738 25744
rect 17788 24410 17816 26386
rect 17880 26194 17908 27406
rect 18052 27396 18104 27402
rect 18052 27338 18104 27344
rect 17880 26166 18000 26194
rect 17972 25294 18000 26166
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17788 24138 17816 24346
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17880 23905 17908 24754
rect 17972 24070 18000 25230
rect 18064 24750 18092 27338
rect 18236 26784 18288 26790
rect 18236 26726 18288 26732
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 17866 23896 17922 23905
rect 17866 23831 17922 23840
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17880 23594 17908 23734
rect 17958 23624 18014 23633
rect 17868 23588 17920 23594
rect 17958 23559 17960 23568
rect 17868 23530 17920 23536
rect 18012 23559 18014 23568
rect 17960 23530 18012 23536
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17420 21894 17448 23122
rect 17684 22772 17736 22778
rect 17736 22732 17908 22760
rect 17684 22714 17736 22720
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17512 20398 17540 22170
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 17314 19408 17370 19417
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17236 18902 17264 19382
rect 17314 19343 17370 19352
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17130 17776 17186 17785
rect 17040 17740 17092 17746
rect 17130 17711 17186 17720
rect 17040 17682 17092 17688
rect 17144 17513 17172 17711
rect 17328 17542 17356 19343
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17420 18698 17448 18838
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17512 17592 17540 20334
rect 17604 19786 17632 22442
rect 17880 21876 17908 22732
rect 17958 22536 18014 22545
rect 17958 22471 18014 22480
rect 17972 22137 18000 22471
rect 17958 22128 18014 22137
rect 17958 22063 18014 22072
rect 17972 22030 18000 22063
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17880 21848 18000 21876
rect 18064 21865 18092 24006
rect 17866 21720 17922 21729
rect 17866 21655 17922 21664
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17604 19417 17632 19722
rect 17590 19408 17646 19417
rect 17590 19343 17646 19352
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17420 17564 17540 17592
rect 17316 17536 17368 17542
rect 17130 17504 17186 17513
rect 17316 17478 17368 17484
rect 17130 17439 17186 17448
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 16946 16824 17002 16833
rect 17052 16794 17080 17206
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 16946 16759 16948 16768
rect 17000 16759 17002 16768
rect 17040 16788 17092 16794
rect 16948 16730 17000 16736
rect 17040 16730 17092 16736
rect 17144 16266 17172 17002
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 16960 16238 17172 16266
rect 16960 16046 16988 16238
rect 17038 16144 17094 16153
rect 17038 16079 17094 16088
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16684 13484 16804 13512
rect 16776 13394 16804 13484
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16684 13258 16712 13330
rect 16868 13297 16896 14214
rect 16960 14006 16988 15982
rect 17052 15745 17080 16079
rect 17224 15972 17276 15978
rect 17224 15914 17276 15920
rect 17038 15736 17094 15745
rect 17038 15671 17094 15680
rect 17236 15502 17264 15914
rect 17328 15609 17356 16458
rect 17420 16182 17448 17564
rect 17604 17524 17632 19246
rect 17512 17496 17632 17524
rect 17512 16776 17540 17496
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17604 17066 17632 17274
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17512 16748 17632 16776
rect 17604 16658 17632 16748
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17314 15600 17370 15609
rect 17314 15535 17370 15544
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17052 15008 17080 15098
rect 17132 15020 17184 15026
rect 17052 14980 17132 15008
rect 17132 14962 17184 14968
rect 17236 14498 17264 15438
rect 17314 15056 17370 15065
rect 17314 14991 17370 15000
rect 17328 14958 17356 14991
rect 17316 14952 17368 14958
rect 17420 14940 17448 15982
rect 17512 15570 17540 16594
rect 17590 16144 17646 16153
rect 17590 16079 17646 16088
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17604 15502 17632 16079
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17696 15162 17724 19722
rect 17788 18057 17816 21490
rect 17880 20874 17908 21655
rect 17972 20942 18000 21848
rect 18050 21856 18106 21865
rect 18050 21791 18106 21800
rect 18156 21622 18184 26386
rect 18248 26081 18276 26726
rect 18234 26072 18290 26081
rect 18234 26007 18290 26016
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18340 25906 18368 25978
rect 18328 25900 18380 25906
rect 18328 25842 18380 25848
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18156 21049 18184 21286
rect 18142 21040 18198 21049
rect 18142 20975 18198 20984
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17880 20777 17908 20810
rect 17866 20768 17922 20777
rect 17866 20703 17922 20712
rect 17958 20632 18014 20641
rect 17958 20567 18014 20576
rect 17972 20466 18000 20567
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17880 20318 18092 20346
rect 17880 20262 17908 20318
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17880 18970 17908 19246
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17972 18834 18000 20198
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17958 18728 18014 18737
rect 18064 18714 18092 20318
rect 18156 19530 18184 20975
rect 18248 19689 18276 25094
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18340 23050 18368 24550
rect 18328 23044 18380 23050
rect 18328 22986 18380 22992
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 18234 19680 18290 19689
rect 18234 19615 18290 19624
rect 18156 19502 18276 19530
rect 18142 19408 18198 19417
rect 18142 19343 18144 19352
rect 18196 19343 18198 19352
rect 18144 19314 18196 19320
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18156 18902 18184 19178
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18248 18834 18276 19502
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18064 18686 18184 18714
rect 17958 18663 18014 18672
rect 17972 18630 18000 18663
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 18352 18012 18358
rect 17958 18320 17960 18329
rect 18012 18320 18014 18329
rect 17958 18255 18014 18264
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17972 17882 18000 18158
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17788 17066 17816 17546
rect 17880 17134 17908 17546
rect 17960 17536 18012 17542
rect 17958 17504 17960 17513
rect 18012 17504 18014 17513
rect 17958 17439 18014 17448
rect 17868 17128 17920 17134
rect 17960 17128 18012 17134
rect 17868 17070 17920 17076
rect 17958 17096 17960 17105
rect 18012 17096 18014 17105
rect 17776 17060 17828 17066
rect 17958 17031 18014 17040
rect 17776 17002 17828 17008
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17788 16130 17816 16594
rect 17788 16102 18000 16130
rect 17788 15473 17816 16102
rect 17972 16046 18000 16102
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17774 15464 17830 15473
rect 17774 15399 17830 15408
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17500 15088 17552 15094
rect 17552 15048 17632 15076
rect 17500 15030 17552 15036
rect 17420 14912 17533 14940
rect 17316 14894 17368 14900
rect 17505 14770 17533 14912
rect 17604 14770 17632 15048
rect 17880 14958 17908 15982
rect 18064 14958 18092 18566
rect 18156 15745 18184 18686
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18142 15736 18198 15745
rect 18142 15671 18198 15680
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17505 14742 17540 14770
rect 17604 14742 18000 14770
rect 17512 14634 17540 14742
rect 17512 14606 17632 14634
rect 17604 14600 17632 14606
rect 17604 14572 17816 14600
rect 17144 14470 17264 14498
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17500 14544 17552 14550
rect 17788 14532 17816 14572
rect 17972 14550 18000 14742
rect 17960 14544 18012 14550
rect 17788 14504 17908 14532
rect 17500 14486 17552 14492
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16946 13560 17002 13569
rect 16946 13495 17002 13504
rect 16960 13326 16988 13495
rect 16948 13320 17000 13326
rect 16854 13288 16910 13297
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16672 13252 16724 13258
rect 16948 13262 17000 13268
rect 16854 13223 16910 13232
rect 16672 13194 16724 13200
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 12850 16344 13126
rect 16408 12986 16436 13194
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 15948 12566 16068 12594
rect 15934 12472 15990 12481
rect 15934 12407 15990 12416
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15948 11506 15976 12407
rect 15856 11478 15976 11506
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15856 11218 15884 11478
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15580 10764 15700 10792
rect 15476 10736 15528 10742
rect 15580 10724 15608 10764
rect 15856 10742 15884 11018
rect 15528 10696 15608 10724
rect 15844 10736 15896 10742
rect 15476 10678 15528 10684
rect 15844 10678 15896 10684
rect 15750 10432 15806 10441
rect 15750 10367 15806 10376
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15672 9761 15700 10134
rect 15658 9752 15714 9761
rect 15658 9687 15714 9696
rect 15660 9512 15712 9518
rect 15580 9472 15660 9500
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 8566 15516 8910
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15580 8294 15608 9472
rect 15660 9454 15712 9460
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15488 8266 15608 8294
rect 15488 7410 15516 8266
rect 15566 7576 15622 7585
rect 15566 7511 15622 7520
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15474 7032 15530 7041
rect 15474 6967 15530 6976
rect 15488 6633 15516 6967
rect 15474 6624 15530 6633
rect 15474 6559 15530 6568
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15304 6208 15516 6236
rect 15382 5672 15438 5681
rect 15382 5607 15438 5616
rect 15198 5536 15254 5545
rect 15198 5471 15254 5480
rect 15198 5400 15254 5409
rect 15198 5335 15200 5344
rect 15252 5335 15254 5344
rect 15200 5306 15252 5312
rect 15198 4856 15254 4865
rect 15198 4791 15254 4800
rect 15212 4486 15240 4791
rect 15290 4720 15346 4729
rect 15290 4655 15292 4664
rect 15344 4655 15346 4664
rect 15292 4626 15344 4632
rect 15200 4480 15252 4486
rect 15106 4448 15162 4457
rect 15200 4422 15252 4428
rect 15106 4383 15162 4392
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15120 3942 15148 4014
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15212 3534 15240 3946
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15396 3194 15424 5607
rect 15488 3534 15516 6208
rect 15580 4146 15608 7511
rect 15672 7041 15700 9114
rect 15658 7032 15714 7041
rect 15658 6967 15714 6976
rect 15672 6798 15700 6967
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15658 6352 15714 6361
rect 15658 6287 15714 6296
rect 15672 5545 15700 6287
rect 15658 5536 15714 5545
rect 15658 5471 15714 5480
rect 15764 5370 15792 10367
rect 16040 10112 16068 12566
rect 15856 10084 16068 10112
rect 15856 9897 15884 10084
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15842 9888 15898 9897
rect 15842 9823 15898 9832
rect 15856 8430 15884 9823
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15856 7002 15884 7346
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 5642 15884 6734
rect 15844 5636 15896 5642
rect 15844 5578 15896 5584
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15764 4486 15792 5170
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15752 4480 15804 4486
rect 15856 4457 15884 4558
rect 15752 4422 15804 4428
rect 15842 4448 15898 4457
rect 15842 4383 15898 4392
rect 15856 4146 15884 4383
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15856 4049 15884 4082
rect 15842 4040 15898 4049
rect 15568 4004 15620 4010
rect 15842 3975 15898 3984
rect 15568 3946 15620 3952
rect 15580 3913 15608 3946
rect 15566 3904 15622 3913
rect 15566 3839 15622 3848
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15014 2136 15070 2145
rect 15014 2071 15070 2080
rect 15212 1494 15240 2382
rect 15488 2281 15516 3334
rect 15672 2774 15700 3402
rect 15856 3058 15884 3975
rect 15948 3942 15976 9930
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16040 9761 16068 9862
rect 16026 9752 16082 9761
rect 16026 9687 16082 9696
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16040 9518 16068 9590
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16132 8922 16160 12718
rect 16224 12702 16344 12730
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 11665 16252 12582
rect 16210 11656 16266 11665
rect 16210 11591 16266 11600
rect 16316 11540 16344 12702
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16224 11512 16344 11540
rect 16224 10588 16252 11512
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16316 10742 16344 11290
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16224 10560 16344 10588
rect 16210 10160 16266 10169
rect 16316 10130 16344 10560
rect 16210 10095 16266 10104
rect 16304 10124 16356 10130
rect 16224 9926 16252 10095
rect 16304 10066 16356 10072
rect 16302 10024 16358 10033
rect 16302 9959 16304 9968
rect 16356 9959 16358 9968
rect 16304 9930 16356 9936
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16316 9654 16344 9930
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16408 9500 16436 12174
rect 16500 11694 16528 12650
rect 16592 12306 16620 13126
rect 16670 13016 16726 13025
rect 17052 13002 17080 14282
rect 16670 12951 16726 12960
rect 16868 12974 17080 13002
rect 16684 12753 16712 12951
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16670 12744 16726 12753
rect 16670 12679 16726 12688
rect 16776 12481 16804 12854
rect 16762 12472 16818 12481
rect 16762 12407 16818 12416
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16868 12050 16896 12974
rect 17040 12912 17092 12918
rect 17144 12900 17172 14470
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 13569 17264 14350
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17222 13560 17278 13569
rect 17222 13495 17278 13504
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17092 12872 17172 12900
rect 17040 12854 17092 12860
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 12646 17080 12718
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 16868 12022 16988 12050
rect 16856 11892 16908 11898
rect 16684 11852 16856 11880
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 10130 16528 11494
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16592 11082 16620 11290
rect 16580 11076 16632 11082
rect 16684 11064 16712 11852
rect 16856 11834 16908 11840
rect 16764 11280 16816 11286
rect 16816 11240 16896 11268
rect 16764 11222 16816 11228
rect 16684 11036 16804 11064
rect 16580 11018 16632 11024
rect 16670 10976 16726 10985
rect 16670 10911 16726 10920
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16500 9586 16528 10066
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16316 9472 16436 9500
rect 16210 9344 16266 9353
rect 16210 9279 16266 9288
rect 16040 8894 16160 8922
rect 16040 7721 16068 8894
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16026 7712 16082 7721
rect 16026 7647 16082 7656
rect 16132 7410 16160 8774
rect 16224 8673 16252 9279
rect 16210 8664 16266 8673
rect 16210 8599 16266 8608
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16224 7206 16252 8599
rect 16316 7834 16344 9472
rect 16486 9072 16542 9081
rect 16486 9007 16542 9016
rect 16500 8906 16528 9007
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16486 8664 16542 8673
rect 16486 8599 16488 8608
rect 16540 8599 16542 8608
rect 16488 8570 16540 8576
rect 16592 8514 16620 10474
rect 16684 9994 16712 10911
rect 16776 10169 16804 11036
rect 16762 10160 16818 10169
rect 16762 10095 16818 10104
rect 16762 10024 16818 10033
rect 16672 9988 16724 9994
rect 16762 9959 16818 9968
rect 16672 9930 16724 9936
rect 16776 9761 16804 9959
rect 16762 9752 16818 9761
rect 16762 9687 16818 9696
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16776 9500 16804 9590
rect 16868 9586 16896 11240
rect 16960 10742 16988 12022
rect 17052 11218 17080 12242
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16776 9472 16813 9500
rect 16785 9432 16813 9472
rect 16776 9404 16813 9432
rect 16776 9042 16804 9404
rect 16960 9081 16988 10678
rect 16946 9072 17002 9081
rect 16764 9036 16816 9042
rect 16946 9007 17002 9016
rect 16764 8978 16816 8984
rect 17052 8922 17080 11154
rect 16500 8486 16620 8514
rect 16684 8894 17080 8922
rect 16396 8424 16448 8430
rect 16394 8392 16396 8401
rect 16448 8392 16450 8401
rect 16394 8327 16450 8336
rect 16316 7806 16436 7834
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 5710 16160 6598
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16118 5536 16174 5545
rect 16118 5471 16174 5480
rect 16132 5234 16160 5471
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 16224 3641 16252 6734
rect 16316 5234 16344 7686
rect 16408 5681 16436 7806
rect 16500 7546 16528 8486
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16592 6633 16620 8366
rect 16684 7954 16712 8894
rect 17144 8809 17172 12872
rect 17236 12288 17264 13330
rect 17328 12866 17356 13806
rect 17420 13308 17448 14486
rect 17512 14278 17540 14486
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17604 13870 17632 14418
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17500 13320 17552 13326
rect 17420 13280 17500 13308
rect 17500 13262 17552 13268
rect 17328 12838 17540 12866
rect 17512 12782 17540 12838
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17590 12744 17646 12753
rect 17236 12260 17448 12288
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 11218 17356 12106
rect 17316 11212 17368 11218
rect 17420 11200 17448 12260
rect 17512 11898 17540 12718
rect 17590 12679 17646 12688
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17604 11694 17632 12679
rect 17696 12434 17724 14282
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17788 13734 17816 14214
rect 17880 14006 17908 14504
rect 17960 14486 18012 14492
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18064 14396 18092 14486
rect 17972 14368 18092 14396
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 12918 17908 13670
rect 17972 13258 18000 14368
rect 18156 14328 18184 15098
rect 18248 14328 18276 18022
rect 18340 17241 18368 22646
rect 18432 19961 18460 28966
rect 18524 27470 18552 30262
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18708 29646 18736 29786
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18616 28150 18644 28902
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18708 27146 18736 29582
rect 18616 27118 18736 27146
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18524 21622 18552 26998
rect 18616 24596 18644 27118
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18708 26382 18736 26930
rect 18800 26450 18828 30534
rect 18880 29708 18932 29714
rect 18880 29650 18932 29656
rect 18892 29102 18920 29650
rect 19352 29594 19380 31758
rect 19444 31482 19472 36722
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19996 30666 20024 31078
rect 19984 30660 20036 30666
rect 19984 30602 20036 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19352 29572 20024 29594
rect 19352 29566 19524 29572
rect 19576 29566 20024 29572
rect 19524 29514 19576 29520
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19524 29300 19576 29306
rect 19524 29242 19576 29248
rect 18972 29232 19024 29238
rect 18972 29174 19024 29180
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18708 25294 18736 26318
rect 18892 25786 18920 29038
rect 18984 28762 19012 29174
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 18972 28756 19024 28762
rect 18972 28698 19024 28704
rect 19064 28688 19116 28694
rect 19064 28630 19116 28636
rect 19076 28558 19104 28630
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 19154 28520 19210 28529
rect 19352 28506 19380 29038
rect 19154 28455 19156 28464
rect 19208 28455 19210 28464
rect 19260 28478 19380 28506
rect 19156 28426 19208 28432
rect 19064 28416 19116 28422
rect 19064 28358 19116 28364
rect 18970 28248 19026 28257
rect 18970 28183 19026 28192
rect 18984 28150 19012 28183
rect 18972 28144 19024 28150
rect 18972 28086 19024 28092
rect 19076 27062 19104 28358
rect 19260 28218 19288 28478
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 19156 27464 19208 27470
rect 19156 27406 19208 27412
rect 19064 27056 19116 27062
rect 19064 26998 19116 27004
rect 18892 25758 19012 25786
rect 18880 25696 18932 25702
rect 18880 25638 18932 25644
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18800 24954 18828 25094
rect 18788 24948 18840 24954
rect 18788 24890 18840 24896
rect 18696 24608 18748 24614
rect 18616 24576 18696 24596
rect 18748 24576 18750 24585
rect 18616 24568 18694 24576
rect 18694 24511 18750 24520
rect 18892 24342 18920 25638
rect 18984 25362 19012 25758
rect 18972 25356 19024 25362
rect 18972 25298 19024 25304
rect 18984 24750 19012 25298
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18696 24200 18748 24206
rect 18748 24160 18828 24188
rect 18696 24142 18748 24148
rect 18696 22704 18748 22710
rect 18616 22664 18696 22692
rect 18616 22234 18644 22664
rect 18696 22646 18748 22652
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18708 22409 18736 22510
rect 18694 22400 18750 22409
rect 18694 22335 18750 22344
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18800 22137 18828 24160
rect 19168 23361 19196 27406
rect 19352 27062 19380 28358
rect 19444 28014 19472 29174
rect 19536 28937 19564 29242
rect 19996 29186 20024 29566
rect 19812 29158 20024 29186
rect 19522 28928 19578 28937
rect 19522 28863 19578 28872
rect 19812 28529 19840 29158
rect 19984 29028 20036 29034
rect 19984 28970 20036 28976
rect 19798 28520 19854 28529
rect 19798 28455 19854 28464
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19996 27614 20024 28970
rect 20088 28762 20116 37198
rect 20180 35894 20208 37334
rect 20640 37330 20668 39200
rect 20628 37324 20680 37330
rect 20628 37266 20680 37272
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 20916 36854 20944 37198
rect 21928 37108 21956 39200
rect 22572 37330 22600 39200
rect 22744 37460 22796 37466
rect 22744 37402 22796 37408
rect 22560 37324 22612 37330
rect 22560 37266 22612 37272
rect 21928 37080 22140 37108
rect 22112 36922 22140 37080
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 20904 36848 20956 36854
rect 20904 36790 20956 36796
rect 20180 35866 20300 35894
rect 20168 30320 20220 30326
rect 20168 30262 20220 30268
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 20076 28144 20128 28150
rect 20074 28112 20076 28121
rect 20128 28112 20130 28121
rect 20074 28047 20130 28056
rect 19996 27586 20116 27614
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19444 27062 19472 27406
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19432 27056 19484 27062
rect 19432 26998 19484 27004
rect 19430 26888 19486 26897
rect 19430 26823 19486 26832
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19260 24886 19288 26250
rect 19338 25800 19394 25809
rect 19338 25735 19340 25744
rect 19392 25735 19394 25744
rect 19340 25706 19392 25712
rect 19444 25702 19472 26823
rect 19996 26314 20024 27270
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19536 25226 19564 25706
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19812 25362 19840 25434
rect 19800 25356 19852 25362
rect 19800 25298 19852 25304
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19248 24880 19300 24886
rect 19248 24822 19300 24828
rect 19248 24336 19300 24342
rect 19248 24278 19300 24284
rect 19260 23798 19288 24278
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19154 23352 19210 23361
rect 19154 23287 19210 23296
rect 18880 23044 18932 23050
rect 18880 22986 18932 22992
rect 18892 22778 18920 22986
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18878 22264 18934 22273
rect 18878 22199 18934 22208
rect 18786 22128 18842 22137
rect 18786 22063 18842 22072
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 21690 18828 21830
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18524 21457 18552 21558
rect 18510 21448 18566 21457
rect 18510 21383 18566 21392
rect 18708 21078 18736 21626
rect 18788 21412 18840 21418
rect 18788 21354 18840 21360
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18524 20641 18552 20946
rect 18510 20632 18566 20641
rect 18510 20567 18566 20576
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18708 20398 18736 20538
rect 18800 20534 18828 21354
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18696 20392 18748 20398
rect 18616 20352 18696 20380
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18418 19952 18474 19961
rect 18418 19887 18474 19896
rect 18432 19854 18460 19887
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18524 19666 18552 20198
rect 18432 19638 18552 19666
rect 18432 18290 18460 19638
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18524 18358 18552 19450
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18510 18048 18566 18057
rect 18432 17814 18460 18022
rect 18510 17983 18566 17992
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18326 17232 18382 17241
rect 18326 17167 18382 17176
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 14657 18368 14826
rect 18326 14648 18382 14657
rect 18326 14583 18382 14592
rect 18432 14464 18460 17614
rect 18524 17338 18552 17983
rect 18616 17338 18644 20352
rect 18696 20334 18748 20340
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18800 20058 18828 20334
rect 18892 20058 18920 22199
rect 19168 21706 19196 23287
rect 18984 21678 19196 21706
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18984 19938 19012 21678
rect 19352 21486 19380 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19706 24440 19762 24449
rect 19996 24410 20024 24550
rect 19706 24375 19762 24384
rect 19984 24404 20036 24410
rect 19720 24342 19748 24375
rect 19984 24346 20036 24352
rect 19708 24336 19760 24342
rect 19708 24278 19760 24284
rect 19430 24032 19486 24041
rect 19430 23967 19486 23976
rect 19444 23798 19472 23967
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19800 23792 19852 23798
rect 19800 23734 19852 23740
rect 19892 23792 19944 23798
rect 19892 23734 19944 23740
rect 19812 23662 19840 23734
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 19444 22098 19472 23530
rect 19904 23186 19932 23734
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20088 22556 20116 27586
rect 20180 26994 20208 30262
rect 20272 28694 20300 35866
rect 20444 33380 20496 33386
rect 20444 33322 20496 33328
rect 20352 31204 20404 31210
rect 20352 31146 20404 31152
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 20364 28642 20392 31146
rect 20456 29238 20484 33322
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20640 30433 20668 31282
rect 20626 30424 20682 30433
rect 20626 30359 20682 30368
rect 20720 29776 20772 29782
rect 20720 29718 20772 29724
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20628 29232 20680 29238
rect 20628 29174 20680 29180
rect 20364 28614 20484 28642
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20272 28150 20300 28358
rect 20260 28144 20312 28150
rect 20260 28086 20312 28092
rect 20364 26994 20392 28494
rect 20456 27614 20484 28614
rect 20534 28112 20590 28121
rect 20534 28047 20590 28056
rect 20548 28014 20576 28047
rect 20536 28008 20588 28014
rect 20536 27950 20588 27956
rect 20456 27586 20576 27614
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20272 24954 20300 25910
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20168 24744 20220 24750
rect 20166 24712 20168 24721
rect 20220 24712 20222 24721
rect 20166 24647 20222 24656
rect 20272 23032 20300 24890
rect 20456 23338 20484 26726
rect 20548 24342 20576 27586
rect 20536 24336 20588 24342
rect 20536 24278 20588 24284
rect 20536 24132 20588 24138
rect 20536 24074 20588 24080
rect 20364 23310 20484 23338
rect 20364 23186 20392 23310
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 20272 23004 20484 23032
rect 20350 22808 20406 22817
rect 20350 22743 20406 22752
rect 20364 22642 20392 22743
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 19522 22536 19578 22545
rect 20088 22528 20300 22556
rect 19522 22471 19578 22480
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19536 21978 19564 22471
rect 20074 22264 20130 22273
rect 20074 22199 20076 22208
rect 20128 22199 20130 22208
rect 20076 22170 20128 22176
rect 19444 21950 19564 21978
rect 19444 21729 19472 21950
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19430 21720 19486 21729
rect 19574 21723 19882 21732
rect 19430 21655 19486 21664
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 19340 21480 19392 21486
rect 19062 21448 19118 21457
rect 19340 21422 19392 21428
rect 19062 21383 19118 21392
rect 19076 20262 19104 21383
rect 19522 21312 19578 21321
rect 19260 21270 19522 21298
rect 19156 20800 19208 20806
rect 19154 20768 19156 20777
rect 19208 20768 19210 20777
rect 19154 20703 19210 20712
rect 19260 20602 19288 21270
rect 19522 21247 19578 21256
rect 19352 21134 20024 21162
rect 19352 21078 19380 21134
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 19444 20924 19472 21014
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19352 20896 19472 20924
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19352 20482 19380 20896
rect 19812 20874 19840 20946
rect 19524 20868 19576 20874
rect 19444 20828 19524 20856
rect 19444 20777 19472 20828
rect 19524 20810 19576 20816
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19430 20768 19486 20777
rect 19430 20703 19486 20712
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19430 20632 19486 20641
rect 19574 20635 19882 20644
rect 19996 20641 20024 21134
rect 20180 20777 20208 21558
rect 20272 21486 20300 22528
rect 20456 22522 20484 23004
rect 20364 22494 20484 22522
rect 20260 21480 20312 21486
rect 20260 21422 20312 21428
rect 20166 20768 20222 20777
rect 20166 20703 20222 20712
rect 19982 20632 20038 20641
rect 19430 20567 19432 20576
rect 19484 20567 19486 20576
rect 19892 20596 19944 20602
rect 19432 20538 19484 20544
rect 20272 20584 20300 21422
rect 20364 20874 20392 22494
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 20364 20777 20392 20810
rect 20350 20768 20406 20777
rect 20350 20703 20406 20712
rect 19982 20567 20038 20576
rect 19892 20538 19944 20544
rect 20180 20556 20300 20584
rect 19168 20454 19380 20482
rect 19616 20460 19668 20466
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19168 20074 19196 20454
rect 19444 20420 19616 20448
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 18708 19910 19012 19938
rect 19076 20046 19196 20074
rect 18708 19281 18736 19910
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18800 19446 18828 19654
rect 18984 19514 19012 19722
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 19076 19360 19104 20046
rect 19260 19825 19288 20198
rect 19444 19990 19472 20420
rect 19616 20402 19668 20408
rect 19904 20210 19932 20538
rect 20076 20528 20128 20534
rect 20180 20516 20208 20556
rect 20456 20534 20484 22170
rect 20548 21298 20576 24074
rect 20640 22438 20668 29174
rect 20732 27606 20760 29718
rect 20916 29646 20944 36790
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 22376 36780 22428 36786
rect 22376 36722 22428 36728
rect 21284 36650 21312 36722
rect 21272 36644 21324 36650
rect 21272 36586 21324 36592
rect 21180 33312 21232 33318
rect 21180 33254 21232 33260
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21088 29096 21140 29102
rect 21088 29038 21140 29044
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20824 28558 20852 28902
rect 20812 28552 20864 28558
rect 20812 28494 20864 28500
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20732 24274 20760 26862
rect 20824 26518 20852 27474
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20824 25906 20852 26454
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20824 24886 20852 25842
rect 21100 25770 21128 29038
rect 21192 25906 21220 33254
rect 21284 30258 21312 36586
rect 22388 36378 22416 36722
rect 21916 36372 21968 36378
rect 21916 36314 21968 36320
rect 22376 36372 22428 36378
rect 22376 36314 22428 36320
rect 21548 36100 21600 36106
rect 21548 36042 21600 36048
rect 21560 31754 21588 36042
rect 21928 31754 21956 36314
rect 22100 33992 22152 33998
rect 22100 33934 22152 33940
rect 21560 31726 21680 31754
rect 21364 30796 21416 30802
rect 21364 30738 21416 30744
rect 21376 30326 21404 30738
rect 21364 30320 21416 30326
rect 21416 30280 21496 30308
rect 21364 30262 21416 30268
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 21468 27606 21496 30280
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 21456 27600 21508 27606
rect 21456 27542 21508 27548
rect 21560 27538 21588 28358
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21284 26432 21312 27066
rect 21376 27010 21404 27270
rect 21468 27130 21496 27338
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21376 26982 21496 27010
rect 21284 26404 21404 26432
rect 21376 26314 21404 26404
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21088 25764 21140 25770
rect 21088 25706 21140 25712
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 24886 21036 25638
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 21376 24682 21404 26250
rect 21364 24676 21416 24682
rect 21364 24618 21416 24624
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20732 22545 20760 24210
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20824 22710 20852 23258
rect 20916 23050 20944 23598
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20718 22536 20774 22545
rect 20718 22471 20774 22480
rect 20812 22500 20864 22506
rect 20812 22442 20864 22448
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20548 21270 20668 21298
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20128 20488 20208 20516
rect 20444 20528 20496 20534
rect 20076 20470 20128 20476
rect 20444 20470 20496 20476
rect 20352 20450 20404 20456
rect 20352 20392 20404 20398
rect 19984 20324 20036 20330
rect 20364 20312 20392 20392
rect 20036 20284 20392 20312
rect 19984 20266 20036 20272
rect 19904 20182 20300 20210
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19628 19922 19656 19994
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19246 19816 19302 19825
rect 19706 19816 19762 19825
rect 19352 19786 19706 19802
rect 19246 19751 19302 19760
rect 19340 19780 19706 19786
rect 19392 19774 19706 19780
rect 19706 19751 19762 19760
rect 19340 19722 19392 19728
rect 19904 19700 19932 19926
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19444 19672 19932 19700
rect 19444 19553 19472 19672
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19430 19544 19486 19553
rect 19574 19547 19882 19556
rect 19430 19479 19486 19488
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19616 19440 19668 19446
rect 19536 19400 19616 19428
rect 19076 19332 19288 19360
rect 18880 19304 18932 19310
rect 18694 19272 18750 19281
rect 18880 19246 18932 19252
rect 18972 19304 19024 19310
rect 19154 19272 19210 19281
rect 18972 19246 19024 19252
rect 18694 19207 18750 19216
rect 18786 19000 18842 19009
rect 18786 18935 18842 18944
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18512 17128 18564 17134
rect 18564 17088 18644 17116
rect 18512 17070 18564 17076
rect 18510 16688 18566 16697
rect 18510 16623 18566 16632
rect 18064 14300 18184 14328
rect 18237 14300 18276 14328
rect 18340 14436 18460 14464
rect 18064 13938 18092 14300
rect 18237 14260 18265 14300
rect 18156 14232 18265 14260
rect 18156 13938 18184 14232
rect 18340 14090 18368 14436
rect 18524 14396 18552 16623
rect 18616 16590 18644 17088
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18248 14062 18368 14090
rect 18432 14368 18552 14396
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18248 13818 18276 14062
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18156 13790 18276 13818
rect 18340 13818 18368 13942
rect 18432 13938 18460 14368
rect 18510 14240 18566 14249
rect 18510 14175 18566 14184
rect 18524 14006 18552 14175
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18510 13832 18566 13841
rect 18340 13802 18460 13818
rect 18340 13796 18472 13802
rect 18340 13790 18420 13796
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18064 13138 18092 13738
rect 17972 13110 18092 13138
rect 18156 13138 18184 13790
rect 18510 13767 18566 13776
rect 18420 13738 18472 13744
rect 18524 13734 18552 13767
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18340 13376 18368 13670
rect 18616 13444 18644 16118
rect 18708 14890 18736 18226
rect 18800 17954 18828 18935
rect 18892 18426 18920 19246
rect 18984 18970 19012 19246
rect 19076 19230 19154 19258
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18972 18760 19024 18766
rect 18970 18728 18972 18737
rect 19024 18728 19026 18737
rect 18970 18663 19026 18672
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18984 18222 19012 18566
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18880 18080 18932 18086
rect 18932 18040 19012 18068
rect 18880 18022 18932 18028
rect 18800 17926 18920 17954
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18800 16182 18828 17682
rect 18892 17134 18920 17926
rect 18984 17814 19012 18040
rect 19076 17954 19104 19230
rect 19154 19207 19210 19216
rect 19154 19136 19210 19145
rect 19154 19071 19210 19080
rect 19168 18601 19196 19071
rect 19260 18698 19288 19332
rect 19338 19000 19394 19009
rect 19338 18935 19394 18944
rect 19352 18834 19380 18935
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19340 18624 19392 18630
rect 19154 18592 19210 18601
rect 19154 18527 19210 18536
rect 19260 18572 19340 18578
rect 19536 18612 19564 19400
rect 19616 19382 19668 19388
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19628 18834 19656 19246
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19720 18698 19748 19178
rect 19996 18970 20024 19450
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19977 18692 20029 18698
rect 19977 18634 20029 18640
rect 19260 18566 19392 18572
rect 19444 18584 19564 18612
rect 19260 18550 19380 18566
rect 19260 18442 19288 18550
rect 19168 18414 19288 18442
rect 19444 18426 19472 18584
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18420 19484 18426
rect 19168 18154 19196 18414
rect 19432 18362 19484 18368
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 19616 18352 19668 18358
rect 19616 18294 19668 18300
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19076 17926 19196 17954
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 19064 17264 19116 17270
rect 19168 17241 19196 17926
rect 19260 17626 19288 18294
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19260 17598 19380 17626
rect 19536 17610 19564 18022
rect 19628 17882 19656 18294
rect 19996 18272 20024 18634
rect 19904 18244 20024 18272
rect 19904 17882 19932 18244
rect 20088 17898 20116 19858
rect 20166 19816 20222 19825
rect 20166 19751 20222 19760
rect 20180 19514 20208 19751
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20272 19378 20300 20182
rect 20352 19984 20404 19990
rect 20352 19926 20404 19932
rect 20442 19952 20498 19961
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20166 19000 20222 19009
rect 20166 18935 20222 18944
rect 20364 18952 20392 19926
rect 20442 19887 20498 19896
rect 20456 19514 20484 19887
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20548 19394 20576 21082
rect 20640 20505 20668 21270
rect 20732 21010 20760 21422
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20626 20496 20682 20505
rect 20626 20431 20682 20440
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20456 19366 20576 19394
rect 20640 19378 20668 19450
rect 20628 19372 20680 19378
rect 20456 19310 20484 19366
rect 20732 19360 20760 20198
rect 20824 19990 20852 22442
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 21008 19938 21036 24278
rect 21100 23662 21128 24550
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 21192 21554 21220 24346
rect 21284 23526 21312 24346
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21468 23254 21496 26982
rect 21560 24750 21588 27474
rect 21652 26353 21680 31726
rect 21744 31726 21956 31754
rect 21638 26344 21694 26353
rect 21638 26279 21694 26288
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 24818 21680 25774
rect 21640 24812 21692 24818
rect 21640 24754 21692 24760
rect 21548 24744 21600 24750
rect 21548 24686 21600 24692
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21548 24336 21600 24342
rect 21548 24278 21600 24284
rect 21560 23254 21588 24278
rect 21652 23798 21680 24550
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 21456 23248 21508 23254
rect 21456 23190 21508 23196
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 21560 23050 21588 23190
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21270 22536 21326 22545
rect 21270 22471 21326 22480
rect 21284 22438 21312 22471
rect 21272 22432 21324 22438
rect 21272 22374 21324 22380
rect 21456 22432 21508 22438
rect 21456 22374 21508 22380
rect 21364 22092 21416 22098
rect 21364 22034 21416 22040
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21284 21690 21312 21898
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21088 21344 21140 21350
rect 21376 21321 21404 22034
rect 21088 21286 21140 21292
rect 21362 21312 21418 21321
rect 21100 20058 21128 21286
rect 21362 21247 21418 21256
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21008 19910 21128 19938
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20732 19332 20852 19360
rect 20628 19314 20680 19320
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20626 19272 20682 19281
rect 20444 19168 20496 19174
rect 20442 19136 20444 19145
rect 20496 19136 20498 19145
rect 20442 19071 20498 19080
rect 20180 18748 20208 18935
rect 20364 18924 20484 18952
rect 20350 18864 20406 18873
rect 20350 18799 20406 18808
rect 20180 18737 20300 18748
rect 20180 18728 20314 18737
rect 20180 18720 20258 18728
rect 20258 18663 20314 18672
rect 20364 18612 20392 18799
rect 20272 18584 20392 18612
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 19996 17870 20116 17898
rect 19996 17796 20024 17870
rect 19989 17768 20024 17796
rect 19989 17728 20017 17768
rect 19989 17700 20024 17728
rect 19996 17626 20024 17700
rect 19064 17206 19116 17212
rect 19154 17232 19210 17241
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18878 16688 18934 16697
rect 18878 16623 18934 16632
rect 18892 16454 18920 16623
rect 19076 16522 19104 17206
rect 19154 17167 19210 17176
rect 19352 17184 19380 17598
rect 19524 17604 19576 17610
rect 19996 17598 20116 17626
rect 19524 17546 19576 17552
rect 19984 17536 20036 17542
rect 19982 17504 19984 17513
rect 20036 17504 20038 17513
rect 19574 17436 19882 17445
rect 19982 17439 20038 17448
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19982 17368 20038 17377
rect 19982 17303 20038 17312
rect 19614 17232 19670 17241
rect 19352 17156 19472 17184
rect 19996 17218 20024 17303
rect 20088 17270 20116 17598
rect 20180 17513 20208 18022
rect 20166 17504 20222 17513
rect 20166 17439 20222 17448
rect 19614 17167 19670 17176
rect 19720 17190 20024 17218
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20168 17196 20220 17202
rect 19338 17096 19394 17105
rect 19338 17031 19394 17040
rect 19352 16833 19380 17031
rect 19338 16824 19394 16833
rect 19338 16759 19394 16768
rect 19444 16574 19472 17156
rect 19522 16824 19578 16833
rect 19522 16759 19578 16768
rect 19168 16546 19472 16574
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18878 16280 18934 16289
rect 18878 16215 18934 16224
rect 19062 16280 19118 16289
rect 19062 16215 19118 16224
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18892 16046 18920 16215
rect 18880 16040 18932 16046
rect 19076 16017 19104 16215
rect 18880 15982 18932 15988
rect 19062 16008 19118 16017
rect 19062 15943 19118 15952
rect 19062 15736 19118 15745
rect 19062 15671 19118 15680
rect 18972 15564 19024 15570
rect 19076 15552 19104 15671
rect 19024 15524 19104 15552
rect 18972 15506 19024 15512
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18800 14618 18828 14894
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18708 14498 18736 14554
rect 18708 14470 18744 14498
rect 18716 14328 18744 14470
rect 18708 14300 18744 14328
rect 18708 13841 18736 14300
rect 18694 13832 18750 13841
rect 18694 13767 18750 13776
rect 18616 13416 18828 13444
rect 18340 13348 18736 13376
rect 18708 13258 18736 13348
rect 18236 13252 18288 13258
rect 18604 13252 18656 13258
rect 18288 13212 18460 13240
rect 18236 13194 18288 13200
rect 18156 13110 18276 13138
rect 17868 12912 17920 12918
rect 17972 12900 18000 13110
rect 18248 12918 18276 13110
rect 18236 12912 18288 12918
rect 17972 12872 18092 12900
rect 17868 12854 17920 12860
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17958 12744 18014 12753
rect 17696 12406 17816 12434
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17696 12170 17724 12310
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17420 11172 17632 11200
rect 17316 11154 17368 11160
rect 17406 11112 17462 11121
rect 17406 11047 17462 11056
rect 17500 11076 17552 11082
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17236 10266 17264 10542
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17328 10062 17356 10542
rect 17420 10198 17448 11047
rect 17500 11018 17552 11024
rect 17512 10248 17540 11018
rect 17604 10418 17632 11172
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17696 10810 17724 10911
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17788 10520 17816 12406
rect 17880 12374 17908 12718
rect 17958 12679 18014 12688
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17972 12186 18000 12679
rect 18064 12306 18092 12872
rect 18236 12854 18288 12860
rect 18326 12744 18382 12753
rect 18156 12702 18326 12730
rect 18156 12646 18184 12702
rect 18432 12714 18460 13212
rect 18604 13194 18656 13200
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18616 12730 18644 13194
rect 18326 12679 18382 12688
rect 18420 12708 18472 12714
rect 18616 12702 18736 12730
rect 18420 12650 18472 12656
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17880 10810 17908 12174
rect 17972 12158 18092 12186
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17972 10674 18000 11766
rect 18064 11082 18092 12158
rect 18340 11898 18368 12582
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18328 11756 18380 11762
rect 18380 11716 18460 11744
rect 18328 11698 18380 11704
rect 18236 11688 18288 11694
rect 18234 11656 18236 11665
rect 18432 11665 18460 11716
rect 18288 11656 18290 11665
rect 18234 11591 18290 11600
rect 18418 11656 18474 11665
rect 18418 11591 18474 11600
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18052 11076 18104 11082
rect 18052 11018 18104 11024
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17788 10492 17908 10520
rect 17604 10390 17816 10418
rect 17788 10266 17816 10390
rect 17684 10260 17736 10266
rect 17512 10220 17632 10248
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17236 9761 17264 9862
rect 17222 9752 17278 9761
rect 17222 9687 17278 9696
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 16946 8800 17002 8809
rect 17130 8800 17186 8809
rect 17002 8758 17080 8786
rect 16946 8735 17002 8744
rect 16762 8664 16818 8673
rect 16762 8599 16818 8608
rect 17052 8616 17080 8758
rect 17130 8735 17186 8744
rect 17132 8628 17184 8634
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16394 5672 16450 5681
rect 16394 5607 16450 5616
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16408 4622 16436 5607
rect 16500 5545 16528 6258
rect 16486 5536 16542 5545
rect 16486 5471 16542 5480
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16500 4826 16528 5306
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16408 3641 16436 4111
rect 16592 3738 16620 6326
rect 16684 4826 16712 7754
rect 16776 6633 16804 8599
rect 17052 8588 17132 8616
rect 17132 8570 17184 8576
rect 16854 8392 16910 8401
rect 16854 8327 16910 8336
rect 16868 7954 16896 8327
rect 17236 8106 17264 9522
rect 17420 9110 17448 9862
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17406 8800 17462 8809
rect 17406 8735 17462 8744
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17328 8430 17356 8502
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17314 8120 17370 8129
rect 17236 8078 17314 8106
rect 17314 8055 17370 8064
rect 17420 8022 17448 8735
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 16960 7546 16988 7958
rect 17512 7886 17540 9998
rect 17604 9704 17632 10220
rect 17684 10202 17736 10208
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17696 10112 17724 10202
rect 17776 10124 17828 10130
rect 17696 10084 17776 10112
rect 17776 10066 17828 10072
rect 17604 9676 17816 9704
rect 17682 9616 17738 9625
rect 17682 9551 17738 9560
rect 17696 9194 17724 9551
rect 17788 9330 17816 9676
rect 17880 9674 17908 10492
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17972 9926 18000 10202
rect 18064 10169 18092 11018
rect 18050 10160 18106 10169
rect 18050 10095 18106 10104
rect 18156 9976 18184 11494
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18248 10985 18276 11018
rect 18234 10976 18290 10985
rect 18234 10911 18290 10920
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18248 10266 18276 10610
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18340 10044 18368 10610
rect 18432 10606 18460 11494
rect 18524 11014 18552 12106
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18524 10606 18552 10746
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18340 10016 18460 10044
rect 18156 9948 18368 9976
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 18052 9920 18104 9926
rect 18104 9868 18184 9874
rect 18052 9862 18184 9868
rect 18064 9846 18184 9862
rect 17880 9646 18092 9674
rect 17788 9302 18000 9330
rect 17696 9166 17908 9194
rect 17592 9036 17644 9042
rect 17644 8996 17724 9024
rect 17592 8978 17644 8984
rect 17696 8906 17724 8996
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17038 7576 17094 7585
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16948 7540 17000 7546
rect 17604 7562 17632 8298
rect 17094 7534 17632 7562
rect 17038 7511 17094 7520
rect 16948 7482 17000 7488
rect 16762 6624 16818 6633
rect 16762 6559 16818 6568
rect 16868 6361 16896 7482
rect 17040 7336 17092 7342
rect 17092 7296 17172 7324
rect 17040 7278 17092 7284
rect 17144 7154 17172 7296
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17144 7126 17264 7154
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17052 6746 17080 6938
rect 17144 6866 17172 6938
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17052 6718 17172 6746
rect 17144 6390 17172 6718
rect 17132 6384 17184 6390
rect 16854 6352 16910 6361
rect 17132 6326 17184 6332
rect 16854 6287 16910 6296
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16868 5574 16896 5646
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16762 5264 16818 5273
rect 16762 5199 16818 5208
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16776 4758 16804 5199
rect 16764 4752 16816 4758
rect 16670 4720 16726 4729
rect 16764 4694 16816 4700
rect 16670 4655 16672 4664
rect 16724 4655 16726 4664
rect 16672 4626 16724 4632
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16210 3632 16266 3641
rect 16210 3567 16266 3576
rect 16394 3632 16450 3641
rect 16394 3567 16450 3576
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 3398 16620 3470
rect 16580 3392 16632 3398
rect 16580 3334 16632 3340
rect 16592 3233 16620 3334
rect 16302 3224 16358 3233
rect 16302 3159 16358 3168
rect 16578 3224 16634 3233
rect 16578 3159 16634 3168
rect 16316 3058 16344 3159
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 15580 2746 15700 2774
rect 15474 2272 15530 2281
rect 15474 2207 15530 2216
rect 15580 1562 15608 2746
rect 15568 1556 15620 1562
rect 15568 1498 15620 1504
rect 15200 1488 15252 1494
rect 15200 1430 15252 1436
rect 16132 800 16160 2994
rect 16684 2825 16712 4082
rect 16960 3602 16988 6190
rect 17038 5944 17094 5953
rect 17038 5879 17040 5888
rect 17092 5879 17094 5888
rect 17040 5850 17092 5856
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 17052 4434 17080 4694
rect 17052 4406 17172 4434
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17052 4185 17080 4218
rect 17038 4176 17094 4185
rect 17038 4111 17094 4120
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16868 3466 16896 3538
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16764 2848 16816 2854
rect 16670 2816 16726 2825
rect 16764 2790 16816 2796
rect 16670 2751 16726 2760
rect 16776 800 16804 2790
rect 16868 2378 16896 2858
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 17144 1698 17172 4406
rect 17236 4282 17264 7126
rect 17328 6440 17356 7239
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17512 6633 17540 6802
rect 17498 6624 17554 6633
rect 17498 6559 17554 6568
rect 17328 6412 17448 6440
rect 17420 5522 17448 6412
rect 17498 6352 17554 6361
rect 17604 6322 17632 7534
rect 17498 6287 17554 6296
rect 17592 6316 17644 6322
rect 17512 6118 17540 6287
rect 17592 6258 17644 6264
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17498 5808 17554 5817
rect 17498 5743 17554 5752
rect 17328 5494 17448 5522
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17328 4010 17356 5494
rect 17512 5409 17540 5743
rect 17498 5400 17554 5409
rect 17408 5364 17460 5370
rect 17498 5335 17554 5344
rect 17408 5306 17460 5312
rect 17420 4758 17448 5306
rect 17500 5160 17552 5166
rect 17500 5102 17552 5108
rect 17512 5001 17540 5102
rect 17498 4992 17554 5001
rect 17498 4927 17554 4936
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17604 4486 17632 6258
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17512 4146 17540 4422
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17696 4010 17724 8842
rect 17880 8430 17908 9166
rect 17868 8424 17920 8430
rect 17972 8401 18000 9302
rect 17868 8366 17920 8372
rect 17958 8392 18014 8401
rect 17958 8327 18014 8336
rect 17774 8120 17830 8129
rect 17774 8055 17776 8064
rect 17828 8055 17830 8064
rect 17776 8026 17828 8032
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17776 7744 17828 7750
rect 17972 7732 18000 7890
rect 18064 7800 18092 9646
rect 18156 7868 18184 9846
rect 18340 9654 18368 9948
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18432 9602 18460 10016
rect 18524 9994 18552 10066
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18248 9518 18276 9590
rect 18432 9574 18552 9602
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 9110 18368 9386
rect 18328 9104 18380 9110
rect 18234 9072 18290 9081
rect 18328 9046 18380 9052
rect 18234 9007 18290 9016
rect 18248 8566 18276 9007
rect 18432 8786 18460 9454
rect 18340 8758 18460 8786
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18156 7840 18276 7868
rect 18064 7772 18184 7800
rect 17972 7704 18092 7732
rect 17776 7686 17828 7692
rect 17788 6322 17816 7686
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17880 7206 17908 7414
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17868 7200 17920 7206
rect 17972 7177 18000 7278
rect 17868 7142 17920 7148
rect 17958 7168 18014 7177
rect 17958 7103 18014 7112
rect 17868 6996 17920 7002
rect 17920 6956 18000 6984
rect 17868 6938 17920 6944
rect 17866 6760 17922 6769
rect 17866 6695 17922 6704
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17880 5914 17908 6695
rect 17972 6644 18000 6956
rect 18064 6866 18092 7704
rect 18156 7478 18184 7772
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 18248 7342 18276 7840
rect 18340 7800 18368 8758
rect 18524 8650 18552 9574
rect 18616 9518 18644 12582
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 8809 18644 9454
rect 18708 9178 18736 12702
rect 18800 12646 18828 13416
rect 18892 13410 18920 15302
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 18984 14822 19012 15030
rect 19076 15026 19104 15524
rect 19168 15366 19196 16546
rect 19536 16522 19564 16759
rect 19628 16538 19656 17167
rect 19720 16658 19748 17190
rect 20168 17138 20220 17144
rect 20180 16776 20208 17138
rect 20272 16946 20300 18584
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20364 17241 20392 18294
rect 20456 18154 20484 18924
rect 20548 18834 20576 19246
rect 20626 19207 20682 19216
rect 20536 18828 20588 18834
rect 20536 18770 20588 18776
rect 20640 18408 20668 19207
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18630 20760 19110
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20824 18426 20852 19332
rect 20916 18873 20944 19790
rect 20902 18864 20958 18873
rect 20902 18799 20958 18808
rect 21100 18714 21128 19910
rect 21192 19854 21220 20334
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21284 19786 21312 20198
rect 21376 20097 21404 21247
rect 21468 21146 21496 22374
rect 21638 22128 21694 22137
rect 21638 22063 21694 22072
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21362 20088 21418 20097
rect 21362 20023 21418 20032
rect 21468 19972 21496 20742
rect 21376 19944 21496 19972
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 20916 18686 21128 18714
rect 20548 18380 20668 18408
rect 20812 18420 20864 18426
rect 20444 18148 20496 18154
rect 20444 18090 20496 18096
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20456 17513 20484 17750
rect 20442 17504 20498 17513
rect 20442 17439 20498 17448
rect 20350 17232 20406 17241
rect 20350 17167 20406 17176
rect 20272 16918 20484 16946
rect 20088 16748 20208 16776
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19812 16538 19840 16594
rect 19524 16516 19576 16522
rect 19444 16476 19524 16504
rect 19246 16280 19302 16289
rect 19302 16238 19380 16266
rect 19246 16215 19302 16224
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19154 15192 19210 15201
rect 19154 15127 19156 15136
rect 19208 15127 19210 15136
rect 19156 15098 19208 15104
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 19168 14532 19196 14962
rect 19260 14958 19288 16118
rect 19352 16096 19380 16238
rect 19444 16232 19472 16476
rect 19628 16510 19840 16538
rect 19984 16516 20036 16522
rect 19524 16458 19576 16464
rect 19984 16458 20036 16464
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19444 16204 19564 16232
rect 19432 16108 19484 16114
rect 19352 16068 19432 16096
rect 19432 16050 19484 16056
rect 19536 15416 19564 16204
rect 19996 16182 20024 16458
rect 19800 16176 19852 16182
rect 19984 16176 20036 16182
rect 19852 16136 19932 16164
rect 19800 16118 19852 16124
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19352 15388 19564 15416
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19076 14504 19196 14532
rect 19076 14006 19104 14504
rect 19352 14464 19380 15388
rect 19628 15348 19656 16050
rect 19904 15366 19932 16136
rect 19984 16118 20036 16124
rect 19984 15904 20036 15910
rect 20088 15892 20116 16748
rect 20166 16688 20222 16697
rect 20456 16674 20484 16918
rect 20166 16623 20222 16632
rect 20272 16646 20484 16674
rect 20548 16658 20576 18380
rect 20812 18362 20864 18368
rect 20628 18284 20680 18290
rect 20680 18244 20852 18272
rect 20628 18226 20680 18232
rect 20824 18086 20852 18244
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20812 17740 20864 17746
rect 20916 17728 20944 18686
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20864 17700 20944 17728
rect 20812 17682 20864 17688
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20718 17232 20774 17241
rect 20718 17167 20774 17176
rect 20626 16688 20682 16697
rect 20536 16652 20588 16658
rect 20036 15864 20116 15892
rect 19984 15846 20036 15852
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 19444 15320 19656 15348
rect 19892 15360 19944 15366
rect 19444 15201 19472 15320
rect 19892 15302 19944 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19430 15192 19486 15201
rect 19574 15195 19882 15204
rect 19982 15192 20038 15201
rect 19430 15127 19486 15136
rect 19720 15136 19982 15144
rect 19720 15127 20038 15136
rect 20088 15144 20116 15370
rect 20180 15337 20208 16623
rect 20272 15502 20300 16646
rect 20732 16658 20760 17167
rect 20626 16623 20682 16632
rect 20720 16652 20772 16658
rect 20536 16594 20588 16600
rect 20352 16516 20404 16522
rect 20352 16458 20404 16464
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20166 15328 20222 15337
rect 20166 15263 20222 15272
rect 19720 15116 20024 15127
rect 20088 15116 20208 15144
rect 19432 15088 19484 15094
rect 19616 15088 19668 15094
rect 19484 15048 19616 15076
rect 19432 15030 19484 15036
rect 19616 15030 19668 15036
rect 19720 14890 19748 15116
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19904 14550 19932 14894
rect 19892 14544 19944 14550
rect 19892 14486 19944 14492
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19168 14436 19380 14464
rect 19168 14006 19196 14436
rect 19996 14362 20024 14486
rect 19444 14334 20024 14362
rect 19340 14272 19392 14278
rect 19338 14240 19340 14249
rect 19392 14240 19394 14249
rect 19338 14175 19394 14184
rect 19444 14113 19472 14334
rect 20088 14260 20116 14962
rect 20180 14770 20208 15116
rect 20364 14958 20392 16458
rect 20442 16416 20498 16425
rect 20442 16351 20498 16360
rect 20456 16114 20484 16351
rect 20534 16144 20590 16153
rect 20444 16108 20496 16114
rect 20534 16079 20590 16088
rect 20640 16096 20668 16623
rect 20720 16594 20772 16600
rect 20720 16108 20772 16114
rect 20444 16050 20496 16056
rect 20548 15586 20576 16079
rect 20640 16068 20720 16096
rect 20720 16050 20772 16056
rect 20456 15558 20576 15586
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20180 14742 20300 14770
rect 20272 14396 20300 14742
rect 20456 14550 20484 15558
rect 20824 15502 20852 17546
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20916 16182 20944 17206
rect 21008 16640 21036 18566
rect 21088 18148 21140 18154
rect 21088 18090 21140 18096
rect 21100 17241 21128 18090
rect 21192 17610 21220 19654
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21284 18834 21312 19246
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21086 17232 21142 17241
rect 21086 17167 21142 17176
rect 21008 16612 21220 16640
rect 21088 16516 21140 16522
rect 21088 16458 21140 16464
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20994 16144 21050 16153
rect 20994 16079 21050 16088
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20536 15496 20588 15502
rect 20812 15496 20864 15502
rect 20536 15438 20588 15444
rect 20626 15464 20682 15473
rect 20548 15094 20576 15438
rect 20810 15464 20812 15473
rect 20864 15464 20866 15473
rect 20682 15422 20760 15450
rect 20626 15399 20682 15408
rect 20536 15088 20588 15094
rect 20536 15030 20588 15036
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20548 14482 20576 14826
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20180 14368 20300 14396
rect 20180 14328 20208 14368
rect 20180 14300 20209 14328
rect 20181 14260 20209 14300
rect 19996 14232 20116 14260
rect 20173 14232 20209 14260
rect 20260 14272 20312 14278
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19430 14104 19486 14113
rect 19574 14107 19882 14116
rect 19430 14039 19486 14048
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 18892 13382 19104 13410
rect 19168 13394 19196 13806
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18892 13161 18920 13262
rect 19076 13258 19104 13382
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 18878 13152 18934 13161
rect 18878 13087 18934 13096
rect 18984 12714 19012 13194
rect 19062 13152 19118 13161
rect 19062 13087 19118 13096
rect 19076 12782 19104 13087
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 19076 12458 19104 12718
rect 18892 12430 19104 12458
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11150 18828 12106
rect 18788 11144 18840 11150
rect 18786 11112 18788 11121
rect 18840 11112 18842 11121
rect 18786 11047 18842 11056
rect 18892 10996 18920 12430
rect 19168 12073 19196 12718
rect 19154 12064 19210 12073
rect 19154 11999 19210 12008
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18984 11626 19012 11834
rect 19076 11801 19104 11834
rect 19062 11792 19118 11801
rect 19062 11727 19118 11736
rect 19062 11656 19118 11665
rect 18972 11620 19024 11626
rect 19260 11642 19288 13330
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19352 11830 19380 13194
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19118 11614 19288 11642
rect 19062 11591 19118 11600
rect 18972 11562 19024 11568
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 18800 10968 18920 10996
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18800 9042 18828 10968
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 18892 9897 18920 10678
rect 18878 9888 18934 9897
rect 18878 9823 18934 9832
rect 18984 9738 19012 11018
rect 19260 10985 19288 11086
rect 19246 10976 19302 10985
rect 19246 10911 19302 10920
rect 19352 10742 19380 11290
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19076 10198 19104 10542
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19168 9926 19196 10066
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19260 9738 19288 10678
rect 19338 9888 19394 9897
rect 19338 9823 19394 9832
rect 18892 9710 19012 9738
rect 19076 9710 19288 9738
rect 18892 9518 18920 9710
rect 19076 9674 19104 9710
rect 18984 9646 19104 9674
rect 19352 9654 19380 9823
rect 19248 9648 19300 9654
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18984 9466 19012 9646
rect 19248 9590 19300 9596
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 18984 9438 19196 9466
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18984 8906 19012 8978
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 18602 8800 18658 8809
rect 18602 8735 18658 8744
rect 18432 8622 18552 8650
rect 18432 8090 18460 8622
rect 18512 8560 18564 8566
rect 18564 8520 18828 8548
rect 18512 8502 18564 8508
rect 18696 8424 18748 8430
rect 18602 8392 18658 8401
rect 18696 8366 18748 8372
rect 18602 8327 18658 8336
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18524 8022 18552 8230
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18340 7772 18460 7800
rect 18326 7712 18382 7721
rect 18326 7647 18382 7656
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 18156 6934 18184 7210
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 18052 6860 18104 6866
rect 18340 6848 18368 7647
rect 18432 6914 18460 7772
rect 18510 7712 18566 7721
rect 18616 7698 18644 8327
rect 18708 8294 18736 8366
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18800 8072 18828 8520
rect 19076 8514 19104 8842
rect 18984 8486 19104 8514
rect 18878 8392 18934 8401
rect 18878 8327 18934 8336
rect 18892 8265 18920 8327
rect 18984 8294 19012 8486
rect 19064 8424 19116 8430
rect 19062 8392 19064 8401
rect 19116 8392 19118 8401
rect 19062 8327 19118 8336
rect 18984 8266 19104 8294
rect 18878 8256 18934 8265
rect 18878 8191 18934 8200
rect 18880 8084 18932 8090
rect 18800 8044 18880 8072
rect 18880 8026 18932 8032
rect 19076 7936 19104 8266
rect 18984 7908 19104 7936
rect 18616 7670 18920 7698
rect 18510 7647 18566 7656
rect 18524 7546 18552 7647
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18524 7274 18552 7346
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18616 7041 18644 7346
rect 18800 7206 18828 7482
rect 18892 7206 18920 7670
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18602 7032 18658 7041
rect 18602 6967 18658 6976
rect 18432 6886 18736 6914
rect 18340 6820 18552 6848
rect 18052 6802 18104 6808
rect 18418 6760 18474 6769
rect 18418 6695 18474 6704
rect 17972 6616 18092 6644
rect 17958 6488 18014 6497
rect 18064 6474 18092 6616
rect 18064 6446 18368 6474
rect 17958 6423 18014 6432
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17880 5642 17908 5714
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17788 4758 17816 5170
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 17788 4214 17816 4558
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17880 4146 17908 5034
rect 17972 4865 18000 6423
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18050 5944 18106 5953
rect 18050 5879 18106 5888
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3602 17816 3878
rect 18064 3738 18092 5879
rect 18156 5370 18184 6258
rect 18234 5808 18290 5817
rect 18234 5743 18290 5752
rect 18248 5710 18276 5743
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18156 5137 18184 5170
rect 18142 5128 18198 5137
rect 18248 5098 18276 5646
rect 18142 5063 18198 5072
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18340 4622 18368 6446
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18236 4208 18288 4214
rect 18156 4156 18236 4162
rect 18156 4150 18288 4156
rect 18156 4134 18276 4150
rect 18432 4146 18460 6695
rect 18420 4140 18472 4146
rect 18156 3942 18184 4134
rect 18420 4082 18472 4088
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17224 1964 17276 1970
rect 17224 1906 17276 1912
rect 17132 1692 17184 1698
rect 17132 1634 17184 1640
rect 17236 1630 17264 1906
rect 17224 1624 17276 1630
rect 17224 1566 17276 1572
rect 17328 1222 17356 3334
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17316 1216 17368 1222
rect 17316 1158 17368 1164
rect 17420 800 17448 2382
rect 17512 1737 17540 2790
rect 17788 2038 17816 3538
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 17498 1728 17554 1737
rect 17498 1663 17554 1672
rect 17972 1290 18000 3470
rect 18064 3058 18092 3470
rect 18248 3126 18276 3606
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18340 3058 18368 3878
rect 18432 3534 18460 3878
rect 18524 3738 18552 6820
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6633 18644 6734
rect 18602 6624 18658 6633
rect 18602 6559 18658 6568
rect 18616 6322 18644 6559
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18708 5914 18736 6886
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18786 6488 18842 6497
rect 18892 6458 18920 6734
rect 18786 6423 18842 6432
rect 18880 6452 18932 6458
rect 18800 6338 18828 6423
rect 18880 6394 18932 6400
rect 18800 6310 18920 6338
rect 18892 5914 18920 6310
rect 18696 5908 18748 5914
rect 18696 5850 18748 5856
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18708 5409 18736 5646
rect 18694 5400 18750 5409
rect 18694 5335 18750 5344
rect 18800 5216 18828 5646
rect 18708 5188 18828 5216
rect 18604 5160 18656 5166
rect 18708 5148 18736 5188
rect 18656 5120 18736 5148
rect 18604 5102 18656 5108
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18800 3369 18828 5034
rect 18786 3360 18842 3369
rect 18786 3295 18842 3304
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18892 2582 18920 5850
rect 18984 5030 19012 7908
rect 19062 7848 19118 7857
rect 19062 7783 19118 7792
rect 19076 7410 19104 7783
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 19076 6730 19104 6938
rect 19064 6724 19116 6730
rect 19064 6666 19116 6672
rect 19062 6624 19118 6633
rect 19062 6559 19118 6568
rect 19076 6322 19104 6559
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 19062 5536 19118 5545
rect 19062 5471 19118 5480
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18984 2825 19012 2994
rect 19076 2854 19104 5471
rect 19168 5302 19196 9438
rect 19260 8634 19288 9590
rect 19340 8900 19392 8906
rect 19444 8888 19472 13738
rect 19536 13258 19564 13738
rect 19904 13258 19932 13942
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19892 13252 19944 13258
rect 19892 13194 19944 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19720 12594 19748 12718
rect 19800 12708 19852 12714
rect 19996 12696 20024 14232
rect 20173 14090 20201 14232
rect 20260 14214 20312 14220
rect 20350 14240 20406 14249
rect 20076 14068 20128 14074
rect 20173 14062 20208 14090
rect 20076 14010 20128 14016
rect 19852 12668 20024 12696
rect 19800 12650 19852 12656
rect 19720 12566 20024 12594
rect 19996 12073 20024 12566
rect 19982 12064 20038 12073
rect 19574 11996 19882 12005
rect 19982 11999 20038 12008
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19628 11762 19656 11834
rect 19800 11824 19852 11830
rect 19720 11784 19800 11812
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19536 11082 19564 11698
rect 19628 11150 19656 11698
rect 19720 11354 19748 11784
rect 19800 11766 19852 11772
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19800 11280 19852 11286
rect 19984 11280 20036 11286
rect 19852 11240 19984 11268
rect 19800 11222 19852 11228
rect 19984 11222 20036 11228
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19984 11076 20036 11082
rect 19984 11018 20036 11024
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10792 20024 11018
rect 19904 10764 20024 10792
rect 19904 10248 19932 10764
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19812 10220 19932 10248
rect 19812 10044 19840 10220
rect 19892 10056 19944 10062
rect 19812 10016 19892 10044
rect 19892 9998 19944 10004
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19708 9648 19760 9654
rect 19760 9608 19840 9636
rect 19708 9590 19760 9596
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19628 9178 19656 9386
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19720 9081 19748 9454
rect 19812 9450 19840 9608
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19706 9072 19762 9081
rect 19706 9007 19762 9016
rect 19996 8974 20024 10542
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19392 8860 19472 8888
rect 19340 8842 19392 8848
rect 19536 8820 19564 8910
rect 20088 8820 20116 14010
rect 20180 11898 20208 14062
rect 20272 13410 20300 14214
rect 20350 14175 20406 14184
rect 20364 13705 20392 14175
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20350 13696 20406 13705
rect 20350 13631 20406 13640
rect 20272 13382 20392 13410
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20272 11393 20300 13262
rect 20364 12345 20392 13382
rect 20350 12336 20406 12345
rect 20350 12271 20406 12280
rect 20258 11384 20314 11393
rect 20258 11319 20314 11328
rect 20456 11200 20484 13874
rect 20640 13841 20668 13942
rect 20626 13832 20682 13841
rect 20626 13767 20682 13776
rect 20536 13456 20588 13462
rect 20536 13398 20588 13404
rect 20548 13258 20576 13398
rect 20626 13288 20682 13297
rect 20536 13252 20588 13258
rect 20626 13223 20682 13232
rect 20536 13194 20588 13200
rect 20640 12918 20668 13223
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20180 11172 20484 11200
rect 20180 11082 20208 11172
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20260 11076 20312 11082
rect 20260 11018 20312 11024
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 20180 9625 20208 10678
rect 20166 9616 20222 9625
rect 20166 9551 20222 9560
rect 20272 9500 20300 11018
rect 20350 10976 20406 10985
rect 20350 10911 20406 10920
rect 20364 10674 20392 10911
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 19444 8792 19564 8820
rect 19996 8792 20116 8820
rect 20180 9472 20300 9500
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19444 8514 19472 8792
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19260 8486 19472 8514
rect 19260 8004 19288 8486
rect 19996 8412 20024 8792
rect 20180 8650 20208 9472
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20173 8622 20208 8650
rect 20272 8634 20300 8842
rect 20364 8650 20392 10406
rect 20456 10130 20484 11172
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20456 9897 20484 10066
rect 20442 9888 20498 9897
rect 20442 9823 20498 9832
rect 20548 9432 20576 12854
rect 20732 12832 20760 15422
rect 20810 15399 20866 15408
rect 20824 15373 20852 15399
rect 20916 15337 20944 15982
rect 20902 15328 20958 15337
rect 20902 15263 20958 15272
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20824 13682 20852 15030
rect 20916 14793 20944 15030
rect 20902 14784 20958 14793
rect 20902 14719 20958 14728
rect 20902 14512 20958 14521
rect 21008 14498 21036 16079
rect 21100 14521 21128 16458
rect 20958 14470 21036 14498
rect 21086 14512 21142 14521
rect 20902 14447 20958 14456
rect 21086 14447 21142 14456
rect 21192 14362 21220 16612
rect 21284 16153 21312 18634
rect 21376 18154 21404 19944
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21468 18222 21496 18362
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21376 17513 21404 17750
rect 21362 17504 21418 17513
rect 21362 17439 21418 17448
rect 21362 17096 21418 17105
rect 21362 17031 21418 17040
rect 21376 16833 21404 17031
rect 21362 16824 21418 16833
rect 21362 16759 21418 16768
rect 21560 16232 21588 21490
rect 21652 20346 21680 22063
rect 21744 20466 21772 31726
rect 22112 30190 22140 33934
rect 22560 32564 22612 32570
rect 22560 32506 22612 32512
rect 22572 30326 22600 32506
rect 22560 30320 22612 30326
rect 22560 30262 22612 30268
rect 22100 30184 22152 30190
rect 22100 30126 22152 30132
rect 21916 28688 21968 28694
rect 21916 28630 21968 28636
rect 21928 28558 21956 28630
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 22098 28520 22154 28529
rect 22098 28455 22154 28464
rect 22112 28150 22140 28455
rect 22100 28144 22152 28150
rect 22100 28086 22152 28092
rect 22468 28008 22520 28014
rect 22468 27950 22520 27956
rect 21916 27600 21968 27606
rect 21916 27542 21968 27548
rect 21928 26926 21956 27542
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 21916 26920 21968 26926
rect 21916 26862 21968 26868
rect 21824 26852 21876 26858
rect 21824 26794 21876 26800
rect 21836 26738 21864 26794
rect 21836 26710 21956 26738
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21836 24206 21864 25842
rect 21928 24342 21956 26710
rect 22020 26217 22048 26930
rect 22388 26586 22416 27338
rect 22480 27062 22508 27950
rect 22756 27146 22784 37402
rect 23216 37244 23244 39200
rect 23216 37216 23520 37244
rect 23492 36922 23520 37216
rect 24504 37126 24532 39200
rect 24584 37256 24636 37262
rect 24584 37198 24636 37204
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 22836 30660 22888 30666
rect 22836 30602 22888 30608
rect 22848 29850 22876 30602
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 23400 28762 23428 36722
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 24504 36174 24532 36314
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 23572 33924 23624 33930
rect 23572 33866 23624 33872
rect 23584 29238 23612 33866
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23676 33522 23704 33798
rect 23664 33516 23716 33522
rect 23664 33458 23716 33464
rect 24504 29646 24532 36110
rect 24596 33658 24624 37198
rect 25148 37126 25176 39200
rect 25320 37256 25372 37262
rect 25320 37198 25372 37204
rect 26240 37256 26292 37262
rect 26240 37198 26292 37204
rect 25136 37120 25188 37126
rect 25136 37062 25188 37068
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 24780 33998 24808 36858
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 25332 33153 25360 37198
rect 26252 35894 26280 37198
rect 26436 37126 26464 39200
rect 27080 37194 27108 39200
rect 27528 37256 27580 37262
rect 27528 37198 27580 37204
rect 26976 37188 27028 37194
rect 26976 37130 27028 37136
rect 27068 37188 27120 37194
rect 27068 37130 27120 37136
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 26988 36786 27016 37130
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 26252 35866 26372 35894
rect 25318 33144 25374 33153
rect 25318 33079 25374 33088
rect 25320 32768 25372 32774
rect 25320 32710 25372 32716
rect 25332 30598 25360 32710
rect 25320 30592 25372 30598
rect 25320 30534 25372 30540
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 24032 29504 24084 29510
rect 24032 29446 24084 29452
rect 23952 29238 23980 29446
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23664 29232 23716 29238
rect 23664 29174 23716 29180
rect 23940 29232 23992 29238
rect 23940 29174 23992 29180
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 23676 28234 23704 29174
rect 23940 29096 23992 29102
rect 23940 29038 23992 29044
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23676 28218 23796 28234
rect 23676 28212 23808 28218
rect 23676 28206 23756 28212
rect 23756 28154 23808 28160
rect 22756 27118 22876 27146
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22744 27056 22796 27062
rect 22744 26998 22796 27004
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22204 26450 22232 26522
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22112 26330 22140 26386
rect 22284 26376 22336 26382
rect 22112 26302 22232 26330
rect 22284 26318 22336 26324
rect 22006 26208 22062 26217
rect 22006 26143 22062 26152
rect 22204 25702 22232 26302
rect 22296 25809 22324 26318
rect 22282 25800 22338 25809
rect 22282 25735 22338 25744
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 22204 25362 22232 25638
rect 22296 25498 22324 25735
rect 22480 25673 22508 26998
rect 22756 26042 22784 26998
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22652 25764 22704 25770
rect 22652 25706 22704 25712
rect 22466 25664 22522 25673
rect 22466 25599 22522 25608
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22192 25356 22244 25362
rect 22192 25298 22244 25304
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21836 23338 21864 23802
rect 21928 23497 21956 24006
rect 21914 23488 21970 23497
rect 21914 23423 21970 23432
rect 21836 23310 22048 23338
rect 22020 23186 22048 23310
rect 22008 23180 22060 23186
rect 22008 23122 22060 23128
rect 21914 23080 21970 23089
rect 21914 23015 21916 23024
rect 21968 23015 21970 23024
rect 21916 22986 21968 22992
rect 21822 22672 21878 22681
rect 21822 22607 21878 22616
rect 21836 20505 21864 22607
rect 21928 22506 21956 22986
rect 22112 22778 22140 24142
rect 22100 22772 22152 22778
rect 22100 22714 22152 22720
rect 22204 22506 22232 25298
rect 22284 25220 22336 25226
rect 22284 25162 22336 25168
rect 22296 24954 22324 25162
rect 22284 24948 22336 24954
rect 22284 24890 22336 24896
rect 22282 24712 22338 24721
rect 22282 24647 22338 24656
rect 22296 24614 22324 24647
rect 22284 24608 22336 24614
rect 22284 24550 22336 24556
rect 22388 24342 22416 25298
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 22388 24206 22416 24278
rect 22376 24200 22428 24206
rect 22376 24142 22428 24148
rect 22284 23792 22336 23798
rect 22480 23769 22508 25162
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22284 23734 22336 23740
rect 22466 23760 22522 23769
rect 21916 22500 21968 22506
rect 21916 22442 21968 22448
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22296 22098 22324 23734
rect 22466 23695 22522 23704
rect 22376 23588 22428 23594
rect 22376 23530 22428 23536
rect 22388 22574 22416 23530
rect 22480 22930 22508 23695
rect 22572 23050 22600 24006
rect 22560 23044 22612 23050
rect 22664 23032 22692 25706
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 22756 23662 22784 24618
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22744 23044 22796 23050
rect 22664 23004 22744 23032
rect 22560 22986 22612 22992
rect 22744 22986 22796 22992
rect 22480 22902 22692 22930
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 21914 21720 21970 21729
rect 21914 21655 21970 21664
rect 21928 21622 21956 21655
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21822 20496 21878 20505
rect 21732 20460 21784 20466
rect 21822 20431 21878 20440
rect 21732 20402 21784 20408
rect 21824 20392 21876 20398
rect 21652 20318 21772 20346
rect 21824 20334 21876 20340
rect 21640 19848 21692 19854
rect 21640 19790 21692 19796
rect 21652 19689 21680 19790
rect 21638 19680 21694 19689
rect 21638 19615 21694 19624
rect 21640 19236 21692 19242
rect 21640 19178 21692 19184
rect 21652 18465 21680 19178
rect 21638 18456 21694 18465
rect 21638 18391 21694 18400
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21376 16204 21588 16232
rect 21270 16144 21326 16153
rect 21270 16079 21326 16088
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21008 14334 21220 14362
rect 21008 13938 21036 14334
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 13864 20956 13870
rect 20902 13832 20904 13841
rect 20956 13832 20958 13841
rect 20902 13767 20958 13776
rect 21100 13784 21128 14214
rect 21192 14074 21220 14214
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21100 13756 21220 13784
rect 21086 13696 21142 13705
rect 20824 13654 20944 13682
rect 20916 13530 20944 13654
rect 21086 13631 21142 13640
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20824 13326 20852 13466
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20902 13288 20958 13297
rect 20902 13223 20958 13232
rect 20916 13190 20944 13223
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20732 12804 20852 12832
rect 20824 12714 20852 12804
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20626 12064 20682 12073
rect 20626 11999 20682 12008
rect 20640 11762 20668 11999
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20732 11506 20760 12650
rect 20904 12368 20956 12374
rect 20810 12336 20866 12345
rect 20904 12310 20956 12316
rect 20810 12271 20866 12280
rect 20824 11608 20852 12271
rect 20916 12170 20944 12310
rect 20904 12164 20956 12170
rect 20904 12106 20956 12112
rect 20902 12064 20958 12073
rect 20902 11999 20958 12008
rect 20916 11801 20944 11999
rect 21008 11898 21036 13330
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21100 11830 21128 13631
rect 21192 12782 21220 13756
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 21088 11824 21140 11830
rect 20902 11792 20958 11801
rect 21088 11766 21140 11772
rect 20902 11727 20958 11736
rect 20824 11580 21128 11608
rect 20732 11478 20852 11506
rect 20718 11384 20774 11393
rect 20718 11319 20774 11328
rect 20628 11212 20680 11218
rect 20732 11200 20760 11319
rect 20680 11172 20760 11200
rect 20628 11154 20680 11160
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 10742 20760 11018
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20628 10600 20680 10606
rect 20824 10588 20852 11478
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 20916 10724 20944 11290
rect 20916 10696 21036 10724
rect 21008 10606 21036 10696
rect 20628 10542 20680 10548
rect 20732 10560 20852 10588
rect 20996 10600 21048 10606
rect 20640 10441 20668 10542
rect 20626 10432 20682 10441
rect 20626 10367 20682 10376
rect 20626 9888 20682 9897
rect 20732 9874 20760 10560
rect 20996 10542 21048 10548
rect 20994 10432 21050 10441
rect 20994 10367 21050 10376
rect 20810 10296 20866 10305
rect 20810 10231 20866 10240
rect 20824 10062 20852 10231
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20626 9823 20682 9832
rect 20724 9846 20760 9874
rect 20640 9500 20668 9823
rect 20724 9738 20752 9846
rect 20724 9710 20944 9738
rect 20916 9586 20944 9710
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20640 9472 20852 9500
rect 20456 9404 20576 9432
rect 20456 8820 20484 9404
rect 20718 9208 20774 9217
rect 20628 9172 20680 9178
rect 20718 9143 20720 9152
rect 20628 9114 20680 9120
rect 20772 9143 20774 9152
rect 20720 9114 20772 9120
rect 20456 8792 20576 8820
rect 20260 8628 20312 8634
rect 20173 8480 20201 8622
rect 20364 8622 20484 8650
rect 20260 8570 20312 8576
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20173 8452 20208 8480
rect 19904 8384 20024 8412
rect 19800 8356 19852 8362
rect 19444 8316 19800 8344
rect 19340 8288 19392 8294
rect 19444 8242 19472 8316
rect 19800 8298 19852 8304
rect 19392 8236 19472 8242
rect 19340 8230 19472 8236
rect 19352 8214 19472 8230
rect 19260 7976 19334 8004
rect 19306 7936 19334 7976
rect 19904 7954 19932 8384
rect 19982 8256 20038 8265
rect 19982 8191 20038 8200
rect 19996 7970 20024 8191
rect 19260 7908 19334 7936
rect 19892 7948 19944 7954
rect 19260 7460 19288 7908
rect 19996 7942 20116 7970
rect 19892 7890 19944 7896
rect 19616 7812 19668 7818
rect 19444 7772 19616 7800
rect 19444 7721 19472 7772
rect 19616 7754 19668 7760
rect 19984 7744 20036 7750
rect 19430 7712 19486 7721
rect 19984 7686 20036 7692
rect 19430 7647 19486 7656
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19260 7432 19380 7460
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19260 6458 19288 6802
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19156 5296 19208 5302
rect 19156 5238 19208 5244
rect 19260 5098 19288 6054
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19352 4978 19380 7432
rect 19996 7290 20024 7686
rect 20088 7410 20116 7942
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19996 7262 20116 7290
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19996 7041 20024 7142
rect 19982 7032 20038 7041
rect 20088 7002 20116 7262
rect 19982 6967 20038 6976
rect 20076 6996 20128 7002
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19432 6656 19484 6662
rect 19628 6644 19656 6734
rect 19484 6616 19656 6644
rect 19432 6598 19484 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19708 6452 19760 6458
rect 19760 6412 19932 6440
rect 19708 6394 19760 6400
rect 19614 6352 19670 6361
rect 19614 6287 19616 6296
rect 19668 6287 19670 6296
rect 19798 6352 19854 6361
rect 19798 6287 19854 6296
rect 19616 6258 19668 6264
rect 19430 5808 19486 5817
rect 19812 5778 19840 6287
rect 19904 5778 19932 6412
rect 19996 6322 20024 6967
rect 20076 6938 20128 6944
rect 20180 6866 20208 8452
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20272 6746 20300 7958
rect 20088 6718 20300 6746
rect 20088 6390 20116 6718
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20258 6352 20314 6361
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 20180 6118 20208 6326
rect 20258 6287 20260 6296
rect 20312 6287 20314 6296
rect 20260 6258 20312 6264
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20364 5914 20392 8502
rect 20456 6474 20484 8622
rect 20548 6662 20576 8792
rect 20640 7274 20668 9114
rect 20824 8906 20852 9472
rect 20902 9480 20958 9489
rect 20902 9415 20958 9424
rect 20916 9382 20944 9415
rect 20904 9376 20956 9382
rect 21008 9353 21036 10367
rect 21100 10169 21128 11580
rect 21192 11354 21220 12310
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21086 10160 21142 10169
rect 21086 10095 21142 10104
rect 21100 10062 21128 10095
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21180 9920 21232 9926
rect 21086 9888 21142 9897
rect 21180 9862 21232 9868
rect 21086 9823 21142 9832
rect 20904 9318 20956 9324
rect 20994 9344 21050 9353
rect 20994 9279 21050 9288
rect 21100 8945 21128 9823
rect 21192 9654 21220 9862
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21178 9208 21234 9217
rect 21178 9143 21180 9152
rect 21232 9143 21234 9152
rect 21180 9114 21232 9120
rect 21086 8936 21142 8945
rect 20812 8900 20864 8906
rect 21086 8871 21142 8880
rect 21180 8900 21232 8906
rect 20812 8842 20864 8848
rect 21180 8842 21232 8848
rect 20902 8800 20958 8809
rect 20902 8735 20958 8744
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20732 8022 20760 8191
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20718 7712 20774 7721
rect 20718 7647 20774 7656
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20732 6798 20760 7647
rect 20824 7478 20852 8434
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20812 6724 20864 6730
rect 20812 6666 20864 6672
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20626 6624 20682 6633
rect 20626 6559 20682 6568
rect 20456 6446 20576 6474
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20456 6118 20484 6258
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 19996 5817 20024 5850
rect 19982 5808 20038 5817
rect 19430 5743 19486 5752
rect 19800 5772 19852 5778
rect 19444 5352 19472 5743
rect 19800 5714 19852 5720
rect 19892 5772 19944 5778
rect 20456 5794 20484 6054
rect 19982 5743 20038 5752
rect 20364 5766 20484 5794
rect 19892 5714 19944 5720
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20088 5574 20116 5646
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19982 5400 20038 5409
rect 19444 5324 19656 5352
rect 19982 5335 20038 5344
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19260 4950 19380 4978
rect 19154 4448 19210 4457
rect 19154 4383 19210 4392
rect 19168 3942 19196 4383
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 19168 3233 19196 3674
rect 19260 3534 19288 4950
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19352 4264 19380 4558
rect 19444 4486 19472 5102
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4554 19564 4966
rect 19628 4622 19656 5324
rect 19996 5030 20024 5335
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 19432 4480 19484 4486
rect 19432 4422 19484 4428
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4276 19484 4282
rect 19352 4236 19432 4264
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19154 3224 19210 3233
rect 19154 3159 19210 3168
rect 19156 3052 19208 3058
rect 19156 2994 19208 3000
rect 19064 2848 19116 2854
rect 18970 2816 19026 2825
rect 19064 2790 19116 2796
rect 18970 2751 19026 2760
rect 19168 2650 19196 2994
rect 19260 2650 19288 3334
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 19062 2544 19118 2553
rect 19062 2479 19118 2488
rect 19246 2544 19302 2553
rect 19352 2514 19380 4236
rect 19432 4218 19484 4224
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19444 2650 19472 4082
rect 19536 4049 19564 4082
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 19890 4040 19946 4049
rect 19996 4010 20024 4422
rect 19890 3975 19946 3984
rect 19984 4004 20036 4010
rect 19904 3738 19932 3975
rect 19984 3946 20036 3952
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19984 3392 20036 3398
rect 20180 3346 20208 4490
rect 20272 3505 20300 5170
rect 20258 3496 20314 3505
rect 20258 3431 20314 3440
rect 19984 3334 20036 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19246 2479 19302 2488
rect 19340 2508 19392 2514
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 17960 1284 18012 1290
rect 17960 1226 18012 1232
rect 18708 800 18736 2382
rect 19076 2038 19104 2479
rect 19260 2145 19288 2479
rect 19340 2450 19392 2456
rect 19536 2292 19564 3130
rect 19996 3058 20024 3334
rect 20088 3318 20208 3346
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19352 2264 19564 2292
rect 19246 2136 19302 2145
rect 19246 2071 19302 2080
rect 19064 2032 19116 2038
rect 19064 1974 19116 1980
rect 19352 800 19380 2264
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2382
rect 20088 2038 20116 3318
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 20180 2106 20208 3130
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 20076 2032 20128 2038
rect 20076 1974 20128 1980
rect 20272 1873 20300 3431
rect 20364 2514 20392 5766
rect 20548 5216 20576 6446
rect 20640 5794 20668 6559
rect 20824 6497 20852 6666
rect 20810 6488 20866 6497
rect 20810 6423 20866 6432
rect 20916 6390 20944 8735
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21100 7886 21128 8230
rect 21192 8129 21220 8842
rect 21178 8120 21234 8129
rect 21178 8055 21234 8064
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21088 7880 21140 7886
rect 20994 7848 21050 7857
rect 21088 7822 21140 7828
rect 21192 7818 21220 7890
rect 20994 7783 21050 7792
rect 21180 7812 21232 7818
rect 21008 7750 21036 7783
rect 21180 7754 21232 7760
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 21088 7268 21140 7274
rect 21088 7210 21140 7216
rect 20996 6792 21048 6798
rect 21100 6769 21128 7210
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 20996 6734 21048 6740
rect 21086 6760 21142 6769
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20732 5914 20760 6326
rect 21008 6186 21036 6734
rect 21086 6695 21142 6704
rect 21192 6458 21220 6802
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21180 6316 21232 6322
rect 21100 6276 21180 6304
rect 20996 6180 21048 6186
rect 20996 6122 21048 6128
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20994 5808 21050 5817
rect 20640 5766 20944 5794
rect 20812 5704 20864 5710
rect 20810 5672 20812 5681
rect 20864 5672 20866 5681
rect 20810 5607 20866 5616
rect 20718 5536 20774 5545
rect 20718 5471 20774 5480
rect 20548 5188 20668 5216
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20456 2378 20484 4966
rect 20548 2417 20576 5034
rect 20640 4486 20668 5188
rect 20732 4593 20760 5471
rect 20916 5409 20944 5766
rect 20994 5743 21050 5752
rect 21008 5710 21036 5743
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20902 5400 20958 5409
rect 20902 5335 20958 5344
rect 20810 5264 20866 5273
rect 20810 5199 20866 5208
rect 20824 5166 20852 5199
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20812 4616 20864 4622
rect 20718 4584 20774 4593
rect 20812 4558 20864 4564
rect 20718 4519 20774 4528
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20732 4214 20760 4422
rect 20720 4208 20772 4214
rect 20626 4176 20682 4185
rect 20720 4150 20772 4156
rect 20626 4111 20682 4120
rect 20640 3738 20668 4111
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20626 3632 20682 3641
rect 20626 3567 20682 3576
rect 20640 3534 20668 3567
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20534 2408 20590 2417
rect 20444 2372 20496 2378
rect 20534 2343 20590 2352
rect 20444 2314 20496 2320
rect 20258 1864 20314 1873
rect 20258 1799 20314 1808
rect 20732 1358 20760 3878
rect 20824 2310 20852 4558
rect 21100 4554 21128 6276
rect 21180 6258 21232 6264
rect 21178 5808 21234 5817
rect 21178 5743 21180 5752
rect 21232 5743 21234 5752
rect 21180 5714 21232 5720
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20916 2922 20944 4082
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21008 3058 21036 3878
rect 21192 3534 21220 4558
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 21100 2582 21128 3402
rect 21284 2774 21312 15302
rect 21376 15065 21404 16204
rect 21546 16144 21602 16153
rect 21546 16079 21602 16088
rect 21560 15688 21588 16079
rect 21652 16046 21680 18158
rect 21744 16833 21772 20318
rect 21836 17082 21864 20334
rect 21928 18873 21956 20946
rect 22020 20398 22048 21490
rect 22112 21486 22140 21898
rect 22204 21570 22232 21966
rect 22204 21542 22324 21570
rect 22100 21480 22152 21486
rect 22192 21480 22244 21486
rect 22100 21422 22152 21428
rect 22190 21448 22192 21457
rect 22244 21448 22246 21457
rect 22190 21383 22246 21392
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22204 21146 22232 21286
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22296 21026 22324 21542
rect 22572 21400 22600 22510
rect 22664 21978 22692 22902
rect 22756 22817 22784 22986
rect 22742 22808 22798 22817
rect 22742 22743 22798 22752
rect 22848 22094 22876 27118
rect 23296 27056 23348 27062
rect 23296 26998 23348 27004
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 22940 22234 22968 26318
rect 23018 26208 23074 26217
rect 23018 26143 23074 26152
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 22848 22066 22968 22094
rect 22664 21950 22784 21978
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21729 22692 21830
rect 22650 21720 22706 21729
rect 22650 21655 22706 21664
rect 22572 21372 22692 21400
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22558 21312 22614 21321
rect 22112 20998 22324 21026
rect 22112 20942 22140 20998
rect 22100 20936 22152 20942
rect 22480 20890 22508 21286
rect 22558 21247 22614 21256
rect 22572 20942 22600 21247
rect 22100 20878 22152 20884
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22008 18896 22060 18902
rect 21914 18864 21970 18873
rect 22008 18838 22060 18844
rect 21914 18799 21970 18808
rect 22020 18290 22048 18838
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 22112 18222 22140 20878
rect 22296 20862 22508 20890
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 19514 22232 20742
rect 22296 20398 22324 20862
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22388 20534 22416 20742
rect 22376 20528 22428 20534
rect 22468 20528 22520 20534
rect 22376 20470 22428 20476
rect 22466 20496 22468 20505
rect 22520 20496 22522 20505
rect 22466 20431 22522 20440
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22374 20360 22430 20369
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 22296 19122 22324 20334
rect 22374 20295 22430 20304
rect 22558 20360 22614 20369
rect 22558 20295 22614 20304
rect 22388 19961 22416 20295
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22374 19952 22430 19961
rect 22374 19887 22430 19896
rect 22480 19786 22508 19994
rect 22572 19786 22600 20295
rect 22468 19780 22520 19786
rect 22468 19722 22520 19728
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22480 19446 22508 19722
rect 22468 19440 22520 19446
rect 22468 19382 22520 19388
rect 22296 19094 22508 19122
rect 22480 18834 22508 19094
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22480 18358 22508 18770
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21916 17808 21968 17814
rect 21916 17750 21968 17756
rect 21928 17202 21956 17750
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17377 22140 17478
rect 22296 17377 22324 17614
rect 22572 17513 22600 17614
rect 22558 17504 22614 17513
rect 22558 17439 22614 17448
rect 22098 17368 22154 17377
rect 22098 17303 22154 17312
rect 22282 17368 22338 17377
rect 22282 17303 22338 17312
rect 22192 17264 22244 17270
rect 22244 17224 22416 17252
rect 22192 17206 22244 17212
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 21836 17054 21956 17082
rect 21730 16824 21786 16833
rect 21730 16759 21786 16768
rect 21928 16674 21956 17054
rect 22098 16824 22154 16833
rect 22098 16759 22154 16768
rect 22282 16824 22338 16833
rect 22282 16759 22338 16768
rect 21744 16646 21956 16674
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21560 15660 21680 15688
rect 21546 15600 21602 15609
rect 21546 15535 21602 15544
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21362 15056 21418 15065
rect 21362 14991 21418 15000
rect 21376 12238 21404 14991
rect 21468 13530 21496 15370
rect 21560 14906 21588 15535
rect 21652 15026 21680 15660
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21560 14878 21680 14906
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21560 14521 21588 14554
rect 21652 14532 21680 14878
rect 21744 14657 21772 16646
rect 22112 16574 22140 16759
rect 22190 16688 22246 16697
rect 22296 16658 22324 16759
rect 22190 16623 22246 16632
rect 22284 16652 22336 16658
rect 21836 16546 22140 16574
rect 21836 15978 21864 16546
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22112 16182 22140 16390
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21824 15972 21876 15978
rect 21824 15914 21876 15920
rect 21928 15552 21956 15982
rect 22112 15706 22140 15982
rect 22204 15706 22232 16623
rect 22284 16594 22336 16600
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22284 15564 22336 15570
rect 21928 15524 22284 15552
rect 22284 15506 22336 15512
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 21916 15088 21968 15094
rect 21914 15056 21916 15065
rect 21968 15056 21970 15065
rect 21914 14991 21970 15000
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21730 14648 21786 14657
rect 21730 14583 21786 14592
rect 21546 14512 21602 14521
rect 21652 14504 21772 14532
rect 21546 14447 21602 14456
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 14006 21588 14282
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21652 13394 21680 14350
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21744 13274 21772 14504
rect 21836 14278 21864 14894
rect 22020 14600 22048 15302
rect 22204 15094 22232 15302
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22388 14958 22416 17224
rect 22664 17134 22692 21372
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22756 16658 22784 21950
rect 22834 21584 22890 21593
rect 22834 21519 22890 21528
rect 22940 21536 22968 22066
rect 23032 22001 23060 26143
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23018 21992 23074 22001
rect 23018 21927 23074 21936
rect 23032 21729 23060 21927
rect 23018 21720 23074 21729
rect 23018 21655 23074 21664
rect 23020 21548 23072 21554
rect 22848 20942 22876 21519
rect 22940 21508 23020 21536
rect 23020 21490 23072 21496
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 22940 20505 22968 20946
rect 23032 20874 23060 21490
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 22926 20496 22982 20505
rect 22926 20431 22982 20440
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22928 20324 22980 20330
rect 22928 20266 22980 20272
rect 22848 17921 22876 20266
rect 22940 19786 22968 20266
rect 23032 20262 23060 20402
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22928 18828 22980 18834
rect 22980 18788 23060 18816
rect 22928 18770 22980 18776
rect 23032 17921 23060 18788
rect 22834 17912 22890 17921
rect 22834 17847 22890 17856
rect 23018 17912 23074 17921
rect 23018 17847 23074 17856
rect 22848 17513 22876 17847
rect 22834 17504 22890 17513
rect 22834 17439 22890 17448
rect 22848 17202 22876 17439
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22940 16697 22968 16730
rect 22926 16688 22982 16697
rect 22744 16652 22796 16658
rect 22926 16623 22982 16632
rect 22744 16594 22796 16600
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22848 16454 22876 16526
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22744 15632 22796 15638
rect 22742 15600 22744 15609
rect 22796 15600 22798 15609
rect 22742 15535 22798 15544
rect 23032 15552 23060 17847
rect 23124 17678 23152 25842
rect 23216 24954 23244 26386
rect 23204 24948 23256 24954
rect 23204 24890 23256 24896
rect 23216 24410 23244 24890
rect 23204 24404 23256 24410
rect 23204 24346 23256 24352
rect 23216 23798 23244 24346
rect 23204 23792 23256 23798
rect 23204 23734 23256 23740
rect 23308 22545 23336 26998
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23400 26042 23428 26182
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23756 25832 23808 25838
rect 23756 25774 23808 25780
rect 23480 24880 23532 24886
rect 23480 24822 23532 24828
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23400 24274 23428 24686
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23294 22536 23350 22545
rect 23294 22471 23350 22480
rect 23400 22438 23428 23258
rect 23388 22432 23440 22438
rect 23202 22400 23258 22409
rect 23388 22374 23440 22380
rect 23202 22335 23258 22344
rect 23216 21962 23244 22335
rect 23294 22128 23350 22137
rect 23294 22063 23350 22072
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23202 21720 23258 21729
rect 23202 21655 23258 21664
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23112 17264 23164 17270
rect 23112 17206 23164 17212
rect 23124 16794 23152 17206
rect 23216 17202 23244 21655
rect 23308 21457 23336 22063
rect 23388 21956 23440 21962
rect 23388 21898 23440 21904
rect 23294 21448 23350 21457
rect 23294 21383 23350 21392
rect 23308 17678 23336 21383
rect 23400 20058 23428 21898
rect 23492 21690 23520 24822
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23676 23866 23704 24074
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23584 23361 23612 23666
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23570 23352 23626 23361
rect 23570 23287 23626 23296
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23584 22216 23612 22986
rect 23676 22710 23704 23462
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23584 22188 23704 22216
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23492 20466 23520 21490
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23400 19718 23428 19994
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23492 18766 23520 20198
rect 23584 19666 23612 22034
rect 23676 20058 23704 22188
rect 23768 22098 23796 25774
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23860 21672 23888 28494
rect 23952 23798 23980 29038
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 22234 23980 22646
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23768 21644 23888 21672
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23768 19938 23796 21644
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 21078 23888 21490
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23938 20632 23994 20641
rect 23938 20567 23994 20576
rect 23848 20392 23900 20398
rect 23848 20334 23900 20340
rect 23676 19910 23796 19938
rect 23676 19786 23704 19910
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23584 19638 23704 19666
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23570 18320 23626 18329
rect 23570 18255 23626 18264
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23308 17105 23336 17478
rect 23294 17096 23350 17105
rect 23294 17031 23350 17040
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23216 16182 23244 16730
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23112 16040 23164 16046
rect 23110 16008 23112 16017
rect 23164 16008 23166 16017
rect 23110 15943 23166 15952
rect 23124 15745 23152 15943
rect 23110 15736 23166 15745
rect 23110 15671 23166 15680
rect 23032 15524 23152 15552
rect 22652 15496 22704 15502
rect 22466 15464 22522 15473
rect 22652 15438 22704 15444
rect 22466 15399 22522 15408
rect 22560 15428 22612 15434
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22282 14784 22338 14793
rect 22282 14719 22338 14728
rect 22100 14612 22152 14618
rect 22020 14572 22100 14600
rect 21824 14272 21876 14278
rect 22020 14249 22048 14572
rect 22100 14554 22152 14560
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 21824 14214 21876 14220
rect 22006 14240 22062 14249
rect 22006 14175 22062 14184
rect 21822 14104 21878 14113
rect 21822 14039 21878 14048
rect 21836 13938 21864 14039
rect 21916 14000 21968 14006
rect 22112 13954 22140 14350
rect 22296 14346 22324 14719
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22282 14104 22338 14113
rect 22282 14039 22284 14048
rect 22336 14039 22338 14048
rect 22284 14010 22336 14016
rect 21916 13942 21968 13948
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21836 13705 21864 13874
rect 21928 13734 21956 13942
rect 22020 13926 22140 13954
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 21916 13728 21968 13734
rect 21822 13696 21878 13705
rect 21916 13670 21968 13676
rect 21822 13631 21878 13640
rect 21560 13246 21772 13274
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21362 11656 21418 11665
rect 21362 11591 21418 11600
rect 21376 11150 21404 11591
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21376 8974 21404 11086
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21376 8634 21404 8774
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21362 8120 21418 8129
rect 21362 8055 21418 8064
rect 21376 7274 21404 8055
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21362 6216 21418 6225
rect 21362 6151 21364 6160
rect 21416 6151 21418 6160
rect 21364 6122 21416 6128
rect 21362 4720 21418 4729
rect 21362 4655 21418 4664
rect 21376 4554 21404 4655
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21468 4146 21496 12854
rect 21560 10742 21588 13246
rect 21914 13152 21970 13161
rect 21914 13087 21970 13096
rect 21928 12918 21956 13087
rect 21916 12912 21968 12918
rect 21730 12880 21786 12889
rect 21916 12854 21968 12860
rect 21730 12815 21732 12824
rect 21784 12815 21786 12824
rect 21732 12786 21784 12792
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21652 10266 21680 12650
rect 22020 12288 22048 13926
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 13705 22140 13806
rect 22098 13696 22154 13705
rect 22098 13631 22154 13640
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 21836 12260 22048 12288
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21744 11665 21772 11698
rect 21730 11656 21786 11665
rect 21730 11591 21786 11600
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21548 9648 21600 9654
rect 21546 9616 21548 9625
rect 21600 9616 21602 9625
rect 21546 9551 21602 9560
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21560 9382 21588 9454
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21548 9104 21600 9110
rect 21546 9072 21548 9081
rect 21600 9072 21602 9081
rect 21546 9007 21602 9016
rect 21652 8838 21680 9522
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21560 8129 21588 8366
rect 21546 8120 21602 8129
rect 21546 8055 21602 8064
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21560 7478 21588 7822
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21652 7410 21680 8774
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21744 7313 21772 11591
rect 21836 9994 21864 12260
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11898 21956 12038
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21914 11792 21970 11801
rect 21914 11727 21916 11736
rect 21968 11727 21970 11736
rect 21916 11698 21968 11704
rect 22020 11529 22048 12106
rect 22112 11830 22140 13330
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22006 11520 22062 11529
rect 22006 11455 22062 11464
rect 22204 11354 22232 13942
rect 22388 13841 22416 14282
rect 22480 13870 22508 15399
rect 22560 15370 22612 15376
rect 22572 14074 22600 15370
rect 22664 14482 22692 15438
rect 22928 15428 22980 15434
rect 22928 15370 22980 15376
rect 23020 15428 23072 15434
rect 23020 15370 23072 15376
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 14278 22784 14350
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22744 13932 22796 13938
rect 22572 13892 22744 13920
rect 22468 13864 22520 13870
rect 22374 13832 22430 13841
rect 22468 13806 22520 13812
rect 22374 13767 22430 13776
rect 22572 13716 22600 13892
rect 22744 13874 22796 13880
rect 22388 13688 22600 13716
rect 22650 13696 22706 13705
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22296 12986 22324 13330
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22388 12889 22416 13688
rect 22650 13631 22706 13640
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22374 12880 22430 12889
rect 22480 12866 22508 13126
rect 22572 12986 22600 13194
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22558 12880 22614 12889
rect 22480 12838 22558 12866
rect 22374 12815 22430 12824
rect 22558 12815 22614 12824
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22296 12306 22324 12650
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 22296 11234 22324 11766
rect 22112 11206 22324 11234
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22020 10810 22048 10950
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 22020 10146 22048 10610
rect 21928 10118 22048 10146
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21928 9897 21956 10118
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21914 9888 21970 9897
rect 21914 9823 21970 9832
rect 22020 9738 22048 9998
rect 21836 9710 22048 9738
rect 21836 8401 21864 9710
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21928 9178 21956 9590
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22006 8936 22062 8945
rect 22006 8871 22062 8880
rect 21914 8800 21970 8809
rect 21914 8735 21970 8744
rect 21928 8498 21956 8735
rect 21916 8492 21968 8498
rect 21916 8434 21968 8440
rect 22020 8401 22048 8871
rect 21822 8392 21878 8401
rect 21822 8327 21878 8336
rect 22006 8392 22062 8401
rect 22006 8327 22062 8336
rect 22020 7970 22048 8327
rect 22112 8106 22140 11206
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22204 9382 22232 11086
rect 22282 10432 22338 10441
rect 22282 10367 22338 10376
rect 22296 10130 22324 10367
rect 22388 10266 22416 12718
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22480 10674 22508 11630
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22296 9450 22324 9590
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 22204 9178 22232 9318
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22190 8936 22246 8945
rect 22190 8871 22246 8880
rect 22204 8362 22232 8871
rect 22388 8650 22416 9998
rect 22480 8945 22508 10406
rect 22466 8936 22522 8945
rect 22572 8906 22600 11222
rect 22664 9489 22692 13631
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22756 13025 22784 13262
rect 22742 13016 22798 13025
rect 22742 12951 22798 12960
rect 22744 12912 22796 12918
rect 22744 12854 22796 12860
rect 22756 10810 22784 12854
rect 22744 10804 22796 10810
rect 22744 10746 22796 10752
rect 22650 9480 22706 9489
rect 22706 9438 22784 9466
rect 22650 9415 22706 9424
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22664 8906 22692 9318
rect 22466 8871 22522 8880
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22296 8622 22416 8650
rect 22296 8412 22324 8622
rect 22376 8560 22428 8566
rect 22428 8520 22508 8548
rect 22376 8502 22428 8508
rect 22296 8384 22416 8412
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22112 8078 22232 8106
rect 21836 7942 22048 7970
rect 22098 7984 22154 7993
rect 21730 7304 21786 7313
rect 21730 7239 21786 7248
rect 21836 6322 21864 7942
rect 22098 7919 22154 7928
rect 22112 7886 22140 7919
rect 22008 7880 22060 7886
rect 21914 7848 21970 7857
rect 22008 7822 22060 7828
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21914 7783 21970 7792
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21744 5658 21772 5850
rect 21560 5630 21772 5658
rect 21560 5250 21588 5630
rect 21836 5534 21864 6258
rect 21928 5778 21956 7783
rect 22020 7206 22048 7822
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22098 7032 22154 7041
rect 22098 6967 22154 6976
rect 22006 6896 22062 6905
rect 22006 6831 22062 6840
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 22020 5574 22048 6831
rect 22112 6798 22140 6967
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 21744 5506 21864 5534
rect 22008 5568 22060 5574
rect 22008 5510 22060 5516
rect 21560 5222 21680 5250
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21362 3768 21418 3777
rect 21362 3703 21418 3712
rect 21376 3534 21404 3703
rect 21652 3652 21680 5222
rect 21744 4049 21772 5506
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21836 4622 21864 5170
rect 22112 4978 22140 6598
rect 22204 5794 22232 8078
rect 22282 7304 22338 7313
rect 22282 7239 22338 7248
rect 22296 6934 22324 7239
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22282 6488 22338 6497
rect 22282 6423 22284 6432
rect 22336 6423 22338 6432
rect 22284 6394 22336 6400
rect 22388 6225 22416 8384
rect 22480 8090 22508 8520
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22466 7984 22522 7993
rect 22466 7919 22522 7928
rect 22480 6390 22508 7919
rect 22468 6384 22520 6390
rect 22468 6326 22520 6332
rect 22572 6254 22600 8842
rect 22756 8430 22784 9438
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22848 7993 22876 14214
rect 22940 13025 22968 15370
rect 22926 13016 22982 13025
rect 23032 12986 23060 15370
rect 23124 15094 23152 15524
rect 23204 15428 23256 15434
rect 23204 15370 23256 15376
rect 23216 15201 23244 15370
rect 23202 15192 23258 15201
rect 23202 15127 23258 15136
rect 23308 15094 23336 17031
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23400 16114 23428 16526
rect 23388 16108 23440 16114
rect 23388 16050 23440 16056
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 23124 13938 23152 15030
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23308 14521 23336 14554
rect 23294 14512 23350 14521
rect 23294 14447 23350 14456
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 14074 23336 14214
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23112 13796 23164 13802
rect 23112 13738 23164 13744
rect 23124 13161 23152 13738
rect 23308 13258 23336 14010
rect 23400 13530 23428 14758
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23492 13274 23520 18090
rect 23584 14822 23612 18255
rect 23676 16590 23704 19638
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 23676 14498 23704 15846
rect 23584 14470 23704 14498
rect 23584 13394 23612 14470
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23676 13462 23704 14350
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23296 13252 23348 13258
rect 23492 13246 23704 13274
rect 23296 13194 23348 13200
rect 23110 13152 23166 13161
rect 23110 13087 23166 13096
rect 22926 12951 22982 12960
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23018 12880 23074 12889
rect 23018 12815 23020 12824
rect 23072 12815 23074 12824
rect 23480 12844 23532 12850
rect 23020 12786 23072 12792
rect 23480 12786 23532 12792
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22940 12356 22968 12718
rect 23018 12472 23074 12481
rect 23492 12442 23520 12786
rect 23480 12436 23532 12442
rect 23074 12416 23428 12434
rect 23018 12407 23428 12416
rect 23032 12406 23428 12407
rect 22940 12328 23152 12356
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 22926 11792 22982 11801
rect 22926 11727 22982 11736
rect 22940 11694 22968 11727
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 23032 10266 23060 12106
rect 23124 11694 23152 12328
rect 23400 12322 23428 12406
rect 23480 12378 23532 12384
rect 23400 12294 23520 12322
rect 23204 12164 23256 12170
rect 23204 12106 23256 12112
rect 23216 12073 23244 12106
rect 23202 12064 23258 12073
rect 23202 11999 23258 12008
rect 23112 11688 23164 11694
rect 23112 11630 23164 11636
rect 23124 11082 23152 11630
rect 23216 11150 23244 11999
rect 23492 11830 23520 12294
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23676 11218 23704 13246
rect 23768 12186 23796 19790
rect 23860 18601 23888 20334
rect 23952 19514 23980 20567
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24044 19446 24072 29446
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 24308 28620 24360 28626
rect 24308 28562 24360 28568
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 24136 21554 24164 25978
rect 24228 25906 24256 28018
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 24320 24664 24348 28562
rect 24952 28484 25004 28490
rect 24952 28426 25004 28432
rect 24964 28014 24992 28426
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 24952 28008 25004 28014
rect 24952 27950 25004 27956
rect 24780 27606 24808 27950
rect 25148 27674 25176 28018
rect 25136 27668 25188 27674
rect 25136 27610 25188 27616
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24412 24886 24440 25638
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 24320 24636 24440 24664
rect 24216 21956 24268 21962
rect 24216 21898 24268 21904
rect 24228 21690 24256 21898
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24136 21049 24164 21490
rect 24122 21040 24178 21049
rect 24122 20975 24178 20984
rect 24122 20496 24178 20505
rect 24122 20431 24124 20440
rect 24176 20431 24178 20440
rect 24124 20402 24176 20408
rect 24228 19854 24256 21490
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24320 20369 24348 20402
rect 24306 20360 24362 20369
rect 24306 20295 24362 20304
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24320 19990 24348 20198
rect 24308 19984 24360 19990
rect 24308 19926 24360 19932
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24032 19440 24084 19446
rect 24084 19400 24164 19428
rect 24032 19382 24084 19388
rect 24032 18624 24084 18630
rect 23846 18592 23902 18601
rect 24032 18566 24084 18572
rect 23846 18527 23902 18536
rect 24044 18358 24072 18566
rect 24032 18352 24084 18358
rect 24032 18294 24084 18300
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 23846 17776 23902 17785
rect 23846 17711 23902 17720
rect 23860 17678 23888 17711
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17338 23980 17478
rect 24044 17338 24072 18158
rect 24136 17882 24164 19400
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24124 17536 24176 17542
rect 24124 17478 24176 17484
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23952 16574 23980 17138
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24044 16794 24072 16934
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 23952 16546 24072 16574
rect 24044 14600 24072 16546
rect 24136 16289 24164 17478
rect 24122 16280 24178 16289
rect 24122 16215 24178 16224
rect 24044 14572 24164 14600
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23860 12306 23888 13262
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23952 12209 23980 13670
rect 24044 12986 24072 14418
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 23938 12200 23994 12209
rect 23768 12158 23888 12186
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23768 11558 23796 12038
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23756 11280 23808 11286
rect 23860 11268 23888 12158
rect 23938 12135 23994 12144
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23952 11830 23980 12038
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 24044 11558 24072 11834
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 23808 11240 23888 11268
rect 24136 11234 24164 14572
rect 23756 11222 23808 11228
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 23480 11076 23532 11082
rect 23480 11018 23532 11024
rect 23492 10810 23520 11018
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23662 10704 23718 10713
rect 23112 10668 23164 10674
rect 23662 10639 23718 10648
rect 23112 10610 23164 10616
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23124 9976 23152 10610
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 22940 9948 23152 9976
rect 22834 7984 22890 7993
rect 22834 7919 22890 7928
rect 22836 7472 22888 7478
rect 22650 7440 22706 7449
rect 22836 7414 22888 7420
rect 22650 7375 22706 7384
rect 22560 6248 22612 6254
rect 22374 6216 22430 6225
rect 22560 6190 22612 6196
rect 22374 6151 22430 6160
rect 22466 5808 22522 5817
rect 22204 5766 22416 5794
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22020 4950 22140 4978
rect 22020 4706 22048 4950
rect 22098 4856 22154 4865
rect 22098 4791 22100 4800
rect 22152 4791 22154 4800
rect 22100 4762 22152 4768
rect 22020 4678 22140 4706
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21730 4040 21786 4049
rect 21730 3975 21786 3984
rect 22006 4040 22062 4049
rect 22006 3975 22062 3984
rect 21916 3664 21968 3670
rect 21652 3624 21916 3652
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21456 3392 21508 3398
rect 21456 3334 21508 3340
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21468 3126 21496 3334
rect 21560 3194 21588 3334
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21456 3120 21508 3126
rect 21456 3062 21508 3068
rect 21836 2825 21864 3624
rect 21916 3606 21968 3612
rect 22020 3534 22048 3975
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 21822 2816 21878 2825
rect 21284 2746 21588 2774
rect 21822 2751 21878 2760
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 21560 2446 21588 2746
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20720 1352 20772 1358
rect 20720 1294 20772 1300
rect 21284 800 21312 2314
rect 21928 800 21956 2994
rect 22112 1766 22140 4678
rect 22204 3602 22232 5646
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22296 5030 22324 5170
rect 22284 5024 22336 5030
rect 22282 4992 22284 5001
rect 22336 4992 22338 5001
rect 22282 4927 22338 4936
rect 22388 4758 22416 5766
rect 22466 5743 22522 5752
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22480 4146 22508 5743
rect 22664 5710 22692 7375
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22756 7002 22784 7142
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22296 3398 22324 3470
rect 22284 3392 22336 3398
rect 22284 3334 22336 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 22204 2514 22232 2858
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22296 2009 22324 3334
rect 22282 2000 22338 2009
rect 22282 1935 22338 1944
rect 22664 1902 22692 3334
rect 22652 1896 22704 1902
rect 22652 1838 22704 1844
rect 22756 1834 22784 6598
rect 22848 3194 22876 7414
rect 22940 6361 22968 9948
rect 23216 9450 23244 10134
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23204 9444 23256 9450
rect 23204 9386 23256 9392
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 22926 6352 22982 6361
rect 22926 6287 22982 6296
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22940 5234 22968 6054
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23032 4010 23060 8502
rect 23112 8356 23164 8362
rect 23112 8298 23164 8304
rect 23124 7546 23152 8298
rect 23216 7886 23244 8910
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23124 5846 23152 6054
rect 23112 5840 23164 5846
rect 23112 5782 23164 5788
rect 23110 5128 23166 5137
rect 23110 5063 23166 5072
rect 23124 4214 23152 5063
rect 23112 4208 23164 4214
rect 23112 4150 23164 4156
rect 23020 4004 23072 4010
rect 23020 3946 23072 3952
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23216 2922 23244 7346
rect 23308 6662 23336 9862
rect 23386 8664 23442 8673
rect 23386 8599 23442 8608
rect 23570 8664 23626 8673
rect 23570 8599 23626 8608
rect 23400 8430 23428 8599
rect 23584 8566 23612 8599
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23676 8498 23704 10639
rect 23768 10305 23796 11222
rect 24044 11206 24164 11234
rect 23938 11112 23994 11121
rect 23938 11047 23994 11056
rect 23754 10296 23810 10305
rect 23754 10231 23810 10240
rect 23952 10198 23980 11047
rect 24044 10606 24072 11206
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 23940 10192 23992 10198
rect 23940 10134 23992 10140
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 7886 23428 8230
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23386 6896 23442 6905
rect 23386 6831 23388 6840
rect 23440 6831 23442 6840
rect 23388 6802 23440 6808
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23308 3194 23336 4082
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 23204 2916 23256 2922
rect 23204 2858 23256 2864
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 23308 2689 23336 2790
rect 23294 2680 23350 2689
rect 23294 2615 23350 2624
rect 23294 2544 23350 2553
rect 23294 2479 23350 2488
rect 23308 2446 23336 2479
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 22744 1828 22796 1834
rect 22744 1770 22796 1776
rect 22100 1760 22152 1766
rect 22100 1702 22152 1708
rect 23216 800 23244 2246
rect 23400 1329 23428 5510
rect 23492 4690 23520 8366
rect 23572 8288 23624 8294
rect 23768 8265 23796 8774
rect 23848 8492 23900 8498
rect 23848 8434 23900 8440
rect 23572 8230 23624 8236
rect 23754 8256 23810 8265
rect 23584 7818 23612 8230
rect 23754 8191 23810 8200
rect 23572 7812 23624 7818
rect 23572 7754 23624 7760
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23570 6624 23626 6633
rect 23570 6559 23626 6568
rect 23584 6458 23612 6559
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23768 1630 23796 6734
rect 23860 5914 23888 8434
rect 24044 5953 24072 9930
rect 24030 5944 24086 5953
rect 23848 5908 23900 5914
rect 24030 5879 24086 5888
rect 23848 5850 23900 5856
rect 24136 5370 24164 11086
rect 24228 8022 24256 19790
rect 24306 18864 24362 18873
rect 24306 18799 24362 18808
rect 24320 16182 24348 18799
rect 24308 16176 24360 16182
rect 24308 16118 24360 16124
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24320 13870 24348 14894
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24320 7721 24348 12174
rect 24306 7712 24362 7721
rect 24306 7647 24362 7656
rect 24412 6458 24440 24636
rect 24584 24608 24636 24614
rect 24584 24550 24636 24556
rect 24490 24168 24546 24177
rect 24490 24103 24546 24112
rect 24504 23730 24532 24103
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24504 21078 24532 21966
rect 24492 21072 24544 21078
rect 24492 21014 24544 21020
rect 24492 20256 24544 20262
rect 24492 20198 24544 20204
rect 24504 19854 24532 20198
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 24504 18222 24532 19178
rect 24492 18216 24544 18222
rect 24492 18158 24544 18164
rect 24492 17604 24544 17610
rect 24492 17546 24544 17552
rect 24504 15978 24532 17546
rect 24492 15972 24544 15978
rect 24492 15914 24544 15920
rect 24596 15638 24624 24550
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24688 23186 24716 24006
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24780 22556 24808 27542
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24872 22930 24900 27474
rect 25044 25152 25096 25158
rect 25044 25094 25096 25100
rect 25056 24886 25084 25094
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 24952 24132 25004 24138
rect 24952 24074 25004 24080
rect 24964 23866 24992 24074
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24964 23050 24992 23462
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24872 22902 24992 22930
rect 24860 22568 24912 22574
rect 24688 22528 24860 22556
rect 24688 19310 24716 22528
rect 24860 22510 24912 22516
rect 24964 22409 24992 22902
rect 24950 22400 25006 22409
rect 24950 22335 25006 22344
rect 24858 22264 24914 22273
rect 24858 22199 24914 22208
rect 24872 21690 24900 22199
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24676 18692 24728 18698
rect 24780 18680 24808 20742
rect 24872 19786 24900 20810
rect 24950 20768 25006 20777
rect 24950 20703 25006 20712
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24964 18902 24992 20703
rect 25056 19854 25084 23666
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 25056 19417 25084 19790
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 25148 19310 25176 27610
rect 25240 26897 25268 29174
rect 25332 28626 25360 30534
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 26068 29102 26096 29582
rect 26056 29096 26108 29102
rect 26056 29038 26108 29044
rect 25320 28620 25372 28626
rect 25320 28562 25372 28568
rect 25504 28620 25556 28626
rect 25504 28562 25556 28568
rect 25412 28484 25464 28490
rect 25412 28426 25464 28432
rect 25424 28218 25452 28426
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 25516 27538 25544 28562
rect 26148 28484 26200 28490
rect 26148 28426 26200 28432
rect 25964 28416 26016 28422
rect 25964 28358 26016 28364
rect 25976 28218 26004 28358
rect 25964 28212 26016 28218
rect 25964 28154 26016 28160
rect 25504 27532 25556 27538
rect 25504 27474 25556 27480
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25884 27130 25912 27338
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25226 26888 25282 26897
rect 25226 26823 25282 26832
rect 25792 26450 25820 26930
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25780 26444 25832 26450
rect 25780 26386 25832 26392
rect 25596 26240 25648 26246
rect 25596 26182 25648 26188
rect 25608 25974 25636 26182
rect 25596 25968 25648 25974
rect 25596 25910 25648 25916
rect 25884 24342 25912 26726
rect 25872 24336 25924 24342
rect 25872 24278 25924 24284
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 24952 18896 25004 18902
rect 24952 18838 25004 18844
rect 25136 18692 25188 18698
rect 24780 18652 25136 18680
rect 24676 18634 24728 18640
rect 25136 18634 25188 18640
rect 24688 18601 24716 18634
rect 24674 18592 24730 18601
rect 24674 18527 24730 18536
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24872 17882 24900 18294
rect 25044 18148 25096 18154
rect 25044 18090 25096 18096
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24688 17610 24716 17818
rect 24676 17604 24728 17610
rect 24676 17546 24728 17552
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24688 16046 24716 16458
rect 24780 16182 24808 17546
rect 24950 17504 25006 17513
rect 24950 17439 25006 17448
rect 24858 17368 24914 17377
rect 24858 17303 24914 17312
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24872 16114 24900 17303
rect 24964 17270 24992 17439
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 24964 17105 24992 17206
rect 24950 17096 25006 17105
rect 24950 17031 25006 17040
rect 25056 16833 25084 18090
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25148 17134 25176 17274
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25042 16824 25098 16833
rect 25042 16759 25098 16768
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24872 15745 24900 16050
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24858 15736 24914 15745
rect 24858 15671 24914 15680
rect 24584 15632 24636 15638
rect 24584 15574 24636 15580
rect 24964 15094 24992 15846
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 9636 24532 14758
rect 24596 14278 24624 14894
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24584 14272 24636 14278
rect 24584 14214 24636 14220
rect 24596 14090 24624 14214
rect 24596 14062 24808 14090
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24596 12986 24624 13874
rect 24674 13288 24730 13297
rect 24674 13223 24676 13232
rect 24728 13223 24730 13232
rect 24676 13194 24728 13200
rect 24584 12980 24636 12986
rect 24780 12968 24808 14062
rect 24872 13802 24900 14282
rect 25056 14249 25084 16050
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 25148 15434 25176 15846
rect 25136 15428 25188 15434
rect 25136 15370 25188 15376
rect 25042 14240 25098 14249
rect 25042 14175 25098 14184
rect 24860 13796 24912 13802
rect 24860 13738 24912 13744
rect 24780 12940 24992 12968
rect 24584 12922 24636 12928
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24596 11937 24624 12174
rect 24582 11928 24638 11937
rect 24582 11863 24638 11872
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24596 11529 24624 11630
rect 24582 11520 24638 11529
rect 24582 11455 24638 11464
rect 24688 11234 24716 12174
rect 24596 11206 24716 11234
rect 24596 11150 24624 11206
rect 24780 11150 24808 12786
rect 24872 11354 24900 12786
rect 24964 12306 24992 12940
rect 25240 12850 25268 23802
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25332 20874 25360 21286
rect 25516 21146 25544 22986
rect 25976 22710 26004 28154
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 26068 25158 26096 27270
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 26068 24818 26096 25094
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 25964 22704 26016 22710
rect 25964 22646 26016 22652
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25976 21078 26004 22646
rect 25780 21072 25832 21078
rect 25780 21014 25832 21020
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25596 19984 25648 19990
rect 25596 19926 25648 19932
rect 25410 19680 25466 19689
rect 25410 19615 25466 19624
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25332 18426 25360 19246
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25424 17785 25452 19615
rect 25608 19446 25636 19926
rect 25700 19922 25728 20334
rect 25792 20330 25820 21014
rect 25962 20904 26018 20913
rect 25962 20839 25964 20848
rect 26016 20839 26018 20848
rect 25964 20810 26016 20816
rect 26160 20618 26188 28426
rect 26240 25764 26292 25770
rect 26240 25706 26292 25712
rect 26252 25362 26280 25706
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26252 22710 26280 23462
rect 26240 22704 26292 22710
rect 26240 22646 26292 22652
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26068 20590 26188 20618
rect 25964 20392 26016 20398
rect 25962 20360 25964 20369
rect 26016 20360 26018 20369
rect 25780 20324 25832 20330
rect 25962 20295 26018 20304
rect 25780 20266 25832 20272
rect 26068 20210 26096 20590
rect 26148 20528 26200 20534
rect 26148 20470 26200 20476
rect 25976 20182 26096 20210
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25608 19310 25636 19382
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 25504 18828 25556 18834
rect 25688 18828 25740 18834
rect 25556 18788 25636 18816
rect 25504 18770 25556 18776
rect 25410 17776 25466 17785
rect 25410 17711 25466 17720
rect 25412 17604 25464 17610
rect 25412 17546 25464 17552
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 25332 14793 25360 14962
rect 25318 14784 25374 14793
rect 25318 14719 25374 14728
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 25134 12200 25190 12209
rect 25134 12135 25136 12144
rect 25188 12135 25190 12144
rect 25136 12106 25188 12112
rect 25134 11792 25190 11801
rect 25134 11727 25190 11736
rect 25148 11694 25176 11727
rect 25136 11688 25188 11694
rect 25136 11630 25188 11636
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24584 11008 24636 11014
rect 24584 10950 24636 10956
rect 24596 10033 24624 10950
rect 24582 10024 24638 10033
rect 24582 9959 24638 9968
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24504 9608 24624 9636
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24504 7546 24532 9454
rect 24596 9450 24624 9608
rect 24688 9518 24716 9658
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24674 9208 24730 9217
rect 24674 9143 24730 9152
rect 24582 8664 24638 8673
rect 24582 8599 24638 8608
rect 24596 8498 24624 8599
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24688 8362 24716 9143
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24504 7274 24532 7482
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24492 7268 24544 7274
rect 24492 7210 24544 7216
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 24124 4480 24176 4486
rect 24124 4422 24176 4428
rect 24136 4146 24164 4422
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 23940 3936 23992 3942
rect 23938 3904 23940 3913
rect 23992 3904 23994 3913
rect 23938 3839 23994 3848
rect 24596 3738 24624 7278
rect 24688 7177 24716 7890
rect 24674 7168 24730 7177
rect 24674 7103 24730 7112
rect 24674 6896 24730 6905
rect 24674 6831 24676 6840
rect 24728 6831 24730 6840
rect 24676 6802 24728 6808
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24032 3528 24084 3534
rect 24030 3496 24032 3505
rect 24084 3496 24086 3505
rect 24030 3431 24086 3440
rect 23940 3392 23992 3398
rect 23940 3334 23992 3340
rect 23952 3058 23980 3334
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23756 1624 23808 1630
rect 23756 1566 23808 1572
rect 23386 1320 23442 1329
rect 23386 1255 23442 1264
rect 23860 800 23888 2790
rect 24780 2514 24808 11086
rect 24860 11008 24912 11014
rect 24860 10950 24912 10956
rect 24872 8129 24900 10950
rect 25044 10736 25096 10742
rect 25044 10678 25096 10684
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24858 8120 24914 8129
rect 24858 8055 24914 8064
rect 24964 7750 24992 10542
rect 25056 9722 25084 10678
rect 25148 10606 25176 11154
rect 25136 10600 25188 10606
rect 25136 10542 25188 10548
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 25042 9072 25098 9081
rect 25042 9007 25098 9016
rect 25056 8498 25084 9007
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24858 7576 24914 7585
rect 24858 7511 24860 7520
rect 24912 7511 24914 7520
rect 24860 7482 24912 7488
rect 24964 6118 24992 7686
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24858 5536 24914 5545
rect 24858 5471 24914 5480
rect 24872 2582 24900 5471
rect 25042 2952 25098 2961
rect 25042 2887 25098 2896
rect 25056 2854 25084 2887
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25240 2774 25268 12786
rect 25332 11937 25360 14719
rect 25424 14414 25452 17546
rect 25502 15600 25558 15609
rect 25502 15535 25558 15544
rect 25516 15094 25544 15535
rect 25504 15088 25556 15094
rect 25504 15030 25556 15036
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25318 11928 25374 11937
rect 25318 11863 25374 11872
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 25332 10266 25360 11766
rect 25424 11354 25452 13806
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25424 10606 25452 11086
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25516 10062 25544 13126
rect 25608 11393 25636 18788
rect 25688 18770 25740 18776
rect 25700 18737 25728 18770
rect 25686 18728 25742 18737
rect 25686 18663 25742 18672
rect 25700 18290 25728 18663
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25686 16688 25742 16697
rect 25686 16623 25742 16632
rect 25700 14822 25728 16623
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 25700 14278 25728 14418
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 12714 25728 13194
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25700 11830 25728 12650
rect 25688 11824 25740 11830
rect 25688 11766 25740 11772
rect 25594 11384 25650 11393
rect 25594 11319 25650 11328
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25424 9654 25452 9862
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25608 9586 25636 11319
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25700 10169 25728 10610
rect 25686 10160 25742 10169
rect 25686 10095 25742 10104
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25792 9110 25820 19654
rect 25976 18834 26004 20182
rect 26054 20088 26110 20097
rect 26054 20023 26110 20032
rect 26068 19417 26096 20023
rect 26054 19408 26110 19417
rect 26054 19343 26110 19352
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25976 18358 26004 18634
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25884 15978 25912 16390
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 25870 14512 25926 14521
rect 25870 14447 25926 14456
rect 25884 14346 25912 14447
rect 25976 14385 26004 17818
rect 26068 16522 26096 19343
rect 26160 19009 26188 20470
rect 26252 19825 26280 20878
rect 26344 20602 26372 35866
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26528 27538 26556 29446
rect 26896 28762 26924 33934
rect 26988 29646 27016 36722
rect 27540 34202 27568 37198
rect 27724 37194 27752 39200
rect 27712 37188 27764 37194
rect 27712 37130 27764 37136
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 28644 36922 28672 37062
rect 28632 36916 28684 36922
rect 28632 36858 28684 36864
rect 28736 36802 28764 37062
rect 28460 36774 28764 36802
rect 29012 36786 29040 39200
rect 29656 37126 29684 39200
rect 30944 37330 30972 39200
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 29736 37256 29788 37262
rect 29736 37198 29788 37204
rect 31208 37256 31260 37262
rect 31208 37198 31260 37204
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29000 36780 29052 36786
rect 28460 36582 28488 36774
rect 29000 36722 29052 36728
rect 28724 36712 28776 36718
rect 28724 36654 28776 36660
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28540 36576 28592 36582
rect 28540 36518 28592 36524
rect 28080 35216 28132 35222
rect 28080 35158 28132 35164
rect 27804 34604 27856 34610
rect 27804 34546 27856 34552
rect 27528 34196 27580 34202
rect 27528 34138 27580 34144
rect 27160 32496 27212 32502
rect 27160 32438 27212 32444
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26884 28756 26936 28762
rect 26884 28698 26936 28704
rect 26516 27532 26568 27538
rect 26516 27474 26568 27480
rect 26424 26580 26476 26586
rect 26424 26522 26476 26528
rect 26436 23225 26464 26522
rect 26528 23662 26556 27474
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26620 23730 26648 24754
rect 26608 23724 26660 23730
rect 26608 23666 26660 23672
rect 26516 23656 26568 23662
rect 26516 23598 26568 23604
rect 26422 23216 26478 23225
rect 26422 23151 26478 23160
rect 26620 22658 26648 23666
rect 26712 22778 26740 25162
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 26976 24744 27028 24750
rect 26976 24686 27028 24692
rect 26700 22772 26752 22778
rect 26700 22714 26752 22720
rect 26620 22630 26740 22658
rect 26516 22500 26568 22506
rect 26516 22442 26568 22448
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26436 21554 26464 22102
rect 26528 22098 26556 22442
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26436 19922 26464 21490
rect 26424 19916 26476 19922
rect 26424 19858 26476 19864
rect 26238 19816 26294 19825
rect 26238 19751 26294 19760
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 26436 19446 26464 19654
rect 26424 19440 26476 19446
rect 26424 19382 26476 19388
rect 26146 19000 26202 19009
rect 26146 18935 26202 18944
rect 26424 18964 26476 18970
rect 26160 18766 26188 18935
rect 26424 18906 26476 18912
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26332 18624 26384 18630
rect 26330 18592 26332 18601
rect 26384 18592 26386 18601
rect 26330 18527 26386 18536
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26252 16522 26280 17070
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 26160 15706 26188 16050
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26344 15502 26372 18158
rect 26436 15706 26464 18906
rect 26516 18148 26568 18154
rect 26516 18090 26568 18096
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 26252 15178 26280 15370
rect 26160 15150 26280 15178
rect 26160 14958 26188 15150
rect 26240 15020 26292 15026
rect 26240 14962 26292 14968
rect 26148 14952 26200 14958
rect 26054 14920 26110 14929
rect 26148 14894 26200 14900
rect 26054 14855 26110 14864
rect 25962 14376 26018 14385
rect 25872 14340 25924 14346
rect 25962 14311 26018 14320
rect 25872 14282 25924 14288
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25884 11014 25912 13806
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25872 10532 25924 10538
rect 25872 10474 25924 10480
rect 25884 10062 25912 10474
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25780 9104 25832 9110
rect 25780 9046 25832 9052
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25502 8528 25558 8537
rect 25502 8463 25504 8472
rect 25556 8463 25558 8472
rect 25504 8434 25556 8440
rect 25608 7818 25636 8774
rect 25700 8401 25728 8774
rect 25686 8392 25742 8401
rect 25686 8327 25742 8336
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25976 7478 26004 12718
rect 26068 12434 26096 14855
rect 26252 12714 26280 14962
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26148 12640 26200 12646
rect 26200 12588 26280 12594
rect 26148 12582 26280 12588
rect 26160 12566 26280 12582
rect 26148 12436 26200 12442
rect 26068 12406 26148 12434
rect 26148 12378 26200 12384
rect 26056 12300 26108 12306
rect 26056 12242 26108 12248
rect 26068 12073 26096 12242
rect 26054 12064 26110 12073
rect 26054 11999 26110 12008
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 25964 7472 26016 7478
rect 25964 7414 26016 7420
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25884 3194 25912 6734
rect 26068 3369 26096 11086
rect 26146 10840 26202 10849
rect 26146 10775 26148 10784
rect 26200 10775 26202 10784
rect 26148 10746 26200 10752
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 26160 9518 26188 10542
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 26160 8809 26188 9454
rect 26146 8800 26202 8809
rect 26146 8735 26202 8744
rect 26252 8090 26280 12566
rect 26344 11694 26372 15438
rect 26424 15360 26476 15366
rect 26424 15302 26476 15308
rect 26436 14618 26464 15302
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26528 14346 26556 18090
rect 26620 15434 26648 22374
rect 26712 18442 26740 22630
rect 26988 22098 27016 24686
rect 27080 23089 27108 25094
rect 27066 23080 27122 23089
rect 27066 23015 27122 23024
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 27080 22166 27108 22578
rect 27068 22160 27120 22166
rect 27068 22102 27120 22108
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26884 22024 26936 22030
rect 26882 21992 26884 22001
rect 26936 21992 26938 22001
rect 26882 21927 26938 21936
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27080 20262 27108 20402
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 27080 19553 27108 19654
rect 27066 19544 27122 19553
rect 27066 19479 27122 19488
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 26790 19272 26846 19281
rect 26790 19207 26846 19216
rect 26884 19236 26936 19242
rect 26804 19174 26832 19207
rect 26884 19178 26936 19184
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26804 18766 26832 19110
rect 26896 18970 26924 19178
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26712 18414 26924 18442
rect 26700 18284 26752 18290
rect 26700 18226 26752 18232
rect 26608 15428 26660 15434
rect 26608 15370 26660 15376
rect 26620 15162 26648 15370
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26620 14657 26648 14894
rect 26606 14648 26662 14657
rect 26606 14583 26662 14592
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26608 14340 26660 14346
rect 26608 14282 26660 14288
rect 26422 14240 26478 14249
rect 26422 14175 26478 14184
rect 26436 13938 26464 14175
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26528 13462 26556 14282
rect 26620 14249 26648 14282
rect 26606 14240 26662 14249
rect 26606 14175 26662 14184
rect 26606 14104 26662 14113
rect 26606 14039 26608 14048
rect 26660 14039 26662 14048
rect 26608 14010 26660 14016
rect 26606 13560 26662 13569
rect 26606 13495 26662 13504
rect 26516 13456 26568 13462
rect 26516 13398 26568 13404
rect 26514 12744 26570 12753
rect 26514 12679 26570 12688
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26436 8022 26464 12106
rect 26528 11150 26556 12679
rect 26620 11354 26648 13495
rect 26712 11762 26740 18226
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26712 10674 26740 11698
rect 26804 10985 26832 17614
rect 26896 16153 26924 18414
rect 26882 16144 26938 16153
rect 26882 16079 26938 16088
rect 26988 16017 27016 19382
rect 27068 19236 27120 19242
rect 27068 19178 27120 19184
rect 27080 19145 27108 19178
rect 27066 19136 27122 19145
rect 27066 19071 27122 19080
rect 27068 18964 27120 18970
rect 27068 18906 27120 18912
rect 27080 18329 27108 18906
rect 27066 18320 27122 18329
rect 27066 18255 27122 18264
rect 27172 17954 27200 32438
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27448 29034 27476 30194
rect 27816 29850 27844 34546
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27448 28558 27476 28970
rect 27436 28552 27488 28558
rect 27436 28494 27488 28500
rect 27804 28076 27856 28082
rect 27804 28018 27856 28024
rect 27436 28008 27488 28014
rect 27436 27950 27488 27956
rect 27252 27396 27304 27402
rect 27252 27338 27304 27344
rect 27264 27130 27292 27338
rect 27252 27124 27304 27130
rect 27252 27066 27304 27072
rect 27252 26240 27304 26246
rect 27252 26182 27304 26188
rect 27264 25838 27292 26182
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 27252 25832 27304 25838
rect 27252 25774 27304 25780
rect 27264 25362 27292 25774
rect 27252 25356 27304 25362
rect 27252 25298 27304 25304
rect 27356 24954 27384 25910
rect 27344 24948 27396 24954
rect 27344 24890 27396 24896
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27356 23798 27384 24006
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 27264 21010 27292 23598
rect 27448 21486 27476 27950
rect 27816 27418 27844 28018
rect 27896 27464 27948 27470
rect 27816 27412 27896 27418
rect 27816 27406 27948 27412
rect 27816 27390 27936 27406
rect 27712 26920 27764 26926
rect 27712 26862 27764 26868
rect 27620 26580 27672 26586
rect 27620 26522 27672 26528
rect 27632 25498 27660 26522
rect 27724 26450 27752 26862
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 27528 25492 27580 25498
rect 27528 25434 27580 25440
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 27436 21480 27488 21486
rect 27436 21422 27488 21428
rect 27540 21332 27568 25434
rect 27816 22137 27844 27390
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27908 23186 27936 23598
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 27802 22128 27858 22137
rect 27802 22063 27858 22072
rect 27448 21304 27568 21332
rect 27252 21004 27304 21010
rect 27252 20946 27304 20952
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27264 18442 27292 19790
rect 27356 19446 27384 20198
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 27342 18456 27398 18465
rect 27264 18414 27342 18442
rect 27342 18391 27398 18400
rect 27250 18184 27306 18193
rect 27250 18119 27252 18128
rect 27304 18119 27306 18128
rect 27252 18090 27304 18096
rect 27080 17926 27200 17954
rect 27080 17678 27108 17926
rect 27250 17912 27306 17921
rect 27250 17847 27306 17856
rect 27264 17746 27292 17847
rect 27252 17740 27304 17746
rect 27252 17682 27304 17688
rect 27068 17672 27120 17678
rect 27068 17614 27120 17620
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 27264 17134 27292 17546
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27066 16824 27122 16833
rect 27066 16759 27122 16768
rect 27252 16788 27304 16794
rect 27080 16522 27108 16759
rect 27252 16730 27304 16736
rect 27068 16516 27120 16522
rect 27068 16458 27120 16464
rect 26974 16008 27030 16017
rect 26974 15943 27030 15952
rect 26988 15638 27016 15943
rect 26976 15632 27028 15638
rect 26976 15574 27028 15580
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26790 10976 26846 10985
rect 26790 10911 26846 10920
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26896 10577 26924 14758
rect 26988 12170 27016 15438
rect 27080 15008 27108 16458
rect 27264 16250 27292 16730
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27356 16130 27384 18391
rect 27448 17542 27476 21304
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27816 20534 27844 20878
rect 27804 20528 27856 20534
rect 27896 20528 27948 20534
rect 27804 20470 27856 20476
rect 27894 20496 27896 20505
rect 27948 20496 27950 20505
rect 27894 20431 27950 20440
rect 27712 19984 27764 19990
rect 27710 19952 27712 19961
rect 27764 19952 27766 19961
rect 27710 19887 27766 19896
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27620 19440 27672 19446
rect 27618 19408 27620 19417
rect 27672 19408 27674 19417
rect 27618 19343 27674 19352
rect 27816 18698 27844 19654
rect 27804 18692 27856 18698
rect 27804 18634 27856 18640
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27436 17536 27488 17542
rect 27436 17478 27488 17484
rect 27540 17338 27568 18294
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27436 17332 27488 17338
rect 27436 17274 27488 17280
rect 27528 17332 27580 17338
rect 27528 17274 27580 17280
rect 27448 16794 27476 17274
rect 27528 17128 27580 17134
rect 27526 17096 27528 17105
rect 27580 17096 27582 17105
rect 27526 17031 27582 17040
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27632 16590 27660 18022
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27710 17232 27766 17241
rect 27710 17167 27766 17176
rect 27724 17134 27752 17167
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27724 16590 27752 17070
rect 27908 16776 27936 17682
rect 28000 17490 28028 22986
rect 28092 22778 28120 35158
rect 28552 32434 28580 36518
rect 28736 36242 28764 36654
rect 28724 36236 28776 36242
rect 28724 36178 28776 36184
rect 29748 34746 29776 37198
rect 31220 36378 31248 37198
rect 31588 37108 31616 39200
rect 32232 37466 32260 39200
rect 32220 37460 32272 37466
rect 32220 37402 32272 37408
rect 33048 37256 33100 37262
rect 33048 37198 33100 37204
rect 31760 37120 31812 37126
rect 31588 37080 31760 37108
rect 31760 37062 31812 37068
rect 33060 36718 33088 37198
rect 33520 37126 33548 39200
rect 34164 37330 34192 39200
rect 35452 39114 35480 39200
rect 35544 39114 35572 39222
rect 35452 39086 35572 39114
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34152 37324 34204 37330
rect 34152 37266 34204 37272
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33048 36712 33100 36718
rect 33048 36654 33100 36660
rect 31208 36372 31260 36378
rect 31208 36314 31260 36320
rect 33796 36174 33824 37198
rect 35820 37108 35848 39222
rect 36082 39200 36138 39800
rect 36726 39200 36782 39800
rect 38014 39200 38070 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 36096 37346 36124 39200
rect 36096 37318 36216 37346
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 35900 37120 35952 37126
rect 35820 37080 35900 37108
rect 35900 37062 35952 37068
rect 35900 36780 35952 36786
rect 35900 36722 35952 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 33784 36168 33836 36174
rect 33784 36110 33836 36116
rect 29920 36100 29972 36106
rect 29920 36042 29972 36048
rect 29736 34740 29788 34746
rect 29736 34682 29788 34688
rect 29000 34604 29052 34610
rect 29000 34546 29052 34552
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 28540 32224 28592 32230
rect 28540 32166 28592 32172
rect 28264 24880 28316 24886
rect 28264 24822 28316 24828
rect 28276 24410 28304 24822
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 28184 22094 28212 24142
rect 28552 23254 28580 32166
rect 28816 27056 28868 27062
rect 28816 26998 28868 27004
rect 28828 26586 28856 26998
rect 28908 26852 28960 26858
rect 28908 26794 28960 26800
rect 28816 26580 28868 26586
rect 28816 26522 28868 26528
rect 28724 26376 28776 26382
rect 28724 26318 28776 26324
rect 28736 26042 28764 26318
rect 28724 26036 28776 26042
rect 28724 25978 28776 25984
rect 28920 25974 28948 26794
rect 29012 26790 29040 34546
rect 29000 26784 29052 26790
rect 29000 26726 29052 26732
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 28908 25968 28960 25974
rect 28908 25910 28960 25916
rect 28632 25424 28684 25430
rect 28632 25366 28684 25372
rect 28644 23798 28672 25366
rect 28920 24886 28948 25910
rect 29460 25492 29512 25498
rect 29460 25434 29512 25440
rect 29092 25288 29144 25294
rect 29092 25230 29144 25236
rect 28908 24880 28960 24886
rect 28908 24822 28960 24828
rect 28920 24274 28948 24822
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28632 23792 28684 23798
rect 28632 23734 28684 23740
rect 28920 23662 28948 24210
rect 28908 23656 28960 23662
rect 28908 23598 28960 23604
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28632 23180 28684 23186
rect 28632 23122 28684 23128
rect 28356 23044 28408 23050
rect 28356 22986 28408 22992
rect 28368 22710 28396 22986
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28092 22066 28212 22094
rect 28092 19242 28120 22066
rect 28368 21486 28396 22646
rect 28644 22098 28672 23122
rect 29000 22636 29052 22642
rect 29000 22578 29052 22584
rect 28632 22092 28684 22098
rect 28632 22034 28684 22040
rect 29012 21622 29040 22578
rect 29104 22001 29132 25230
rect 29276 24132 29328 24138
rect 29276 24074 29328 24080
rect 29288 22574 29316 24074
rect 29368 22704 29420 22710
rect 29368 22646 29420 22652
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 29196 22438 29224 22469
rect 29184 22432 29236 22438
rect 29182 22400 29184 22409
rect 29236 22400 29238 22409
rect 29182 22335 29238 22344
rect 29090 21992 29146 22001
rect 29090 21927 29146 21936
rect 28908 21616 28960 21622
rect 28908 21558 28960 21564
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 28816 21344 28868 21350
rect 28630 21312 28686 21321
rect 28816 21286 28868 21292
rect 28630 21247 28686 21256
rect 28644 21010 28672 21247
rect 28828 21146 28856 21286
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28632 21004 28684 21010
rect 28632 20946 28684 20952
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28080 19236 28132 19242
rect 28080 19178 28132 19184
rect 28092 18086 28120 19178
rect 28276 19174 28304 19790
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 28000 17462 28212 17490
rect 27908 16748 28028 16776
rect 27896 16652 27948 16658
rect 27896 16594 27948 16600
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27816 16182 27844 16390
rect 27804 16176 27856 16182
rect 27264 16114 27384 16130
rect 27252 16108 27384 16114
rect 27304 16102 27384 16108
rect 27434 16144 27490 16153
rect 27804 16118 27856 16124
rect 27434 16079 27490 16088
rect 27252 16050 27304 16056
rect 27158 15872 27214 15881
rect 27158 15807 27214 15816
rect 27172 15706 27200 15807
rect 27160 15700 27212 15706
rect 27160 15642 27212 15648
rect 27080 14980 27200 15008
rect 27068 14816 27120 14822
rect 27066 14784 27068 14793
rect 27120 14784 27122 14793
rect 27066 14719 27122 14728
rect 27172 14634 27200 14980
rect 27080 14606 27200 14634
rect 27080 13870 27108 14606
rect 27160 14408 27212 14414
rect 27158 14376 27160 14385
rect 27212 14376 27214 14385
rect 27158 14311 27214 14320
rect 27264 14260 27292 16050
rect 27342 15056 27398 15065
rect 27342 14991 27344 15000
rect 27396 14991 27398 15000
rect 27344 14962 27396 14968
rect 27344 14884 27396 14890
rect 27344 14826 27396 14832
rect 27172 14232 27292 14260
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 27068 13252 27120 13258
rect 27068 13194 27120 13200
rect 27080 12646 27108 13194
rect 27068 12640 27120 12646
rect 27068 12582 27120 12588
rect 27172 12434 27200 14232
rect 27250 13832 27306 13841
rect 27250 13767 27306 13776
rect 27264 13734 27292 13767
rect 27252 13728 27304 13734
rect 27252 13670 27304 13676
rect 27356 12753 27384 14826
rect 27448 14396 27476 16079
rect 27620 15700 27672 15706
rect 27620 15642 27672 15648
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27540 15162 27568 15506
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27632 14550 27660 15642
rect 27804 15632 27856 15638
rect 27804 15574 27856 15580
rect 27712 14952 27764 14958
rect 27712 14894 27764 14900
rect 27724 14618 27752 14894
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27620 14544 27672 14550
rect 27620 14486 27672 14492
rect 27620 14408 27672 14414
rect 27448 14368 27568 14396
rect 27540 12850 27568 14368
rect 27620 14350 27672 14356
rect 27632 13841 27660 14350
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27724 13938 27752 14214
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27618 13832 27674 13841
rect 27618 13767 27674 13776
rect 27724 13682 27752 13874
rect 27632 13654 27752 13682
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 27342 12744 27398 12753
rect 27342 12679 27398 12688
rect 27172 12406 27292 12434
rect 26976 12164 27028 12170
rect 26976 12106 27028 12112
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27068 11824 27120 11830
rect 27068 11766 27120 11772
rect 26976 11620 27028 11626
rect 26976 11562 27028 11568
rect 26882 10568 26938 10577
rect 26882 10503 26938 10512
rect 26988 9042 27016 11562
rect 27080 11354 27108 11766
rect 27172 11626 27200 12038
rect 27264 11762 27292 12406
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27160 11620 27212 11626
rect 27160 11562 27212 11568
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27172 10538 27200 11086
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 27264 8906 27292 10066
rect 27356 9897 27384 12174
rect 27342 9888 27398 9897
rect 27342 9823 27398 9832
rect 27344 9376 27396 9382
rect 27344 9318 27396 9324
rect 27356 8906 27384 9318
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27344 8900 27396 8906
rect 27344 8842 27396 8848
rect 26424 8016 26476 8022
rect 26424 7958 26476 7964
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 26054 3360 26110 3369
rect 26054 3295 26110 3304
rect 25872 3188 25924 3194
rect 25872 3130 25924 3136
rect 25410 3088 25466 3097
rect 25410 3023 25412 3032
rect 25464 3023 25466 3032
rect 25412 2994 25464 3000
rect 25148 2746 25268 2774
rect 25148 2582 25176 2746
rect 26160 2650 26188 7822
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26620 3058 26648 7346
rect 27264 6866 27292 8842
rect 27632 8838 27660 13654
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27724 11218 27752 12038
rect 27712 11212 27764 11218
rect 27712 11154 27764 11160
rect 27816 10198 27844 15574
rect 27908 14278 27936 16594
rect 28000 15450 28028 16748
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 28092 15978 28120 16390
rect 28080 15972 28132 15978
rect 28080 15914 28132 15920
rect 28000 15422 28120 15450
rect 28184 15434 28212 17462
rect 28460 17116 28488 20334
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28552 17270 28580 19654
rect 28828 19446 28856 21082
rect 28920 20602 28948 21558
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28816 19440 28868 19446
rect 28868 19388 28948 19394
rect 28816 19382 28948 19388
rect 28828 19366 28948 19382
rect 28632 18760 28684 18766
rect 28632 18702 28684 18708
rect 28540 17264 28592 17270
rect 28540 17206 28592 17212
rect 28460 17088 28580 17116
rect 28446 16960 28502 16969
rect 28446 16895 28502 16904
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28264 16176 28316 16182
rect 28264 16118 28316 16124
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 27896 14272 27948 14278
rect 27896 14214 27948 14220
rect 28000 13433 28028 15302
rect 27986 13424 28042 13433
rect 27986 13359 28042 13368
rect 27988 12912 28040 12918
rect 27988 12854 28040 12860
rect 28000 12374 28028 12854
rect 28092 12782 28120 15422
rect 28172 15428 28224 15434
rect 28172 15370 28224 15376
rect 28170 14376 28226 14385
rect 28170 14311 28172 14320
rect 28224 14311 28226 14320
rect 28172 14282 28224 14288
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 27988 12368 28040 12374
rect 27988 12310 28040 12316
rect 27896 11008 27948 11014
rect 27896 10950 27948 10956
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 27908 9994 27936 10950
rect 28184 10742 28212 13262
rect 28276 12209 28304 16118
rect 28368 15570 28396 16730
rect 28460 16590 28488 16895
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28368 15094 28396 15506
rect 28460 15434 28488 15846
rect 28448 15428 28500 15434
rect 28448 15370 28500 15376
rect 28356 15088 28408 15094
rect 28356 15030 28408 15036
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 28356 14272 28408 14278
rect 28356 14214 28408 14220
rect 28262 12200 28318 12209
rect 28262 12135 28318 12144
rect 28368 11082 28396 14214
rect 28460 13326 28488 14350
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28552 11626 28580 17088
rect 28644 16425 28672 18702
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28736 17649 28764 18566
rect 28828 18057 28856 18566
rect 28814 18048 28870 18057
rect 28814 17983 28870 17992
rect 28722 17640 28778 17649
rect 28722 17575 28778 17584
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 16726 28856 17478
rect 28920 17066 28948 19366
rect 29012 18714 29040 20402
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29104 18834 29132 19654
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 29012 18686 29132 18714
rect 29000 18216 29052 18222
rect 29000 18158 29052 18164
rect 29012 17134 29040 18158
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 28908 17060 28960 17066
rect 28908 17002 28960 17008
rect 29104 16946 29132 18686
rect 29196 18193 29224 22335
rect 29276 21412 29328 21418
rect 29276 21354 29328 21360
rect 29288 20806 29316 21354
rect 29380 21146 29408 22646
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29276 20800 29328 20806
rect 29276 20742 29328 20748
rect 29472 20534 29500 25434
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29748 23118 29776 23530
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29552 22568 29604 22574
rect 29552 22510 29604 22516
rect 29564 22438 29592 22510
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 29644 21004 29696 21010
rect 29644 20946 29696 20952
rect 29552 20800 29604 20806
rect 29552 20742 29604 20748
rect 29460 20528 29512 20534
rect 29460 20470 29512 20476
rect 29472 19310 29500 20470
rect 29460 19304 29512 19310
rect 29460 19246 29512 19252
rect 29368 18692 29420 18698
rect 29368 18634 29420 18640
rect 29182 18184 29238 18193
rect 29182 18119 29238 18128
rect 29184 18080 29236 18086
rect 29236 18057 29316 18068
rect 29236 18048 29330 18057
rect 29236 18040 29274 18048
rect 29184 18022 29236 18028
rect 29274 17983 29330 17992
rect 29182 17912 29238 17921
rect 29182 17847 29238 17856
rect 29012 16918 29132 16946
rect 28816 16720 28868 16726
rect 28816 16662 28868 16668
rect 28630 16416 28686 16425
rect 29012 16402 29040 16918
rect 29092 16584 29144 16590
rect 29090 16552 29092 16561
rect 29144 16552 29146 16561
rect 29090 16487 29146 16496
rect 29012 16374 29132 16402
rect 28630 16351 28686 16360
rect 28644 13326 28672 16351
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 28816 15428 28868 15434
rect 28816 15370 28868 15376
rect 28724 15088 28776 15094
rect 28724 15030 28776 15036
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28356 11076 28408 11082
rect 28356 11018 28408 11024
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 28736 9654 28764 15030
rect 28828 14521 28856 15370
rect 28814 14512 28870 14521
rect 28814 14447 28870 14456
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28920 14074 28948 14214
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28920 12617 28948 13126
rect 28906 12608 28962 12617
rect 28906 12543 28962 12552
rect 28724 9648 28776 9654
rect 28724 9590 28776 9596
rect 28816 9580 28868 9586
rect 28816 9522 28868 9528
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 28828 3126 28856 9522
rect 29012 8634 29040 15982
rect 29104 15978 29132 16374
rect 29196 16182 29224 17847
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29092 15972 29144 15978
rect 29092 15914 29144 15920
rect 29184 15972 29236 15978
rect 29184 15914 29236 15920
rect 29090 15192 29146 15201
rect 29090 15127 29146 15136
rect 29104 13977 29132 15127
rect 29196 14958 29224 15914
rect 29276 15496 29328 15502
rect 29276 15438 29328 15444
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 29090 13968 29146 13977
rect 29090 13903 29146 13912
rect 29196 12986 29224 14894
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 29288 11257 29316 15438
rect 29380 13870 29408 18634
rect 29458 18184 29514 18193
rect 29458 18119 29460 18128
rect 29512 18119 29514 18128
rect 29460 18090 29512 18096
rect 29564 16182 29592 20742
rect 29656 16726 29684 20946
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29748 20466 29776 20878
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29748 18358 29776 20198
rect 29840 19446 29868 26726
rect 29932 25498 29960 36042
rect 35532 35624 35584 35630
rect 35532 35566 35584 35572
rect 34520 35488 34572 35494
rect 34520 35430 34572 35436
rect 34532 33522 34560 35430
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34520 33516 34572 33522
rect 34520 33458 34572 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 32404 28688 32456 28694
rect 32404 28630 32456 28636
rect 32036 28416 32088 28422
rect 32036 28358 32088 28364
rect 30748 27940 30800 27946
rect 30748 27882 30800 27888
rect 30760 27130 30788 27882
rect 30748 27124 30800 27130
rect 30748 27066 30800 27072
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30852 26314 30880 27066
rect 32048 26926 32076 28358
rect 32036 26920 32088 26926
rect 32036 26862 32088 26868
rect 30840 26308 30892 26314
rect 30840 26250 30892 26256
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 29920 25492 29972 25498
rect 29920 25434 29972 25440
rect 30564 24064 30616 24070
rect 30564 24006 30616 24012
rect 30576 23798 30604 24006
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30564 23316 30616 23322
rect 30564 23258 30616 23264
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 30024 19786 30052 20266
rect 29920 19780 29972 19786
rect 29920 19722 29972 19728
rect 30012 19780 30064 19786
rect 30012 19722 30064 19728
rect 29932 19514 29960 19722
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29828 19440 29880 19446
rect 29828 19382 29880 19388
rect 29736 18352 29788 18358
rect 29736 18294 29788 18300
rect 29840 18170 29868 19382
rect 29932 18834 29960 19450
rect 30196 19440 30248 19446
rect 30196 19382 30248 19388
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30012 18896 30064 18902
rect 30012 18838 30064 18844
rect 29920 18828 29972 18834
rect 29920 18770 29972 18776
rect 29920 18692 29972 18698
rect 29920 18634 29972 18640
rect 29932 18426 29960 18634
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 30024 18222 30052 18838
rect 30116 18290 30144 19246
rect 30208 18902 30236 19382
rect 30196 18896 30248 18902
rect 30196 18838 30248 18844
rect 30104 18284 30156 18290
rect 30104 18226 30156 18232
rect 29748 18142 29868 18170
rect 30012 18216 30064 18222
rect 30012 18158 30064 18164
rect 29644 16720 29696 16726
rect 29644 16662 29696 16668
rect 29748 16454 29776 18142
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 29828 17808 29880 17814
rect 29828 17750 29880 17756
rect 29840 17610 29868 17750
rect 30208 17746 30236 18022
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 30012 17604 30064 17610
rect 30012 17546 30064 17552
rect 29736 16448 29788 16454
rect 29736 16390 29788 16396
rect 29552 16176 29604 16182
rect 29552 16118 29604 16124
rect 29564 14482 29592 16118
rect 30024 16046 30052 17546
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30012 16040 30064 16046
rect 30012 15982 30064 15988
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29840 14822 29868 15438
rect 29828 14816 29880 14822
rect 29828 14758 29880 14764
rect 29552 14476 29604 14482
rect 29552 14418 29604 14424
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29736 14272 29788 14278
rect 29736 14214 29788 14220
rect 29748 14074 29776 14214
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29368 13864 29420 13870
rect 29368 13806 29420 13812
rect 29380 13530 29408 13806
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29932 13326 29960 14350
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29274 11248 29330 11257
rect 29274 11183 29330 11192
rect 29748 9518 29776 13262
rect 30116 10266 30144 17070
rect 30300 16658 30328 23054
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 30392 19786 30420 20810
rect 30380 19780 30432 19786
rect 30380 19722 30432 19728
rect 30576 19446 30604 23258
rect 30668 22166 30696 23598
rect 30656 22160 30708 22166
rect 30656 22102 30708 22108
rect 30380 19440 30432 19446
rect 30564 19440 30616 19446
rect 30432 19388 30512 19394
rect 30380 19382 30512 19388
rect 30564 19382 30616 19388
rect 30392 19366 30512 19382
rect 30380 18080 30432 18086
rect 30380 18022 30432 18028
rect 30392 17542 30420 18022
rect 30484 17610 30512 19366
rect 30668 19310 30696 22102
rect 30760 21690 30788 23734
rect 30852 23662 30880 25842
rect 30840 23656 30892 23662
rect 30840 23598 30892 23604
rect 30748 21684 30800 21690
rect 30748 21626 30800 21632
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 30656 19304 30708 19310
rect 30656 19246 30708 19252
rect 31404 18834 31432 19722
rect 31484 19712 31536 19718
rect 31484 19654 31536 19660
rect 31496 19378 31524 19654
rect 31484 19372 31536 19378
rect 31484 19314 31536 19320
rect 31392 18828 31444 18834
rect 31392 18770 31444 18776
rect 31300 18692 31352 18698
rect 31300 18634 31352 18640
rect 30564 18284 30616 18290
rect 30564 18226 30616 18232
rect 30840 18284 30892 18290
rect 30840 18226 30892 18232
rect 30472 17604 30524 17610
rect 30472 17546 30524 17552
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30576 17338 30604 18226
rect 30852 18057 30880 18226
rect 31312 18193 31340 18634
rect 31298 18184 31354 18193
rect 31298 18119 31354 18128
rect 30838 18048 30894 18057
rect 30838 17983 30894 17992
rect 30748 17876 30800 17882
rect 30748 17818 30800 17824
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30472 16448 30524 16454
rect 30472 16390 30524 16396
rect 30484 16182 30512 16390
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30564 15360 30616 15366
rect 30564 15302 30616 15308
rect 30380 15020 30432 15026
rect 30380 14962 30432 14968
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30300 14074 30328 14418
rect 30288 14068 30340 14074
rect 30288 14010 30340 14016
rect 30392 13977 30420 14962
rect 30472 14272 30524 14278
rect 30472 14214 30524 14220
rect 30484 14006 30512 14214
rect 30472 14000 30524 14006
rect 30378 13968 30434 13977
rect 30472 13942 30524 13948
rect 30378 13903 30434 13912
rect 30576 13802 30604 15302
rect 30564 13796 30616 13802
rect 30564 13738 30616 13744
rect 30378 13016 30434 13025
rect 30378 12951 30380 12960
rect 30432 12951 30434 12960
rect 30380 12922 30432 12928
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 29736 9512 29788 9518
rect 29736 9454 29788 9460
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 25136 2576 25188 2582
rect 25136 2518 25188 2524
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 24504 800 24532 2382
rect 25792 800 25820 2382
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 26436 800 26464 2314
rect 26620 1494 26648 2994
rect 26608 1488 26660 1494
rect 26608 1430 26660 1436
rect 27724 800 27752 2994
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28368 800 28396 2246
rect 28460 2106 28488 2382
rect 28448 2100 28500 2106
rect 28448 2042 28500 2048
rect 28828 2038 28856 3062
rect 28908 2916 28960 2922
rect 28908 2858 28960 2864
rect 28920 2378 28948 2858
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 29748 2310 29776 8434
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30392 3194 30420 6734
rect 30380 3188 30432 3194
rect 30380 3130 30432 3136
rect 30668 2774 30696 17478
rect 30760 17066 30788 17818
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31128 17202 31156 17614
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 30748 17060 30800 17066
rect 30748 17002 30800 17008
rect 30840 16720 30892 16726
rect 30840 16662 30892 16668
rect 30852 16114 30880 16662
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 31128 16250 31156 16390
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 30840 16108 30892 16114
rect 30840 16050 30892 16056
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31128 15026 31156 16050
rect 31404 15638 31432 18770
rect 31576 17264 31628 17270
rect 31576 17206 31628 17212
rect 31588 16250 31616 17206
rect 31576 16244 31628 16250
rect 31576 16186 31628 16192
rect 31392 15632 31444 15638
rect 31392 15574 31444 15580
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 31128 14346 31156 14962
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31220 14346 31248 14758
rect 31404 14482 31432 15574
rect 31392 14476 31444 14482
rect 31392 14418 31444 14424
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 31208 14340 31260 14346
rect 31208 14282 31260 14288
rect 30840 12912 30892 12918
rect 30840 12854 30892 12860
rect 30748 12776 30800 12782
rect 30748 12718 30800 12724
rect 30760 12306 30788 12718
rect 30748 12300 30800 12306
rect 30748 12242 30800 12248
rect 30852 8294 30880 12854
rect 31668 12776 31720 12782
rect 31668 12718 31720 12724
rect 31024 12708 31076 12714
rect 31024 12650 31076 12656
rect 30840 8288 30892 8294
rect 30840 8230 30892 8236
rect 31036 6866 31064 12650
rect 31680 12238 31708 12718
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31680 11694 31708 12174
rect 31668 11688 31720 11694
rect 31668 11630 31720 11636
rect 31024 6860 31076 6866
rect 31024 6802 31076 6808
rect 32416 5234 32444 28630
rect 33796 24206 33824 32370
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35544 32026 35572 35566
rect 35912 34746 35940 36722
rect 35900 34740 35952 34746
rect 35900 34682 35952 34688
rect 35532 32020 35584 32026
rect 35532 31962 35584 31968
rect 33876 31816 33928 31822
rect 33876 31758 33928 31764
rect 33888 26042 33916 31758
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33876 26036 33928 26042
rect 33876 25978 33928 25984
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33796 22030 33824 24142
rect 36096 23526 36124 37198
rect 36188 36174 36216 37318
rect 36740 37262 36768 39200
rect 36818 38856 36874 38865
rect 36818 38791 36874 38800
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 36544 37188 36596 37194
rect 36544 37130 36596 37136
rect 36176 36168 36228 36174
rect 36176 36110 36228 36116
rect 36176 36032 36228 36038
rect 36176 35974 36228 35980
rect 36188 32910 36216 35974
rect 36176 32904 36228 32910
rect 36176 32846 36228 32852
rect 36556 26382 36584 37130
rect 36832 36922 36860 38791
rect 37648 37120 37700 37126
rect 37648 37062 37700 37068
rect 36820 36916 36872 36922
rect 36820 36858 36872 36864
rect 37462 36816 37518 36825
rect 37462 36751 37518 36760
rect 37476 36378 37504 36751
rect 37464 36372 37516 36378
rect 37464 36314 37516 36320
rect 37280 35080 37332 35086
rect 37280 35022 37332 35028
rect 37188 34536 37240 34542
rect 37188 34478 37240 34484
rect 37200 34105 37228 34478
rect 37186 34096 37242 34105
rect 37186 34031 37242 34040
rect 37188 31816 37240 31822
rect 37188 31758 37240 31764
rect 37200 31385 37228 31758
rect 37186 31376 37242 31385
rect 37186 31311 37242 31320
rect 37004 29504 37056 29510
rect 37004 29446 37056 29452
rect 37016 28558 37044 29446
rect 37188 29096 37240 29102
rect 37188 29038 37240 29044
rect 37200 28665 37228 29038
rect 37186 28656 37242 28665
rect 37186 28591 37242 28600
rect 37004 28552 37056 28558
rect 37004 28494 37056 28500
rect 36544 26376 36596 26382
rect 36544 26318 36596 26324
rect 36556 25362 36584 26318
rect 36544 25356 36596 25362
rect 36544 25298 36596 25304
rect 36084 23520 36136 23526
rect 36084 23462 36136 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 33784 22024 33836 22030
rect 33784 21966 33836 21972
rect 32680 21956 32732 21962
rect 32680 21898 32732 21904
rect 32692 18766 32720 21898
rect 33600 21888 33652 21894
rect 33600 21830 33652 21836
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 33508 16788 33560 16794
rect 33508 16730 33560 16736
rect 33520 15706 33548 16730
rect 33508 15700 33560 15706
rect 33508 15642 33560 15648
rect 32404 5228 32456 5234
rect 32404 5170 32456 5176
rect 31300 4616 31352 4622
rect 31300 4558 31352 4564
rect 31312 4282 31340 4558
rect 31300 4276 31352 4282
rect 31300 4218 31352 4224
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 30668 2746 30788 2774
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 28816 2032 28868 2038
rect 28816 1974 28868 1980
rect 29932 1426 29960 2382
rect 29000 1420 29052 1426
rect 29000 1362 29052 1368
rect 29920 1420 29972 1426
rect 29920 1362 29972 1368
rect 29012 800 29040 1362
rect 30208 1306 30236 2450
rect 30378 2408 30434 2417
rect 30378 2343 30434 2352
rect 30392 2310 30420 2343
rect 30380 2304 30432 2310
rect 30380 2246 30432 2252
rect 30760 2106 30788 2746
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 30748 2100 30800 2106
rect 30748 2042 30800 2048
rect 30208 1278 30328 1306
rect 30300 800 30328 1278
rect 30944 800 30972 2246
rect 32232 800 32260 2246
rect 32876 800 32904 2994
rect 33612 2446 33640 21830
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34532 17678 34560 18566
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 35900 16108 35952 16114
rect 35900 16050 35952 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 33980 8090 34008 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34060 12232 34112 12238
rect 34060 12174 34112 12180
rect 34072 11898 34100 12174
rect 34060 11892 34112 11898
rect 34060 11834 34112 11840
rect 34796 11824 34848 11830
rect 34796 11766 34848 11772
rect 34808 11082 34836 11766
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35912 11082 35940 16050
rect 37200 14414 37228 16594
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 37200 14074 37228 14350
rect 37188 14068 37240 14074
rect 37188 14010 37240 14016
rect 36452 12844 36504 12850
rect 36452 12786 36504 12792
rect 36464 12442 36492 12786
rect 36452 12436 36504 12442
rect 36452 12378 36504 12384
rect 37292 12374 37320 35022
rect 37464 32360 37516 32366
rect 37464 32302 37516 32308
rect 37476 32065 37504 32302
rect 37462 32056 37518 32065
rect 37462 31991 37518 32000
rect 37556 31816 37608 31822
rect 37556 31758 37608 31764
rect 37372 27532 37424 27538
rect 37372 27474 37424 27480
rect 37384 17746 37412 27474
rect 37464 27464 37516 27470
rect 37464 27406 37516 27412
rect 37476 27305 37504 27406
rect 37462 27296 37518 27305
rect 37462 27231 37518 27240
rect 37568 24818 37596 31758
rect 37660 27878 37688 37062
rect 38028 36854 38056 39200
rect 38290 38176 38346 38185
rect 38290 38111 38346 38120
rect 38016 36848 38068 36854
rect 38016 36790 38068 36796
rect 37832 36576 37884 36582
rect 37832 36518 37884 36524
rect 37740 34536 37792 34542
rect 37740 34478 37792 34484
rect 37648 27872 37700 27878
rect 37648 27814 37700 27820
rect 37752 26586 37780 34478
rect 37740 26580 37792 26586
rect 37740 26522 37792 26528
rect 37646 25256 37702 25265
rect 37646 25191 37648 25200
rect 37700 25191 37702 25200
rect 37648 25162 37700 25168
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 37464 24200 37516 24206
rect 37464 24142 37516 24148
rect 37476 23905 37504 24142
rect 37462 23896 37518 23905
rect 37462 23831 37518 23840
rect 37568 22642 37596 24754
rect 37648 24608 37700 24614
rect 37648 24550 37700 24556
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37556 21548 37608 21554
rect 37556 21490 37608 21496
rect 37372 17740 37424 17746
rect 37372 17682 37424 17688
rect 37464 17128 37516 17134
rect 37462 17096 37464 17105
rect 37516 17096 37518 17105
rect 37462 17031 37518 17040
rect 37372 15496 37424 15502
rect 37372 15438 37424 15444
rect 37384 14618 37412 15438
rect 37372 14612 37424 14618
rect 37372 14554 37424 14560
rect 37280 12368 37332 12374
rect 37280 12310 37332 12316
rect 37464 11688 37516 11694
rect 37462 11656 37464 11665
rect 37516 11656 37518 11665
rect 37462 11591 37518 11600
rect 37568 11098 37596 21490
rect 34796 11076 34848 11082
rect 34796 11018 34848 11024
rect 35900 11076 35952 11082
rect 35900 11018 35952 11024
rect 37476 11070 37596 11098
rect 34428 10056 34480 10062
rect 34428 9998 34480 10004
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 34440 3194 34468 9998
rect 34428 3188 34480 3194
rect 34428 3130 34480 3136
rect 34808 2650 34836 11018
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37200 9625 37228 9998
rect 37186 9616 37242 9625
rect 37186 9551 37242 9560
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 37476 7546 37504 11070
rect 37556 9104 37608 9110
rect 37556 9046 37608 9052
rect 37464 7540 37516 7546
rect 37464 7482 37516 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35716 6792 35768 6798
rect 35716 6734 35768 6740
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35728 3670 35756 6734
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 35820 3738 35848 6258
rect 37568 5914 37596 9046
rect 37556 5908 37608 5914
rect 37556 5850 37608 5856
rect 37556 5568 37608 5574
rect 37556 5510 37608 5516
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 35808 3732 35860 3738
rect 35808 3674 35860 3680
rect 35716 3664 35768 3670
rect 35716 3606 35768 3612
rect 36912 3052 36964 3058
rect 36912 2994 36964 3000
rect 36924 2825 36952 2994
rect 36910 2816 36966 2825
rect 34934 2748 35242 2757
rect 36910 2751 36966 2760
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 33520 800 33548 2246
rect 34808 800 34836 2314
rect 35452 800 35480 2314
rect 36728 2304 36780 2310
rect 36728 2246 36780 2252
rect 36740 800 36768 2246
rect 37200 2145 37228 3878
rect 37280 3528 37332 3534
rect 37280 3470 37332 3476
rect 37186 2136 37242 2145
rect 37186 2071 37242 2080
rect 8116 750 8168 756
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12254 200 12310 800
rect 12898 200 12954 800
rect 14186 200 14242 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 17406 200 17462 800
rect 18694 200 18750 800
rect 19338 200 19394 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 21914 200 21970 800
rect 23202 200 23258 800
rect 23846 200 23902 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 26422 200 26478 800
rect 27710 200 27766 800
rect 28354 200 28410 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 32862 200 32918 800
rect 33506 200 33562 800
rect 34794 200 34850 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 37292 105 37320 3470
rect 37568 3058 37596 5510
rect 37556 3052 37608 3058
rect 37556 2994 37608 3000
rect 37660 2514 37688 24550
rect 37740 24200 37792 24206
rect 37740 24142 37792 24148
rect 37752 15570 37780 24142
rect 37844 19854 37872 36518
rect 38198 36136 38254 36145
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 38304 35290 38332 38111
rect 38672 36650 38700 39200
rect 38660 36644 38712 36650
rect 38660 36586 38712 36592
rect 39316 35766 39344 39200
rect 39304 35760 39356 35766
rect 39304 35702 39356 35708
rect 38292 35284 38344 35290
rect 38292 35226 38344 35232
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 38120 33425 38148 33458
rect 38106 33416 38162 33425
rect 38106 33351 38162 33360
rect 38106 30696 38162 30705
rect 38106 30631 38108 30640
rect 38160 30631 38162 30640
rect 38108 30602 38160 30608
rect 38200 30592 38252 30598
rect 38200 30534 38252 30540
rect 38212 27062 38240 30534
rect 38292 29640 38344 29646
rect 38292 29582 38344 29588
rect 38304 29345 38332 29582
rect 38290 29336 38346 29345
rect 38290 29271 38346 29280
rect 38200 27056 38252 27062
rect 38200 26998 38252 27004
rect 38292 26988 38344 26994
rect 38292 26930 38344 26936
rect 38304 26625 38332 26930
rect 38290 26616 38346 26625
rect 38290 26551 38346 26560
rect 38200 26512 38252 26518
rect 38200 26454 38252 26460
rect 38212 25945 38240 26454
rect 38198 25936 38254 25945
rect 38198 25871 38254 25880
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38212 24585 38240 25094
rect 38198 24576 38254 24585
rect 38198 24511 38254 24520
rect 38384 24268 38436 24274
rect 38384 24210 38436 24216
rect 38016 22636 38068 22642
rect 38016 22578 38068 22584
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37844 19378 37872 19790
rect 37924 19508 37976 19514
rect 37924 19450 37976 19456
rect 37832 19372 37884 19378
rect 37832 19314 37884 19320
rect 37740 15564 37792 15570
rect 37740 15506 37792 15512
rect 37752 15026 37780 15506
rect 37740 15020 37792 15026
rect 37740 14962 37792 14968
rect 37936 14414 37964 19450
rect 38028 16250 38056 22578
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38304 21865 38332 21966
rect 38290 21856 38346 21865
rect 38290 21791 38346 21800
rect 38198 21720 38254 21729
rect 38198 21655 38200 21664
rect 38252 21655 38254 21664
rect 38200 21626 38252 21632
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 38120 21185 38148 21490
rect 38106 21176 38162 21185
rect 38106 21111 38162 21120
rect 38292 19848 38344 19854
rect 38290 19816 38292 19825
rect 38344 19816 38346 19825
rect 38290 19751 38346 19760
rect 38292 18760 38344 18766
rect 38292 18702 38344 18708
rect 38304 18465 38332 18702
rect 38290 18456 38346 18465
rect 38290 18391 38346 18400
rect 38108 16516 38160 16522
rect 38108 16458 38160 16464
rect 38120 16425 38148 16458
rect 38106 16416 38162 16425
rect 38106 16351 38162 16360
rect 38016 16244 38068 16250
rect 38016 16186 38068 16192
rect 38200 15360 38252 15366
rect 38200 15302 38252 15308
rect 38212 15065 38240 15302
rect 38198 15056 38254 15065
rect 38198 14991 38254 15000
rect 38016 14816 38068 14822
rect 38016 14758 38068 14764
rect 37924 14408 37976 14414
rect 37924 14350 37976 14356
rect 37740 13932 37792 13938
rect 37740 13874 37792 13880
rect 37752 10062 37780 13874
rect 37740 10056 37792 10062
rect 37740 9998 37792 10004
rect 37752 5710 37780 9998
rect 38028 8974 38056 14758
rect 38198 14376 38254 14385
rect 38198 14311 38254 14320
rect 38212 14278 38240 14311
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 38292 13932 38344 13938
rect 38292 13874 38344 13880
rect 38304 13705 38332 13874
rect 38290 13696 38346 13705
rect 38290 13631 38346 13640
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 38396 10742 38424 24210
rect 38384 10736 38436 10742
rect 38384 10678 38436 10684
rect 38108 10668 38160 10674
rect 38108 10610 38160 10616
rect 38120 10305 38148 10610
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 38292 7880 38344 7886
rect 38292 7822 38344 7828
rect 38304 7585 38332 7822
rect 38290 7576 38346 7585
rect 38290 7511 38346 7520
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38120 6905 38148 7346
rect 38106 6896 38162 6905
rect 38106 6831 38162 6840
rect 38016 6180 38068 6186
rect 38016 6122 38068 6128
rect 37740 5704 37792 5710
rect 37740 5646 37792 5652
rect 38028 4146 38056 6122
rect 38200 5568 38252 5574
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38198 5471 38254 5480
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 38212 4865 38240 4966
rect 38198 4856 38254 4865
rect 38198 4791 38254 4800
rect 38200 4480 38252 4486
rect 38200 4422 38252 4428
rect 38212 4185 38240 4422
rect 38198 4176 38254 4185
rect 38016 4140 38068 4146
rect 38198 4111 38254 4120
rect 38016 4082 38068 4088
rect 39304 3528 39356 3534
rect 39304 3470 39356 3476
rect 38292 3460 38344 3466
rect 38292 3402 38344 3408
rect 38016 2848 38068 2854
rect 38016 2790 38068 2796
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 37384 800 37412 2382
rect 37752 2038 37780 2382
rect 37740 2032 37792 2038
rect 37740 1974 37792 1980
rect 38028 800 38056 2790
rect 37370 200 37426 800
rect 38014 200 38070 800
rect 38304 785 38332 3402
rect 39316 800 39344 3470
rect 38290 776 38346 785
rect 38290 711 38346 720
rect 39302 200 39358 800
rect 37278 96 37334 105
rect 37278 31 37334 40
<< via2 >>
rect 3054 39480 3110 39536
rect 2870 38800 2926 38856
rect 1766 36760 1822 36816
rect 1582 35400 1638 35456
rect 1766 34040 1822 34096
rect 110 23432 166 23488
rect 18 19760 74 19816
rect 1398 30368 1454 30424
rect 1766 32716 1768 32736
rect 1768 32716 1820 32736
rect 1820 32716 1822 32736
rect 1766 32680 1822 32716
rect 1766 32000 1822 32056
rect 1766 30640 1822 30696
rect 1766 29280 1822 29336
rect 1766 27940 1822 27976
rect 1766 27920 1768 27940
rect 1768 27920 1820 27940
rect 1820 27920 1822 27940
rect 1766 27276 1768 27296
rect 1768 27276 1820 27296
rect 1820 27276 1822 27296
rect 1766 27240 1822 27276
rect 1766 25200 1822 25256
rect 3146 37440 3202 37496
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 2042 30368 2098 30424
rect 2042 25064 2098 25120
rect 2594 29008 2650 29064
rect 2318 25916 2320 25936
rect 2320 25916 2372 25936
rect 2372 25916 2374 25936
rect 2318 25880 2374 25916
rect 1490 23024 1546 23080
rect 1582 22480 1638 22536
rect 1950 21528 2006 21584
rect 1766 18400 1822 18456
rect 1674 15680 1730 15736
rect 1398 9596 1400 9616
rect 1400 9596 1452 9616
rect 1452 9596 1454 9616
rect 1398 9560 1454 9596
rect 1766 13676 1768 13696
rect 1768 13676 1820 13696
rect 1820 13676 1822 13696
rect 1766 13640 1822 13676
rect 2686 28464 2742 28520
rect 2410 21800 2466 21856
rect 2410 16632 2466 16688
rect 2226 13096 2282 13152
rect 3054 26016 3110 26072
rect 3054 24792 3110 24848
rect 3238 23704 3294 23760
rect 3422 24556 3424 24576
rect 3424 24556 3476 24576
rect 3476 24556 3478 24576
rect 3422 24520 3478 24556
rect 3054 20848 3110 20904
rect 2870 19352 2926 19408
rect 2502 11872 2558 11928
rect 1766 7540 1822 7576
rect 1766 7520 1768 7540
rect 1768 7520 1820 7540
rect 1820 7520 1822 7540
rect 1674 5480 1730 5536
rect 2318 6432 2374 6488
rect 2318 6332 2320 6352
rect 2320 6332 2372 6352
rect 2372 6332 2374 6352
rect 2318 6296 2374 6332
rect 3698 29960 3754 30016
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4434 30368 4490 30424
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 3330 21256 3386 21312
rect 3238 15680 3294 15736
rect 2870 10240 2926 10296
rect 2410 4256 2466 4312
rect 2962 8744 3018 8800
rect 3698 21936 3754 21992
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4618 28600 4674 28656
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27648 4122 27704
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 26288 4122 26344
rect 4066 25744 4122 25800
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4434 25200 4490 25256
rect 4158 24656 4214 24712
rect 5170 30368 5226 30424
rect 4710 26016 4766 26072
rect 5078 27104 5134 27160
rect 4986 26968 5042 27024
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4066 23860 4122 23896
rect 4066 23840 4068 23860
rect 4068 23840 4120 23860
rect 4120 23840 4122 23860
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3974 21120 4030 21176
rect 4618 21664 4674 21720
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 20440 4122 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 3698 19896 3754 19952
rect 4986 24928 5042 24984
rect 4802 21936 4858 21992
rect 4894 21664 4950 21720
rect 4802 20576 4858 20632
rect 5078 24384 5134 24440
rect 5078 23160 5134 23216
rect 5446 26696 5502 26752
rect 5262 23432 5318 23488
rect 5170 21256 5226 21312
rect 5170 21120 5226 21176
rect 5078 20712 5134 20768
rect 4894 19760 4950 19816
rect 4802 19352 4858 19408
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4710 18536 4766 18592
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4066 17720 4122 17776
rect 3882 16496 3938 16552
rect 3790 12960 3846 13016
rect 3698 12144 3754 12200
rect 3422 11228 3424 11248
rect 3424 11228 3476 11248
rect 3476 11228 3478 11248
rect 3422 11192 3478 11228
rect 3238 10124 3294 10160
rect 3238 10104 3240 10124
rect 3240 10104 3292 10124
rect 3292 10104 3294 10124
rect 3882 12280 3938 12336
rect 4250 17176 4306 17232
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4066 16360 4122 16416
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4526 14048 4582 14104
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4158 12960 4214 13016
rect 4526 12688 4582 12744
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3974 12008 4030 12064
rect 3882 11056 3938 11112
rect 3882 10920 3938 10976
rect 3974 9596 3976 9616
rect 3976 9596 4028 9616
rect 4028 9596 4030 9616
rect 3974 9560 4030 9596
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4434 9832 4490 9888
rect 5170 15952 5226 16008
rect 5078 14728 5134 14784
rect 4802 10920 4858 10976
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 2962 4256 3018 4312
rect 2962 3576 3018 3632
rect 2962 3304 3018 3360
rect 3698 6180 3754 6216
rect 3698 6160 3700 6180
rect 3700 6160 3752 6180
rect 3752 6160 3754 6180
rect 4342 8900 4398 8936
rect 4342 8880 4344 8900
rect 4344 8880 4396 8900
rect 4396 8880 4398 8900
rect 3974 8336 4030 8392
rect 3882 8236 3884 8256
rect 3884 8236 3936 8256
rect 3936 8236 3938 8256
rect 3882 8200 3938 8236
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4066 7248 4122 7304
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4802 6024 4858 6080
rect 4710 5888 4766 5944
rect 3882 5072 3938 5128
rect 3514 3032 3570 3088
rect 3974 4120 4030 4176
rect 3790 3440 3846 3496
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4710 4664 4766 4720
rect 5446 22888 5502 22944
rect 5722 26832 5778 26888
rect 5354 19624 5410 19680
rect 5354 18708 5356 18728
rect 5356 18708 5408 18728
rect 5408 18708 5410 18728
rect 5354 18672 5410 18708
rect 5998 26288 6054 26344
rect 5998 25064 6054 25120
rect 5906 24928 5962 24984
rect 5906 24012 5908 24032
rect 5908 24012 5960 24032
rect 5960 24012 5962 24032
rect 5906 23976 5962 24012
rect 5722 23024 5778 23080
rect 5446 16632 5502 16688
rect 5354 13232 5410 13288
rect 5078 12416 5134 12472
rect 5998 22208 6054 22264
rect 5998 21936 6054 21992
rect 6274 25336 6330 25392
rect 5998 17176 6054 17232
rect 5630 14048 5686 14104
rect 5446 12824 5502 12880
rect 5446 11464 5502 11520
rect 7010 29144 7066 29200
rect 7010 27648 7066 27704
rect 6642 26856 6644 26888
rect 6644 26856 6696 26888
rect 6696 26856 6698 26888
rect 6642 26832 6698 26856
rect 6550 23432 6606 23488
rect 6826 26016 6882 26072
rect 6918 25780 6920 25800
rect 6920 25780 6972 25800
rect 6972 25780 6974 25800
rect 6918 25744 6974 25780
rect 6734 24520 6790 24576
rect 6734 23296 6790 23352
rect 6642 21392 6698 21448
rect 6458 20168 6514 20224
rect 6366 19488 6422 19544
rect 6274 18808 6330 18864
rect 6642 20032 6698 20088
rect 6366 15036 6368 15056
rect 6368 15036 6420 15056
rect 6420 15036 6422 15056
rect 6366 15000 6422 15036
rect 6918 23840 6974 23896
rect 9126 36488 9182 36544
rect 8850 30132 8852 30152
rect 8852 30132 8904 30152
rect 8904 30132 8906 30152
rect 8850 30096 8906 30132
rect 7378 26288 7434 26344
rect 7286 25744 7342 25800
rect 7102 24132 7158 24168
rect 7102 24112 7104 24132
rect 7104 24112 7156 24132
rect 7156 24112 7158 24132
rect 7562 23976 7618 24032
rect 7746 29008 7802 29064
rect 7746 25336 7802 25392
rect 7746 24248 7802 24304
rect 6826 20984 6882 21040
rect 6918 17720 6974 17776
rect 6918 17584 6974 17640
rect 6734 16088 6790 16144
rect 5906 10376 5962 10432
rect 5630 9696 5686 9752
rect 5446 8880 5502 8936
rect 5354 8064 5410 8120
rect 5906 10104 5962 10160
rect 5814 7948 5870 7984
rect 5814 7928 5816 7948
rect 5816 7928 5868 7948
rect 5868 7928 5870 7948
rect 5078 5480 5134 5536
rect 4250 3168 4306 3224
rect 3974 2760 4030 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4618 2524 4620 2544
rect 4620 2524 4672 2544
rect 4672 2524 4674 2544
rect 4618 2488 4674 2524
rect 5354 3052 5410 3088
rect 5354 3032 5356 3052
rect 5356 3032 5408 3052
rect 5408 3032 5410 3052
rect 5998 8200 6054 8256
rect 5722 6160 5778 6216
rect 5262 2624 5318 2680
rect 5538 2896 5594 2952
rect 6090 5344 6146 5400
rect 5998 4120 6054 4176
rect 5170 1808 5226 1864
rect 6274 9424 6330 9480
rect 7470 23704 7526 23760
rect 7286 21936 7342 21992
rect 7102 19216 7158 19272
rect 7194 17856 7250 17912
rect 6826 14340 6882 14376
rect 6826 14320 6828 14340
rect 6828 14320 6880 14340
rect 6880 14320 6882 14340
rect 6826 14184 6882 14240
rect 6734 13504 6790 13560
rect 6918 12960 6974 13016
rect 7010 12144 7066 12200
rect 6734 11192 6790 11248
rect 6642 10648 6698 10704
rect 6458 7384 6514 7440
rect 6826 9288 6882 9344
rect 6826 9052 6828 9072
rect 6828 9052 6880 9072
rect 6880 9052 6882 9072
rect 6826 9016 6882 9052
rect 6458 5616 6514 5672
rect 6550 3984 6606 4040
rect 6366 2760 6422 2816
rect 6090 2216 6146 2272
rect 6550 2896 6606 2952
rect 7562 22072 7618 22128
rect 7470 21664 7526 21720
rect 7470 21256 7526 21312
rect 7378 12008 7434 12064
rect 7562 20440 7618 20496
rect 8298 29280 8354 29336
rect 8666 29280 8722 29336
rect 8850 29280 8906 29336
rect 8206 26868 8208 26888
rect 8208 26868 8260 26888
rect 8260 26868 8262 26888
rect 8206 26832 8262 26868
rect 8482 28076 8538 28112
rect 8482 28056 8484 28076
rect 8484 28056 8536 28076
rect 8536 28056 8538 28076
rect 8390 27376 8446 27432
rect 7838 21664 7894 21720
rect 7654 19352 7710 19408
rect 7746 19252 7748 19272
rect 7748 19252 7800 19272
rect 7800 19252 7802 19272
rect 7746 19216 7802 19252
rect 7838 17992 7894 18048
rect 8114 25200 8170 25256
rect 8114 24384 8170 24440
rect 8114 23432 8170 23488
rect 8022 22208 8078 22264
rect 8022 22072 8078 22128
rect 8482 24248 8538 24304
rect 8758 27648 8814 27704
rect 8758 27412 8760 27432
rect 8760 27412 8812 27432
rect 8812 27412 8814 27432
rect 8758 27376 8814 27412
rect 8850 25744 8906 25800
rect 8206 21120 8262 21176
rect 8206 20712 8262 20768
rect 8666 21936 8722 21992
rect 8574 21800 8630 21856
rect 8206 19080 8262 19136
rect 7562 14728 7618 14784
rect 7194 8608 7250 8664
rect 6826 6432 6882 6488
rect 6918 5616 6974 5672
rect 7102 5364 7158 5400
rect 7102 5344 7104 5364
rect 7104 5344 7156 5364
rect 7156 5344 7158 5364
rect 7378 9968 7434 10024
rect 7286 5208 7342 5264
rect 7286 4528 7342 4584
rect 7010 4392 7066 4448
rect 7286 3984 7342 4040
rect 7562 9152 7618 9208
rect 7470 6976 7526 7032
rect 6826 2488 6882 2544
rect 6458 1400 6514 1456
rect 7930 15408 7986 15464
rect 8666 20304 8722 20360
rect 9402 28500 9404 28520
rect 9404 28500 9456 28520
rect 9456 28500 9458 28520
rect 9402 28464 9458 28500
rect 8942 23840 8998 23896
rect 8850 23432 8906 23488
rect 8850 21936 8906 21992
rect 8666 18400 8722 18456
rect 8574 18164 8576 18184
rect 8576 18164 8628 18184
rect 8628 18164 8630 18184
rect 8574 18128 8630 18164
rect 8574 17992 8630 18048
rect 8574 17312 8630 17368
rect 8206 16768 8262 16824
rect 7838 15156 7894 15192
rect 7838 15136 7840 15156
rect 7840 15136 7892 15156
rect 7892 15136 7894 15156
rect 8022 14864 8078 14920
rect 7746 11872 7802 11928
rect 7746 11736 7802 11792
rect 7930 12008 7986 12064
rect 8206 14728 8262 14784
rect 8114 12552 8170 12608
rect 8574 16632 8630 16688
rect 8758 16360 8814 16416
rect 8850 15816 8906 15872
rect 8574 13368 8630 13424
rect 8390 12164 8446 12200
rect 8390 12144 8392 12164
rect 8392 12144 8444 12164
rect 8444 12144 8446 12164
rect 8390 11600 8446 11656
rect 8206 11464 8262 11520
rect 7930 11056 7986 11112
rect 7838 8608 7894 8664
rect 7746 7384 7802 7440
rect 7930 7420 7932 7440
rect 7932 7420 7984 7440
rect 7984 7420 7986 7440
rect 7930 7384 7986 7420
rect 7746 4664 7802 4720
rect 7746 3848 7802 3904
rect 7930 3712 7986 3768
rect 8298 10668 8354 10704
rect 8298 10648 8300 10668
rect 8300 10648 8352 10668
rect 8352 10648 8354 10668
rect 8206 7656 8262 7712
rect 8114 5616 8170 5672
rect 8574 12280 8630 12336
rect 8574 12008 8630 12064
rect 8666 10920 8722 10976
rect 8574 9832 8630 9888
rect 8758 9696 8814 9752
rect 8482 9424 8538 9480
rect 8482 5344 8538 5400
rect 8298 4800 8354 4856
rect 8758 8608 8814 8664
rect 8666 7792 8722 7848
rect 8758 7520 8814 7576
rect 8666 5752 8722 5808
rect 8666 5344 8722 5400
rect 9126 24928 9182 24984
rect 9126 24692 9128 24712
rect 9128 24692 9180 24712
rect 9180 24692 9182 24712
rect 9126 24656 9182 24692
rect 9310 23296 9366 23352
rect 9862 29960 9918 30016
rect 9770 29552 9826 29608
rect 9954 29688 10010 29744
rect 10138 29416 10194 29472
rect 9678 28192 9734 28248
rect 9586 28056 9642 28112
rect 9586 27648 9642 27704
rect 9494 26560 9550 26616
rect 9954 27648 10010 27704
rect 10598 29960 10654 30016
rect 10598 29824 10654 29880
rect 10782 29824 10838 29880
rect 10782 29572 10838 29608
rect 10782 29552 10784 29572
rect 10784 29552 10836 29572
rect 10836 29552 10838 29572
rect 10506 28736 10562 28792
rect 9770 26152 9826 26208
rect 9586 25064 9642 25120
rect 9126 21392 9182 21448
rect 9310 21256 9366 21312
rect 9034 20576 9090 20632
rect 9218 20576 9274 20632
rect 9862 24928 9918 24984
rect 9678 23976 9734 24032
rect 9770 23024 9826 23080
rect 9678 20304 9734 20360
rect 9586 19896 9642 19952
rect 9494 19760 9550 19816
rect 9034 19352 9090 19408
rect 9586 19216 9642 19272
rect 9494 18944 9550 19000
rect 9218 18536 9274 18592
rect 9034 17856 9090 17912
rect 9402 18128 9458 18184
rect 9126 16632 9182 16688
rect 9218 13640 9274 13696
rect 8942 10104 8998 10160
rect 8942 9696 8998 9752
rect 8850 4936 8906 4992
rect 9218 13232 9274 13288
rect 9310 9424 9366 9480
rect 9034 7520 9090 7576
rect 9034 6704 9090 6760
rect 9126 6568 9182 6624
rect 8206 4256 8262 4312
rect 8206 3168 8262 3224
rect 8482 3984 8538 4040
rect 9310 6296 9366 6352
rect 9586 17312 9642 17368
rect 9494 16224 9550 16280
rect 10230 26832 10286 26888
rect 10046 23840 10102 23896
rect 9954 23704 10010 23760
rect 10046 21664 10102 21720
rect 9954 19352 10010 19408
rect 9862 18536 9918 18592
rect 10230 23976 10286 24032
rect 10782 28464 10838 28520
rect 10690 27648 10746 27704
rect 12070 30368 12126 30424
rect 11886 30252 11942 30288
rect 11886 30232 11888 30252
rect 11888 30232 11940 30252
rect 11940 30232 11942 30252
rect 12254 30096 12310 30152
rect 12162 29144 12218 29200
rect 10966 26424 11022 26480
rect 10506 21800 10562 21856
rect 10782 23296 10838 23352
rect 10506 21528 10562 21584
rect 10690 21528 10746 21584
rect 10230 19760 10286 19816
rect 10138 18808 10194 18864
rect 9862 17040 9918 17096
rect 9678 15308 9680 15328
rect 9680 15308 9732 15328
rect 9732 15308 9734 15328
rect 9678 15272 9734 15308
rect 9586 15136 9642 15192
rect 10046 15272 10102 15328
rect 9862 15136 9918 15192
rect 9494 13232 9550 13288
rect 9494 12860 9496 12880
rect 9496 12860 9548 12880
rect 9548 12860 9550 12880
rect 9494 12824 9550 12860
rect 10046 13912 10102 13968
rect 9494 6568 9550 6624
rect 9034 3984 9090 4040
rect 9034 3576 9090 3632
rect 8390 1944 8446 2000
rect 8298 1672 8354 1728
rect 3514 756 3516 776
rect 3516 756 3568 776
rect 3568 756 3570 776
rect 3514 720 3570 756
rect 9218 3576 9274 3632
rect 9678 10512 9734 10568
rect 9678 8064 9734 8120
rect 9678 7112 9734 7168
rect 9862 8064 9918 8120
rect 9770 4936 9826 4992
rect 9678 4800 9734 4856
rect 9678 3440 9734 3496
rect 10138 11600 10194 11656
rect 10046 9424 10102 9480
rect 10046 6568 10102 6624
rect 10046 5364 10102 5400
rect 10046 5344 10048 5364
rect 10048 5344 10100 5364
rect 10100 5344 10102 5364
rect 10690 21392 10746 21448
rect 10598 19896 10654 19952
rect 11242 26016 11298 26072
rect 11150 25472 11206 25528
rect 11058 24656 11114 24712
rect 11058 24520 11114 24576
rect 11058 23432 11114 23488
rect 11242 23296 11298 23352
rect 11242 22480 11298 22536
rect 10874 21392 10930 21448
rect 10874 20984 10930 21040
rect 11058 21936 11114 21992
rect 10874 19292 10930 19348
rect 10598 14048 10654 14104
rect 10506 13776 10562 13832
rect 10506 10648 10562 10704
rect 11702 24384 11758 24440
rect 11518 22616 11574 22672
rect 11426 22344 11482 22400
rect 11334 21936 11390 21992
rect 11242 21392 11298 21448
rect 11334 19488 11390 19544
rect 11334 19352 11390 19408
rect 11150 19216 11206 19272
rect 11058 18944 11114 19000
rect 10966 18128 11022 18184
rect 10874 17856 10930 17912
rect 10782 17312 10838 17368
rect 10782 16224 10838 16280
rect 10966 15136 11022 15192
rect 11242 17856 11298 17912
rect 11978 26444 12034 26480
rect 11978 26424 11980 26444
rect 11980 26424 12032 26444
rect 12032 26424 12034 26444
rect 12530 28736 12586 28792
rect 12438 28076 12494 28112
rect 12438 28056 12440 28076
rect 12440 28056 12492 28076
rect 12492 28056 12494 28076
rect 13082 29280 13138 29336
rect 13358 28484 13414 28520
rect 13358 28464 13360 28484
rect 13360 28464 13412 28484
rect 13412 28464 13414 28484
rect 13082 27376 13138 27432
rect 12806 26424 12862 26480
rect 12162 23432 12218 23488
rect 11886 21936 11942 21992
rect 11886 21392 11942 21448
rect 11610 19488 11666 19544
rect 11426 15544 11482 15600
rect 10782 14456 10838 14512
rect 10782 12416 10838 12472
rect 10782 11872 10838 11928
rect 10782 10920 10838 10976
rect 10782 10512 10838 10568
rect 11978 20304 12034 20360
rect 11702 17856 11758 17912
rect 12254 23044 12310 23080
rect 12254 23024 12256 23044
rect 12256 23024 12308 23044
rect 12308 23024 12310 23044
rect 12438 22772 12494 22808
rect 12438 22752 12440 22772
rect 12440 22752 12492 22772
rect 12492 22752 12494 22772
rect 12254 22652 12256 22672
rect 12256 22652 12308 22672
rect 12308 22652 12310 22672
rect 12622 23432 12678 23488
rect 12254 22616 12310 22652
rect 12254 22344 12310 22400
rect 12346 20848 12402 20904
rect 12530 20984 12586 21040
rect 12530 20884 12532 20904
rect 12532 20884 12584 20904
rect 12584 20884 12586 20904
rect 12530 20848 12586 20884
rect 11886 19080 11942 19136
rect 11886 18808 11942 18864
rect 11886 18536 11942 18592
rect 11702 17448 11758 17504
rect 11794 17176 11850 17232
rect 11794 15680 11850 15736
rect 12070 18808 12126 18864
rect 12070 18400 12126 18456
rect 12530 19760 12586 19816
rect 12346 18420 12402 18456
rect 12346 18400 12348 18420
rect 12348 18400 12400 18420
rect 12400 18400 12402 18420
rect 12162 17604 12218 17640
rect 12162 17584 12164 17604
rect 12164 17584 12216 17604
rect 12216 17584 12218 17604
rect 12070 17448 12126 17504
rect 12254 16904 12310 16960
rect 12162 16632 12218 16688
rect 12438 17856 12494 17912
rect 12806 22344 12862 22400
rect 12714 22208 12770 22264
rect 12990 24792 13046 24848
rect 13450 26968 13506 27024
rect 13634 26832 13690 26888
rect 13266 23024 13322 23080
rect 13174 22092 13230 22128
rect 13174 22072 13176 22092
rect 13176 22072 13228 22092
rect 13228 22072 13230 22092
rect 13082 21528 13138 21584
rect 12990 21256 13046 21312
rect 12898 19760 12954 19816
rect 12898 18808 12954 18864
rect 13082 19896 13138 19952
rect 13542 26696 13598 26752
rect 13542 23296 13598 23352
rect 13910 24384 13966 24440
rect 13818 23840 13874 23896
rect 13726 23568 13782 23624
rect 13542 22652 13544 22672
rect 13544 22652 13596 22672
rect 13596 22652 13598 22672
rect 13542 22616 13598 22652
rect 13910 22616 13966 22672
rect 13818 21528 13874 21584
rect 13726 21392 13782 21448
rect 13542 20440 13598 20496
rect 13726 20440 13782 20496
rect 13818 19896 13874 19952
rect 13358 18808 13414 18864
rect 13358 18536 13414 18592
rect 12070 16360 12126 16416
rect 11702 15272 11758 15328
rect 11794 14592 11850 14648
rect 11058 12824 11114 12880
rect 11058 11328 11114 11384
rect 11150 10648 11206 10704
rect 11150 10512 11206 10568
rect 11058 9832 11114 9888
rect 10598 8608 10654 8664
rect 10598 7792 10654 7848
rect 10414 6976 10470 7032
rect 10414 6568 10470 6624
rect 10322 5480 10378 5536
rect 10874 9016 10930 9072
rect 10874 8608 10930 8664
rect 11426 13232 11482 13288
rect 11334 10376 11390 10432
rect 11334 10240 11390 10296
rect 11242 9036 11298 9072
rect 11242 9016 11244 9036
rect 11244 9016 11296 9036
rect 11296 9016 11298 9036
rect 11610 13368 11666 13424
rect 11610 12824 11666 12880
rect 11702 11636 11704 11656
rect 11704 11636 11756 11656
rect 11756 11636 11758 11656
rect 11702 11600 11758 11636
rect 11702 10784 11758 10840
rect 11518 10512 11574 10568
rect 11518 10240 11574 10296
rect 11334 8336 11390 8392
rect 10874 6976 10930 7032
rect 11058 6976 11114 7032
rect 10598 6296 10654 6352
rect 10782 6296 10838 6352
rect 10322 3440 10378 3496
rect 10690 3440 10746 3496
rect 11242 5636 11298 5672
rect 11242 5616 11244 5636
rect 11244 5616 11296 5636
rect 11296 5616 11298 5636
rect 11242 5208 11298 5264
rect 11702 9016 11758 9072
rect 12162 15272 12218 15328
rect 12070 14864 12126 14920
rect 11886 13368 11942 13424
rect 11886 10532 11942 10568
rect 11886 10512 11888 10532
rect 11888 10512 11940 10532
rect 11940 10512 11942 10532
rect 12438 15816 12494 15872
rect 12438 14456 12494 14512
rect 12254 13776 12310 13832
rect 12898 17448 12954 17504
rect 12898 17312 12954 17368
rect 12806 15816 12862 15872
rect 12806 15544 12862 15600
rect 12714 14728 12770 14784
rect 12438 12280 12494 12336
rect 12438 11328 12494 11384
rect 12806 12416 12862 12472
rect 13358 17720 13414 17776
rect 13266 17040 13322 17096
rect 13266 16632 13322 16688
rect 13266 15680 13322 15736
rect 13174 15544 13230 15600
rect 13082 15408 13138 15464
rect 13726 19352 13782 19408
rect 13910 18536 13966 18592
rect 13726 17312 13782 17368
rect 13910 16632 13966 16688
rect 13726 15136 13782 15192
rect 13266 13504 13322 13560
rect 12254 10784 12310 10840
rect 12530 10104 12586 10160
rect 11886 9016 11942 9072
rect 11886 8608 11942 8664
rect 12898 10920 12954 10976
rect 12806 10104 12862 10160
rect 12806 9968 12862 10024
rect 13266 12280 13322 12336
rect 13634 13504 13690 13560
rect 14554 27512 14610 27568
rect 16302 30096 16358 30152
rect 15014 29688 15070 29744
rect 14554 24928 14610 24984
rect 14646 24656 14702 24712
rect 14186 20984 14242 21040
rect 14094 19488 14150 19544
rect 14094 19352 14150 19408
rect 14278 17992 14334 18048
rect 14094 17856 14150 17912
rect 14462 23044 14518 23080
rect 14462 23024 14464 23044
rect 14464 23024 14516 23044
rect 14516 23024 14518 23044
rect 14462 22072 14518 22128
rect 14462 20712 14518 20768
rect 14094 17176 14150 17232
rect 14278 17312 14334 17368
rect 14186 16904 14242 16960
rect 14370 17176 14426 17232
rect 14002 14728 14058 14784
rect 13818 13776 13874 13832
rect 13542 11600 13598 11656
rect 13542 11056 13598 11112
rect 13450 10104 13506 10160
rect 13266 8200 13322 8256
rect 12898 7964 12900 7984
rect 12900 7964 12952 7984
rect 12952 7964 12954 7984
rect 12898 7928 12954 7964
rect 11886 6976 11942 7032
rect 11610 5516 11612 5536
rect 11612 5516 11664 5536
rect 11664 5516 11666 5536
rect 11610 5480 11666 5516
rect 12162 6568 12218 6624
rect 11702 5072 11758 5128
rect 10230 2080 10286 2136
rect 10874 2624 10930 2680
rect 10966 2352 11022 2408
rect 12070 4664 12126 4720
rect 12622 6876 12624 6896
rect 12624 6876 12676 6896
rect 12676 6876 12678 6896
rect 12622 6840 12678 6876
rect 12806 6840 12862 6896
rect 12346 5636 12402 5672
rect 12346 5616 12348 5636
rect 12348 5616 12400 5636
rect 12400 5616 12402 5636
rect 12530 5616 12586 5672
rect 12530 5364 12586 5400
rect 12530 5344 12532 5364
rect 12532 5344 12584 5364
rect 12584 5344 12586 5364
rect 12530 4800 12586 4856
rect 12346 4664 12402 4720
rect 12162 4120 12218 4176
rect 12530 3984 12586 4040
rect 12530 3712 12586 3768
rect 12806 4140 12862 4176
rect 12806 4120 12808 4140
rect 12808 4120 12860 4140
rect 12860 4120 12862 4140
rect 13266 7928 13322 7984
rect 13082 5752 13138 5808
rect 13082 5480 13138 5536
rect 13818 12144 13874 12200
rect 13818 11328 13874 11384
rect 14002 11076 14058 11112
rect 14002 11056 14004 11076
rect 14004 11056 14056 11076
rect 14056 11056 14058 11076
rect 13726 10784 13782 10840
rect 14002 10920 14058 10976
rect 13818 9968 13874 10024
rect 13726 9016 13782 9072
rect 13634 8200 13690 8256
rect 14002 9832 14058 9888
rect 14002 8200 14058 8256
rect 13358 5752 13414 5808
rect 12990 3168 13046 3224
rect 13450 4800 13506 4856
rect 13818 7692 13820 7712
rect 13820 7692 13872 7712
rect 13872 7692 13874 7712
rect 13818 7656 13874 7692
rect 13818 7112 13874 7168
rect 13726 4800 13782 4856
rect 13726 4392 13782 4448
rect 14002 6296 14058 6352
rect 14002 5480 14058 5536
rect 14370 15816 14426 15872
rect 14462 13368 14518 13424
rect 14462 12416 14518 12472
rect 14646 15272 14702 15328
rect 14646 14456 14702 14512
rect 14186 10512 14242 10568
rect 14186 10240 14242 10296
rect 14554 12144 14610 12200
rect 14554 11328 14610 11384
rect 14462 10920 14518 10976
rect 14462 10684 14464 10704
rect 14464 10684 14516 10704
rect 14516 10684 14518 10704
rect 14462 10648 14518 10684
rect 14462 10376 14518 10432
rect 14370 9016 14426 9072
rect 15198 26288 15254 26344
rect 15198 26152 15254 26208
rect 15658 29164 15714 29200
rect 15658 29144 15660 29164
rect 15660 29144 15712 29164
rect 15712 29144 15714 29164
rect 15750 29008 15806 29064
rect 15658 26560 15714 26616
rect 15106 23976 15162 24032
rect 15014 20848 15070 20904
rect 14830 19488 14886 19544
rect 14738 12416 14794 12472
rect 14186 8336 14242 8392
rect 14186 7112 14242 7168
rect 14462 7656 14518 7712
rect 15014 15272 15070 15328
rect 15290 23432 15346 23488
rect 15198 21664 15254 21720
rect 15474 25608 15530 25664
rect 15842 25336 15898 25392
rect 15566 22752 15622 22808
rect 15842 24248 15898 24304
rect 16026 23704 16082 23760
rect 15658 22344 15714 22400
rect 15382 21684 15438 21720
rect 15382 21664 15384 21684
rect 15384 21664 15436 21684
rect 15436 21664 15438 21684
rect 15382 20304 15438 20360
rect 15198 19488 15254 19544
rect 15566 20712 15622 20768
rect 15474 18536 15530 18592
rect 15198 16768 15254 16824
rect 15474 16768 15530 16824
rect 15382 15816 15438 15872
rect 15198 13096 15254 13152
rect 14830 10512 14886 10568
rect 15474 13096 15530 13152
rect 15474 11600 15530 11656
rect 15106 10240 15162 10296
rect 14646 6296 14702 6352
rect 14186 4800 14242 4856
rect 14094 3984 14150 4040
rect 14278 3984 14334 4040
rect 14462 4004 14518 4040
rect 14646 4820 14702 4856
rect 14646 4800 14648 4820
rect 14648 4800 14700 4820
rect 14700 4800 14702 4820
rect 14462 3984 14464 4004
rect 14464 3984 14516 4004
rect 14516 3984 14518 4004
rect 14094 3712 14150 3768
rect 14830 7112 14886 7168
rect 15198 8336 15254 8392
rect 15198 7112 15254 7168
rect 15198 6840 15254 6896
rect 15198 6568 15254 6624
rect 15842 14592 15898 14648
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 17498 29416 17554 29472
rect 16026 20848 16082 20904
rect 16118 20712 16174 20768
rect 16026 19896 16082 19952
rect 16118 18536 16174 18592
rect 16118 17720 16174 17776
rect 16118 14592 16174 14648
rect 16578 26968 16634 27024
rect 16394 23840 16450 23896
rect 16762 26424 16818 26480
rect 17406 28328 17462 28384
rect 16946 27648 17002 27704
rect 16854 25472 16910 25528
rect 16670 22752 16726 22808
rect 16578 22616 16634 22672
rect 16486 21664 16542 21720
rect 16394 19760 16450 19816
rect 16302 19488 16358 19544
rect 17590 26832 17646 26888
rect 17222 23604 17224 23624
rect 17224 23604 17276 23624
rect 17276 23604 17278 23624
rect 17222 23568 17278 23604
rect 16670 20712 16726 20768
rect 16670 19352 16726 19408
rect 16946 19488 17002 19544
rect 16394 18264 16450 18320
rect 16578 17720 16634 17776
rect 16486 15680 16542 15736
rect 16302 14728 16358 14784
rect 16486 14728 16542 14784
rect 16210 14456 16266 14512
rect 16486 14456 16542 14512
rect 16762 15544 16818 15600
rect 16670 14728 16726 14784
rect 16394 14184 16450 14240
rect 16486 13912 16542 13968
rect 16118 13232 16174 13288
rect 16394 13640 16450 13696
rect 17130 21392 17186 21448
rect 17682 26288 17738 26344
rect 17682 25744 17738 25800
rect 17866 23840 17922 23896
rect 17958 23588 18014 23624
rect 17958 23568 17960 23588
rect 17960 23568 18012 23588
rect 18012 23568 18014 23588
rect 17314 19352 17370 19408
rect 17130 17720 17186 17776
rect 17958 22480 18014 22536
rect 17958 22072 18014 22128
rect 17866 21664 17922 21720
rect 17590 19352 17646 19408
rect 17130 17448 17186 17504
rect 16946 16788 17002 16824
rect 16946 16768 16948 16788
rect 16948 16768 17000 16788
rect 17000 16768 17002 16788
rect 17038 16088 17094 16144
rect 17038 15680 17094 15736
rect 17314 15544 17370 15600
rect 17314 15000 17370 15056
rect 17590 16088 17646 16144
rect 18050 21800 18106 21856
rect 18234 26016 18290 26072
rect 18142 20984 18198 21040
rect 17866 20712 17922 20768
rect 17958 20576 18014 20632
rect 17958 18672 18014 18728
rect 18234 19624 18290 19680
rect 18142 19372 18198 19408
rect 18142 19352 18144 19372
rect 18144 19352 18196 19372
rect 18196 19352 18198 19372
rect 17958 18300 17960 18320
rect 17960 18300 18012 18320
rect 18012 18300 18014 18320
rect 17958 18264 18014 18300
rect 17774 17992 17830 18048
rect 17958 17484 17960 17504
rect 17960 17484 18012 17504
rect 18012 17484 18014 17504
rect 17958 17448 18014 17484
rect 17958 17076 17960 17096
rect 17960 17076 18012 17096
rect 18012 17076 18014 17096
rect 17958 17040 18014 17076
rect 17774 15408 17830 15464
rect 18142 15680 18198 15736
rect 16946 13504 17002 13560
rect 16854 13232 16910 13288
rect 15934 12416 15990 12472
rect 15750 10376 15806 10432
rect 15658 9696 15714 9752
rect 15566 7520 15622 7576
rect 15474 6976 15530 7032
rect 15474 6568 15530 6624
rect 15382 5616 15438 5672
rect 15198 5480 15254 5536
rect 15198 5364 15254 5400
rect 15198 5344 15200 5364
rect 15200 5344 15252 5364
rect 15252 5344 15254 5364
rect 15198 4800 15254 4856
rect 15290 4684 15346 4720
rect 15290 4664 15292 4684
rect 15292 4664 15344 4684
rect 15344 4664 15346 4684
rect 15106 4392 15162 4448
rect 15658 6976 15714 7032
rect 15658 6296 15714 6352
rect 15658 5480 15714 5536
rect 15842 9832 15898 9888
rect 15842 4392 15898 4448
rect 15842 3984 15898 4040
rect 15566 3848 15622 3904
rect 15014 2080 15070 2136
rect 16026 9696 16082 9752
rect 16210 11600 16266 11656
rect 16210 10104 16266 10160
rect 16302 9988 16358 10024
rect 16302 9968 16304 9988
rect 16304 9968 16356 9988
rect 16356 9968 16358 9988
rect 16670 12960 16726 13016
rect 16670 12688 16726 12744
rect 16762 12416 16818 12472
rect 17222 13504 17278 13560
rect 16670 10920 16726 10976
rect 16210 9288 16266 9344
rect 16026 7656 16082 7712
rect 16210 8608 16266 8664
rect 16486 9016 16542 9072
rect 16486 8628 16542 8664
rect 16486 8608 16488 8628
rect 16488 8608 16540 8628
rect 16540 8608 16542 8628
rect 16762 10104 16818 10160
rect 16762 9968 16818 10024
rect 16762 9696 16818 9752
rect 16946 9016 17002 9072
rect 16394 8372 16396 8392
rect 16396 8372 16448 8392
rect 16448 8372 16450 8392
rect 16394 8336 16450 8372
rect 16118 5480 16174 5536
rect 17590 12688 17646 12744
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19154 28484 19210 28520
rect 19154 28464 19156 28484
rect 19156 28464 19208 28484
rect 19208 28464 19210 28484
rect 18970 28192 19026 28248
rect 18694 24556 18696 24576
rect 18696 24556 18748 24576
rect 18748 24556 18750 24576
rect 18694 24520 18750 24556
rect 18694 22344 18750 22400
rect 19522 28872 19578 28928
rect 19798 28464 19854 28520
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20074 28092 20076 28112
rect 20076 28092 20128 28112
rect 20128 28092 20130 28112
rect 20074 28056 20130 28092
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19430 26832 19486 26888
rect 19338 25764 19394 25800
rect 19338 25744 19340 25764
rect 19340 25744 19392 25764
rect 19392 25744 19394 25764
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19154 23296 19210 23352
rect 18878 22208 18934 22264
rect 18786 22072 18842 22128
rect 18510 21392 18566 21448
rect 18510 20576 18566 20632
rect 18418 19896 18474 19952
rect 18510 17992 18566 18048
rect 18326 17176 18382 17232
rect 18326 14592 18382 14648
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19706 24384 19762 24440
rect 19430 23976 19486 24032
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20626 30368 20682 30424
rect 20534 28056 20590 28112
rect 20166 24692 20168 24712
rect 20168 24692 20220 24712
rect 20220 24692 20222 24712
rect 20166 24656 20222 24692
rect 20350 22752 20406 22808
rect 19522 22480 19578 22536
rect 20074 22228 20130 22264
rect 20074 22208 20076 22228
rect 20076 22208 20128 22228
rect 20128 22208 20130 22228
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19430 21664 19486 21720
rect 19062 21392 19118 21448
rect 19154 20748 19156 20768
rect 19156 20748 19208 20768
rect 19208 20748 19210 20768
rect 19154 20712 19210 20748
rect 19522 21256 19578 21312
rect 19430 20712 19486 20768
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20166 20712 20222 20768
rect 19430 20596 19486 20632
rect 19430 20576 19432 20596
rect 19432 20576 19484 20596
rect 19484 20576 19486 20596
rect 19982 20576 20038 20632
rect 20350 20712 20406 20768
rect 20718 22480 20774 22536
rect 19246 19760 19302 19816
rect 19706 19760 19762 19816
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19430 19488 19486 19544
rect 18694 19216 18750 19272
rect 18786 18944 18842 19000
rect 18510 16632 18566 16688
rect 18510 14184 18566 14240
rect 18510 13776 18566 13832
rect 18970 18708 18972 18728
rect 18972 18708 19024 18728
rect 19024 18708 19026 18728
rect 18970 18672 19026 18708
rect 19154 19216 19210 19272
rect 19154 19080 19210 19136
rect 19338 18944 19394 19000
rect 19154 18536 19210 18592
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20166 19760 20222 19816
rect 20166 18944 20222 19000
rect 20442 19896 20498 19952
rect 20626 20440 20682 20496
rect 21638 26288 21694 26344
rect 21270 22480 21326 22536
rect 21362 21256 21418 21312
rect 20442 19116 20444 19136
rect 20444 19116 20496 19136
rect 20496 19116 20498 19136
rect 20442 19080 20498 19116
rect 20350 18808 20406 18864
rect 20258 18672 20314 18728
rect 18878 16632 18934 16688
rect 19154 17176 19210 17232
rect 19982 17484 19984 17504
rect 19984 17484 20036 17504
rect 20036 17484 20038 17504
rect 19982 17448 20038 17484
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19982 17312 20038 17368
rect 19614 17176 19670 17232
rect 20166 17448 20222 17504
rect 19338 17040 19394 17096
rect 19338 16768 19394 16824
rect 19522 16768 19578 16824
rect 18878 16224 18934 16280
rect 19062 16224 19118 16280
rect 19062 15952 19118 16008
rect 19062 15680 19118 15736
rect 18694 13776 18750 13832
rect 17406 11056 17462 11112
rect 17682 10920 17738 10976
rect 17958 12688 18014 12744
rect 18326 12688 18382 12744
rect 18234 11636 18236 11656
rect 18236 11636 18288 11656
rect 18288 11636 18290 11656
rect 18234 11600 18290 11636
rect 18418 11600 18474 11656
rect 17222 9696 17278 9752
rect 16946 8744 17002 8800
rect 16762 8608 16818 8664
rect 17130 8744 17186 8800
rect 16578 6568 16634 6624
rect 16394 5616 16450 5672
rect 16486 5480 16542 5536
rect 16394 4120 16450 4176
rect 16854 8336 16910 8392
rect 17406 8744 17462 8800
rect 17314 8064 17370 8120
rect 17682 9560 17738 9616
rect 18050 10104 18106 10160
rect 18234 10920 18290 10976
rect 17038 7520 17094 7576
rect 16762 6568 16818 6624
rect 17314 7248 17370 7304
rect 16854 6296 16910 6352
rect 16762 5208 16818 5264
rect 16670 4684 16726 4720
rect 16670 4664 16672 4684
rect 16672 4664 16724 4684
rect 16724 4664 16726 4684
rect 16210 3576 16266 3632
rect 16394 3576 16450 3632
rect 16302 3168 16358 3224
rect 16578 3168 16634 3224
rect 15474 2216 15530 2272
rect 17038 5908 17094 5944
rect 17038 5888 17040 5908
rect 17040 5888 17092 5908
rect 17092 5888 17094 5908
rect 17038 4120 17094 4176
rect 16670 2760 16726 2816
rect 17498 6568 17554 6624
rect 17498 6296 17554 6352
rect 17498 5752 17554 5808
rect 17498 5344 17554 5400
rect 17498 4936 17554 4992
rect 17958 8336 18014 8392
rect 17774 8084 17830 8120
rect 17774 8064 17776 8084
rect 17776 8064 17828 8084
rect 17828 8064 17830 8084
rect 18234 9016 18290 9072
rect 17958 7112 18014 7168
rect 17866 6704 17922 6760
rect 20626 19216 20682 19272
rect 20902 18808 20958 18864
rect 21638 22072 21694 22128
rect 21362 20032 21418 20088
rect 20442 17448 20498 17504
rect 20350 17176 20406 17232
rect 19246 16224 19302 16280
rect 19154 15156 19210 15192
rect 19154 15136 19156 15156
rect 19156 15136 19208 15156
rect 19208 15136 19210 15156
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 20166 16632 20222 16688
rect 20718 17176 20774 17232
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19430 15136 19486 15192
rect 19982 15136 20038 15192
rect 20626 16632 20682 16688
rect 20166 15272 20222 15328
rect 19338 14220 19340 14240
rect 19340 14220 19392 14240
rect 19392 14220 19394 14240
rect 19338 14184 19394 14220
rect 20442 16360 20498 16416
rect 20534 16088 20590 16144
rect 21086 17176 21142 17232
rect 20994 16088 21050 16144
rect 20626 15408 20682 15464
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19430 14048 19486 14104
rect 18878 13096 18934 13152
rect 19062 13096 19118 13152
rect 18786 11092 18788 11112
rect 18788 11092 18840 11112
rect 18840 11092 18842 11112
rect 18786 11056 18842 11092
rect 19154 12008 19210 12064
rect 19062 11736 19118 11792
rect 19062 11600 19118 11656
rect 18878 9832 18934 9888
rect 19246 10920 19302 10976
rect 19338 9832 19394 9888
rect 18602 8744 18658 8800
rect 18602 8336 18658 8392
rect 18326 7656 18382 7712
rect 18510 7656 18566 7712
rect 18878 8336 18934 8392
rect 19062 8372 19064 8392
rect 19064 8372 19116 8392
rect 19116 8372 19118 8392
rect 19062 8336 19118 8372
rect 18878 8200 18934 8256
rect 18602 6976 18658 7032
rect 18418 6704 18474 6760
rect 17958 6432 18014 6488
rect 18050 5888 18106 5944
rect 17958 4800 18014 4856
rect 18234 5752 18290 5808
rect 18142 5072 18198 5128
rect 17498 1672 17554 1728
rect 18602 6568 18658 6624
rect 18786 6432 18842 6488
rect 18694 5344 18750 5400
rect 18786 3304 18842 3360
rect 19062 7792 19118 7848
rect 19062 6568 19118 6624
rect 19062 5480 19118 5536
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19982 12008 20038 12064
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19706 9016 19762 9072
rect 20350 14184 20406 14240
rect 20350 13640 20406 13696
rect 20350 12280 20406 12336
rect 20258 11328 20314 11384
rect 20626 13776 20682 13832
rect 20626 13232 20682 13288
rect 20166 9560 20222 9616
rect 20350 10920 20406 10976
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20442 9832 20498 9888
rect 20810 15444 20812 15464
rect 20812 15444 20864 15464
rect 20864 15444 20866 15464
rect 20810 15408 20866 15444
rect 20902 15272 20958 15328
rect 20902 14728 20958 14784
rect 20902 14456 20958 14512
rect 21086 14456 21142 14512
rect 21362 17448 21418 17504
rect 21362 17040 21418 17096
rect 21362 16768 21418 16824
rect 22098 28464 22154 28520
rect 25318 33088 25374 33144
rect 22006 26152 22062 26208
rect 22282 25744 22338 25800
rect 22466 25608 22522 25664
rect 21914 23432 21970 23488
rect 21914 23044 21970 23080
rect 21914 23024 21916 23044
rect 21916 23024 21968 23044
rect 21968 23024 21970 23044
rect 21822 22616 21878 22672
rect 22282 24656 22338 24712
rect 22466 23704 22522 23760
rect 21914 21664 21970 21720
rect 21822 20440 21878 20496
rect 21638 19624 21694 19680
rect 21638 18400 21694 18456
rect 21270 16088 21326 16144
rect 20902 13812 20904 13832
rect 20904 13812 20956 13832
rect 20956 13812 20958 13832
rect 20902 13776 20958 13812
rect 21086 13640 21142 13696
rect 20902 13232 20958 13288
rect 20626 12008 20682 12064
rect 20810 12280 20866 12336
rect 20902 12008 20958 12064
rect 20902 11736 20958 11792
rect 20718 11328 20774 11384
rect 20626 10376 20682 10432
rect 20626 9832 20682 9888
rect 20994 10376 21050 10432
rect 20810 10240 20866 10296
rect 20718 9172 20774 9208
rect 20718 9152 20720 9172
rect 20720 9152 20772 9172
rect 20772 9152 20774 9172
rect 19982 8200 20038 8256
rect 19430 7656 19486 7712
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19982 6976 20038 7032
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19614 6316 19670 6352
rect 19614 6296 19616 6316
rect 19616 6296 19668 6316
rect 19668 6296 19670 6316
rect 19798 6296 19854 6352
rect 19430 5752 19486 5808
rect 20258 6316 20314 6352
rect 20258 6296 20260 6316
rect 20260 6296 20312 6316
rect 20312 6296 20314 6316
rect 20902 9424 20958 9480
rect 21086 10104 21142 10160
rect 21086 9832 21142 9888
rect 20994 9288 21050 9344
rect 21178 9172 21234 9208
rect 21178 9152 21180 9172
rect 21180 9152 21232 9172
rect 21232 9152 21234 9172
rect 21086 8880 21142 8936
rect 20902 8744 20958 8800
rect 20718 8200 20774 8256
rect 20718 7656 20774 7712
rect 20626 6568 20682 6624
rect 19982 5752 20038 5808
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19982 5344 20038 5400
rect 19154 4392 19210 4448
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19154 3168 19210 3224
rect 18970 2760 19026 2816
rect 19062 2488 19118 2544
rect 19246 2488 19302 2544
rect 19522 3984 19578 4040
rect 19890 3984 19946 4040
rect 20258 3440 20314 3496
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19246 2080 19302 2136
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20810 6432 20866 6488
rect 21178 8064 21234 8120
rect 20994 7792 21050 7848
rect 21086 6704 21142 6760
rect 20810 5652 20812 5672
rect 20812 5652 20864 5672
rect 20864 5652 20866 5672
rect 20810 5616 20866 5652
rect 20718 5480 20774 5536
rect 20994 5752 21050 5808
rect 20902 5344 20958 5400
rect 20810 5208 20866 5264
rect 20718 4528 20774 4584
rect 20626 4120 20682 4176
rect 20626 3576 20682 3632
rect 20534 2352 20590 2408
rect 20258 1808 20314 1864
rect 21178 5772 21234 5808
rect 21178 5752 21180 5772
rect 21180 5752 21232 5772
rect 21232 5752 21234 5772
rect 21546 16088 21602 16144
rect 22190 21428 22192 21448
rect 22192 21428 22244 21448
rect 22244 21428 22246 21448
rect 22190 21392 22246 21428
rect 22742 22752 22798 22808
rect 23018 26152 23074 26208
rect 22650 21664 22706 21720
rect 22558 21256 22614 21312
rect 21914 18808 21970 18864
rect 22466 20476 22468 20496
rect 22468 20476 22520 20496
rect 22520 20476 22522 20496
rect 22466 20440 22522 20476
rect 22374 20304 22430 20360
rect 22558 20304 22614 20360
rect 22374 19896 22430 19952
rect 22558 17448 22614 17504
rect 22098 17312 22154 17368
rect 22282 17312 22338 17368
rect 21730 16768 21786 16824
rect 22098 16768 22154 16824
rect 22282 16768 22338 16824
rect 21546 15544 21602 15600
rect 21362 15000 21418 15056
rect 22190 16632 22246 16688
rect 21914 15036 21916 15056
rect 21916 15036 21968 15056
rect 21968 15036 21970 15056
rect 21914 15000 21970 15036
rect 21730 14592 21786 14648
rect 21546 14456 21602 14512
rect 22834 21528 22890 21584
rect 23018 21936 23074 21992
rect 23018 21664 23074 21720
rect 22926 20440 22982 20496
rect 22834 17856 22890 17912
rect 23018 17856 23074 17912
rect 22834 17448 22890 17504
rect 22926 16632 22982 16688
rect 22742 15580 22744 15600
rect 22744 15580 22796 15600
rect 22796 15580 22798 15600
rect 22742 15544 22798 15580
rect 23294 22480 23350 22536
rect 23202 22344 23258 22400
rect 23294 22072 23350 22128
rect 23202 21664 23258 21720
rect 23294 21392 23350 21448
rect 23570 23296 23626 23352
rect 23938 20576 23994 20632
rect 23570 18264 23626 18320
rect 23294 17040 23350 17096
rect 23110 15988 23112 16008
rect 23112 15988 23164 16008
rect 23164 15988 23166 16008
rect 23110 15952 23166 15988
rect 23110 15680 23166 15736
rect 22466 15408 22522 15464
rect 22282 14728 22338 14784
rect 22006 14184 22062 14240
rect 21822 14048 21878 14104
rect 22282 14068 22338 14104
rect 22282 14048 22284 14068
rect 22284 14048 22336 14068
rect 22336 14048 22338 14068
rect 21822 13640 21878 13696
rect 21362 11600 21418 11656
rect 21362 8064 21418 8120
rect 21362 6180 21418 6216
rect 21362 6160 21364 6180
rect 21364 6160 21416 6180
rect 21416 6160 21418 6180
rect 21362 4664 21418 4720
rect 21914 13096 21970 13152
rect 21730 12844 21786 12880
rect 21730 12824 21732 12844
rect 21732 12824 21784 12844
rect 21784 12824 21786 12844
rect 22098 13640 22154 13696
rect 21730 11600 21786 11656
rect 21546 9596 21548 9616
rect 21548 9596 21600 9616
rect 21600 9596 21602 9616
rect 21546 9560 21602 9596
rect 21546 9052 21548 9072
rect 21548 9052 21600 9072
rect 21600 9052 21602 9072
rect 21546 9016 21602 9052
rect 21546 8064 21602 8120
rect 21914 11756 21970 11792
rect 21914 11736 21916 11756
rect 21916 11736 21968 11756
rect 21968 11736 21970 11756
rect 22006 11464 22062 11520
rect 22374 13776 22430 13832
rect 22650 13640 22706 13696
rect 22374 12824 22430 12880
rect 22558 12824 22614 12880
rect 21914 9832 21970 9888
rect 22006 8880 22062 8936
rect 21914 8744 21970 8800
rect 21822 8336 21878 8392
rect 22006 8336 22062 8392
rect 22282 10376 22338 10432
rect 22190 8880 22246 8936
rect 22466 8880 22522 8936
rect 22742 12960 22798 13016
rect 22650 9424 22706 9480
rect 21730 7248 21786 7304
rect 22098 7928 22154 7984
rect 21914 7792 21970 7848
rect 22098 6976 22154 7032
rect 22006 6840 22062 6896
rect 21362 3712 21418 3768
rect 22282 7248 22338 7304
rect 22282 6452 22338 6488
rect 22282 6432 22284 6452
rect 22284 6432 22336 6452
rect 22336 6432 22338 6452
rect 22466 7928 22522 7984
rect 22926 12960 22982 13016
rect 23202 15136 23258 15192
rect 23294 14456 23350 14512
rect 23110 13096 23166 13152
rect 23018 12844 23074 12880
rect 23018 12824 23020 12844
rect 23020 12824 23072 12844
rect 23072 12824 23074 12844
rect 23018 12416 23074 12472
rect 22926 11736 22982 11792
rect 23202 12008 23258 12064
rect 24122 20984 24178 21040
rect 24122 20460 24178 20496
rect 24122 20440 24124 20460
rect 24124 20440 24176 20460
rect 24176 20440 24178 20460
rect 24306 20304 24362 20360
rect 23846 18536 23902 18592
rect 23846 17720 23902 17776
rect 24122 16224 24178 16280
rect 23938 12144 23994 12200
rect 23662 10648 23718 10704
rect 22834 7928 22890 7984
rect 22650 7384 22706 7440
rect 22374 6160 22430 6216
rect 22098 4820 22154 4856
rect 22098 4800 22100 4820
rect 22100 4800 22152 4820
rect 22152 4800 22154 4820
rect 21730 3984 21786 4040
rect 22006 3984 22062 4040
rect 21822 2760 21878 2816
rect 22282 4972 22284 4992
rect 22284 4972 22336 4992
rect 22336 4972 22338 4992
rect 22282 4936 22338 4972
rect 22466 5752 22522 5808
rect 22282 1944 22338 2000
rect 22926 6296 22982 6352
rect 23110 5072 23166 5128
rect 23386 8608 23442 8664
rect 23570 8608 23626 8664
rect 23938 11056 23994 11112
rect 23754 10240 23810 10296
rect 23386 6860 23442 6896
rect 23386 6840 23388 6860
rect 23388 6840 23440 6860
rect 23440 6840 23442 6860
rect 23294 2624 23350 2680
rect 23294 2488 23350 2544
rect 23754 8200 23810 8256
rect 23570 6568 23626 6624
rect 24030 5888 24086 5944
rect 24306 18808 24362 18864
rect 24306 7656 24362 7712
rect 24490 24112 24546 24168
rect 24950 22344 25006 22400
rect 24858 22208 24914 22264
rect 24950 20712 25006 20768
rect 25042 19352 25098 19408
rect 25226 26832 25282 26888
rect 24674 18536 24730 18592
rect 24950 17448 25006 17504
rect 24858 17312 24914 17368
rect 24950 17040 25006 17096
rect 25042 16768 25098 16824
rect 24858 15680 24914 15736
rect 24674 13252 24730 13288
rect 24674 13232 24676 13252
rect 24676 13232 24728 13252
rect 24728 13232 24730 13252
rect 25042 14184 25098 14240
rect 24582 11872 24638 11928
rect 24582 11464 24638 11520
rect 25410 19624 25466 19680
rect 25962 20868 26018 20904
rect 25962 20848 25964 20868
rect 25964 20848 26016 20868
rect 26016 20848 26018 20868
rect 25962 20340 25964 20360
rect 25964 20340 26016 20360
rect 26016 20340 26018 20360
rect 25962 20304 26018 20340
rect 25410 17720 25466 17776
rect 25318 14728 25374 14784
rect 25134 12164 25190 12200
rect 25134 12144 25136 12164
rect 25136 12144 25188 12164
rect 25188 12144 25190 12164
rect 25134 11736 25190 11792
rect 24582 9968 24638 10024
rect 24674 9152 24730 9208
rect 24582 8608 24638 8664
rect 23938 3884 23940 3904
rect 23940 3884 23992 3904
rect 23992 3884 23994 3904
rect 23938 3848 23994 3884
rect 24674 7112 24730 7168
rect 24674 6860 24730 6896
rect 24674 6840 24676 6860
rect 24676 6840 24728 6860
rect 24728 6840 24730 6860
rect 24030 3476 24032 3496
rect 24032 3476 24084 3496
rect 24084 3476 24086 3496
rect 24030 3440 24086 3476
rect 23386 1264 23442 1320
rect 24858 8064 24914 8120
rect 25042 9016 25098 9072
rect 24858 7540 24914 7576
rect 24858 7520 24860 7540
rect 24860 7520 24912 7540
rect 24912 7520 24914 7540
rect 24858 5480 24914 5536
rect 25042 2896 25098 2952
rect 25502 15544 25558 15600
rect 25318 11872 25374 11928
rect 25686 18672 25742 18728
rect 25686 16632 25742 16688
rect 25594 11328 25650 11384
rect 25686 10104 25742 10160
rect 26054 20032 26110 20088
rect 26054 19352 26110 19408
rect 25870 14456 25926 14512
rect 26422 23160 26478 23216
rect 26238 19760 26294 19816
rect 26146 18944 26202 19000
rect 26330 18572 26332 18592
rect 26332 18572 26384 18592
rect 26384 18572 26386 18592
rect 26330 18536 26386 18572
rect 26054 14864 26110 14920
rect 25962 14320 26018 14376
rect 25502 8492 25558 8528
rect 25502 8472 25504 8492
rect 25504 8472 25556 8492
rect 25556 8472 25558 8492
rect 25686 8336 25742 8392
rect 26054 12008 26110 12064
rect 26146 10804 26202 10840
rect 26146 10784 26148 10804
rect 26148 10784 26200 10804
rect 26200 10784 26202 10804
rect 26146 8744 26202 8800
rect 27066 23024 27122 23080
rect 26882 21972 26884 21992
rect 26884 21972 26936 21992
rect 26936 21972 26938 21992
rect 26882 21936 26938 21972
rect 27066 19488 27122 19544
rect 26790 19216 26846 19272
rect 26606 14592 26662 14648
rect 26422 14184 26478 14240
rect 26606 14184 26662 14240
rect 26606 14068 26662 14104
rect 26606 14048 26608 14068
rect 26608 14048 26660 14068
rect 26660 14048 26662 14068
rect 26606 13504 26662 13560
rect 26514 12688 26570 12744
rect 26882 16088 26938 16144
rect 27066 19080 27122 19136
rect 27066 18264 27122 18320
rect 27802 22072 27858 22128
rect 27342 18400 27398 18456
rect 27250 18148 27306 18184
rect 27250 18128 27252 18148
rect 27252 18128 27304 18148
rect 27304 18128 27306 18148
rect 27250 17856 27306 17912
rect 27066 16768 27122 16824
rect 26974 15952 27030 16008
rect 26790 10920 26846 10976
rect 27894 20476 27896 20496
rect 27896 20476 27948 20496
rect 27948 20476 27950 20496
rect 27894 20440 27950 20476
rect 27710 19932 27712 19952
rect 27712 19932 27764 19952
rect 27764 19932 27766 19952
rect 27710 19896 27766 19932
rect 27618 19388 27620 19408
rect 27620 19388 27672 19408
rect 27672 19388 27674 19408
rect 27618 19352 27674 19388
rect 27526 17076 27528 17096
rect 27528 17076 27580 17096
rect 27580 17076 27582 17096
rect 27526 17040 27582 17076
rect 27710 17176 27766 17232
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 29182 22380 29184 22400
rect 29184 22380 29236 22400
rect 29236 22380 29238 22400
rect 29182 22344 29238 22380
rect 29090 21936 29146 21992
rect 28630 21256 28686 21312
rect 27434 16088 27490 16144
rect 27158 15816 27214 15872
rect 27066 14764 27068 14784
rect 27068 14764 27120 14784
rect 27120 14764 27122 14784
rect 27066 14728 27122 14764
rect 27158 14356 27160 14376
rect 27160 14356 27212 14376
rect 27212 14356 27214 14376
rect 27158 14320 27214 14356
rect 27342 15020 27398 15056
rect 27342 15000 27344 15020
rect 27344 15000 27396 15020
rect 27396 15000 27398 15020
rect 27250 13776 27306 13832
rect 27618 13776 27674 13832
rect 27342 12688 27398 12744
rect 26882 10512 26938 10568
rect 27342 9832 27398 9888
rect 26054 3304 26110 3360
rect 25410 3052 25466 3088
rect 25410 3032 25412 3052
rect 25412 3032 25464 3052
rect 25464 3032 25466 3052
rect 28446 16904 28502 16960
rect 27986 13368 28042 13424
rect 28170 14340 28226 14376
rect 28170 14320 28172 14340
rect 28172 14320 28224 14340
rect 28224 14320 28226 14340
rect 28262 12144 28318 12200
rect 28814 17992 28870 18048
rect 28722 17584 28778 17640
rect 29182 18128 29238 18184
rect 29274 17992 29330 18048
rect 29182 17856 29238 17912
rect 28630 16360 28686 16416
rect 29090 16532 29092 16552
rect 29092 16532 29144 16552
rect 29144 16532 29146 16552
rect 29090 16496 29146 16532
rect 28814 14456 28870 14512
rect 28906 12552 28962 12608
rect 29090 15136 29146 15192
rect 29090 13912 29146 13968
rect 29458 18148 29514 18184
rect 29458 18128 29460 18148
rect 29460 18128 29512 18148
rect 29512 18128 29514 18148
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 29274 11192 29330 11248
rect 31298 18128 31354 18184
rect 30838 17992 30894 18048
rect 30378 13912 30434 13968
rect 30378 12980 30434 13016
rect 30378 12960 30380 12980
rect 30380 12960 30432 12980
rect 30432 12960 30434 12980
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 36818 38800 36874 38856
rect 37462 36760 37518 36816
rect 37186 34040 37242 34096
rect 37186 31320 37242 31376
rect 37186 28600 37242 28656
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 30378 2352 30434 2408
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37462 32000 37518 32056
rect 37462 27240 37518 27296
rect 38290 38120 38346 38176
rect 37646 25220 37702 25256
rect 37646 25200 37648 25220
rect 37648 25200 37700 25220
rect 37700 25200 37702 25220
rect 37462 23840 37518 23896
rect 37462 17076 37464 17096
rect 37464 17076 37516 17096
rect 37516 17076 37518 17096
rect 37462 17040 37518 17076
rect 37462 11636 37464 11656
rect 37464 11636 37516 11656
rect 37516 11636 37518 11656
rect 37462 11600 37518 11636
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 37186 9560 37242 9616
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36910 2760 36966 2816
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37186 2080 37242 2136
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38106 33360 38162 33416
rect 38106 30660 38162 30696
rect 38106 30640 38108 30660
rect 38108 30640 38160 30660
rect 38160 30640 38162 30660
rect 38290 29280 38346 29336
rect 38290 26560 38346 26616
rect 38198 25880 38254 25936
rect 38198 24520 38254 24576
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38290 21800 38346 21856
rect 38198 21684 38254 21720
rect 38198 21664 38200 21684
rect 38200 21664 38252 21684
rect 38252 21664 38254 21684
rect 38106 21120 38162 21176
rect 38290 19796 38292 19816
rect 38292 19796 38344 19816
rect 38344 19796 38346 19816
rect 38290 19760 38346 19796
rect 38290 18400 38346 18456
rect 38106 16360 38162 16416
rect 38198 15000 38254 15056
rect 38198 14320 38254 14376
rect 38290 13640 38346 13696
rect 38198 12280 38254 12336
rect 38106 10240 38162 10296
rect 38198 8880 38254 8936
rect 38290 7520 38346 7576
rect 38106 6840 38162 6896
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 38198 4800 38254 4856
rect 38198 4120 38254 4176
rect 38290 720 38346 776
rect 37278 40 37334 96
<< metal3 >>
rect 200 39538 800 39568
rect 3049 39538 3115 39541
rect 200 39536 3115 39538
rect 200 39480 3054 39536
rect 3110 39480 3115 39536
rect 200 39478 3115 39480
rect 200 39448 800 39478
rect 3049 39475 3115 39478
rect 200 38858 800 38888
rect 2865 38858 2931 38861
rect 200 38856 2931 38858
rect 200 38800 2870 38856
rect 2926 38800 2931 38856
rect 200 38798 2931 38800
rect 200 38768 800 38798
rect 2865 38795 2931 38798
rect 36813 38858 36879 38861
rect 39200 38858 39800 38888
rect 36813 38856 39800 38858
rect 36813 38800 36818 38856
rect 36874 38800 39800 38856
rect 36813 38798 39800 38800
rect 36813 38795 36879 38798
rect 39200 38768 39800 38798
rect 38285 38178 38351 38181
rect 39200 38178 39800 38208
rect 38285 38176 39800 38178
rect 38285 38120 38290 38176
rect 38346 38120 39800 38176
rect 38285 38118 39800 38120
rect 38285 38115 38351 38118
rect 39200 38088 39800 38118
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 3141 37498 3207 37501
rect 200 37496 3207 37498
rect 200 37440 3146 37496
rect 3202 37440 3207 37496
rect 200 37438 3207 37440
rect 200 37408 800 37438
rect 3141 37435 3207 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 200 36818 800 36848
rect 1761 36818 1827 36821
rect 200 36816 1827 36818
rect 200 36760 1766 36816
rect 1822 36760 1827 36816
rect 200 36758 1827 36760
rect 200 36728 800 36758
rect 1761 36755 1827 36758
rect 37457 36818 37523 36821
rect 39200 36818 39800 36848
rect 37457 36816 39800 36818
rect 37457 36760 37462 36816
rect 37518 36760 39800 36816
rect 37457 36758 39800 36760
rect 37457 36755 37523 36758
rect 39200 36728 39800 36758
rect 8518 36484 8524 36548
rect 8588 36546 8594 36548
rect 9121 36546 9187 36549
rect 8588 36544 9187 36546
rect 8588 36488 9126 36544
rect 9182 36488 9187 36544
rect 8588 36486 9187 36488
rect 8588 36484 8594 36486
rect 9121 36483 9187 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 200 35458 800 35488
rect 1577 35458 1643 35461
rect 200 35456 1643 35458
rect 200 35400 1582 35456
rect 1638 35400 1643 35456
rect 200 35398 1643 35400
rect 200 35368 800 35398
rect 1577 35395 1643 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 200 34688 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 37181 34098 37247 34101
rect 39200 34098 39800 34128
rect 37181 34096 39800 34098
rect 37181 34040 37186 34096
rect 37242 34040 39800 34096
rect 37181 34038 39800 34040
rect 37181 34035 37247 34038
rect 39200 34008 39800 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 38101 33418 38167 33421
rect 39200 33418 39800 33448
rect 38101 33416 39800 33418
rect 38101 33360 38106 33416
rect 38162 33360 39800 33416
rect 38101 33358 39800 33360
rect 38101 33355 38167 33358
rect 39200 33328 39800 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 25313 33146 25379 33149
rect 27286 33146 27292 33148
rect 25313 33144 27292 33146
rect 25313 33088 25318 33144
rect 25374 33088 27292 33144
rect 25313 33086 27292 33088
rect 25313 33083 25379 33086
rect 27286 33084 27292 33086
rect 27356 33084 27362 33148
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 37457 32058 37523 32061
rect 39200 32058 39800 32088
rect 37457 32056 39800 32058
rect 37457 32000 37462 32056
rect 37518 32000 39800 32056
rect 37457 31998 39800 32000
rect 37457 31995 37523 31998
rect 39200 31968 39800 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 37181 31378 37247 31381
rect 39200 31378 39800 31408
rect 37181 31376 39800 31378
rect 37181 31320 37186 31376
rect 37242 31320 39800 31376
rect 37181 31318 39800 31320
rect 37181 31315 37247 31318
rect 39200 31288 39800 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 38101 30698 38167 30701
rect 39200 30698 39800 30728
rect 38101 30696 39800 30698
rect 38101 30640 38106 30696
rect 38162 30640 39800 30696
rect 38101 30638 39800 30640
rect 38101 30635 38167 30638
rect 39200 30608 39800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 1158 30364 1164 30428
rect 1228 30426 1234 30428
rect 1393 30426 1459 30429
rect 1228 30424 1459 30426
rect 1228 30368 1398 30424
rect 1454 30368 1459 30424
rect 1228 30366 1459 30368
rect 1228 30364 1234 30366
rect 1393 30363 1459 30366
rect 2037 30428 2103 30429
rect 2037 30424 2084 30428
rect 2148 30426 2154 30428
rect 4429 30426 4495 30429
rect 4838 30426 4844 30428
rect 2037 30368 2042 30424
rect 2037 30364 2084 30368
rect 2148 30366 2194 30426
rect 4429 30424 4844 30426
rect 4429 30368 4434 30424
rect 4490 30368 4844 30424
rect 4429 30366 4844 30368
rect 2148 30364 2154 30366
rect 2037 30363 2103 30364
rect 4429 30363 4495 30366
rect 4838 30364 4844 30366
rect 4908 30364 4914 30428
rect 5165 30426 5231 30429
rect 5390 30426 5396 30428
rect 5165 30424 5396 30426
rect 5165 30368 5170 30424
rect 5226 30368 5396 30424
rect 5165 30366 5396 30368
rect 5165 30363 5231 30366
rect 5390 30364 5396 30366
rect 5460 30364 5466 30428
rect 12065 30426 12131 30429
rect 12750 30426 12756 30428
rect 12065 30424 12756 30426
rect 12065 30368 12070 30424
rect 12126 30368 12756 30424
rect 12065 30366 12756 30368
rect 12065 30363 12131 30366
rect 12750 30364 12756 30366
rect 12820 30364 12826 30428
rect 20621 30426 20687 30429
rect 22686 30426 22692 30428
rect 20621 30424 22692 30426
rect 20621 30368 20626 30424
rect 20682 30368 22692 30424
rect 20621 30366 22692 30368
rect 20621 30363 20687 30366
rect 22686 30364 22692 30366
rect 22756 30364 22762 30428
rect 11881 30290 11947 30293
rect 21582 30290 21588 30292
rect 11881 30288 21588 30290
rect 11881 30232 11886 30288
rect 11942 30232 21588 30288
rect 11881 30230 21588 30232
rect 11881 30227 11947 30230
rect 21582 30228 21588 30230
rect 21652 30228 21658 30292
rect 8845 30154 8911 30157
rect 12249 30154 12315 30157
rect 16297 30156 16363 30157
rect 8845 30152 12315 30154
rect 8845 30096 8850 30152
rect 8906 30096 12254 30152
rect 12310 30096 12315 30152
rect 8845 30094 12315 30096
rect 8845 30091 8911 30094
rect 12249 30091 12315 30094
rect 16246 30092 16252 30156
rect 16316 30154 16363 30156
rect 16316 30152 16408 30154
rect 16358 30096 16408 30152
rect 16316 30094 16408 30096
rect 16316 30092 16363 30094
rect 16297 30091 16363 30092
rect 200 30018 800 30048
rect 3693 30018 3759 30021
rect 200 30016 3759 30018
rect 200 29960 3698 30016
rect 3754 29960 3759 30016
rect 200 29958 3759 29960
rect 200 29928 800 29958
rect 3693 29955 3759 29958
rect 9857 30018 9923 30021
rect 10593 30018 10659 30021
rect 9857 30016 10659 30018
rect 9857 29960 9862 30016
rect 9918 29960 10598 30016
rect 10654 29960 10659 30016
rect 9857 29958 10659 29960
rect 9857 29955 9923 29958
rect 10593 29955 10659 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 10593 29882 10659 29885
rect 10777 29882 10843 29885
rect 10593 29880 10843 29882
rect 10593 29824 10598 29880
rect 10654 29824 10782 29880
rect 10838 29824 10843 29880
rect 10593 29822 10843 29824
rect 10593 29819 10659 29822
rect 10777 29819 10843 29822
rect 9949 29746 10015 29749
rect 15009 29746 15075 29749
rect 9949 29744 15075 29746
rect 9949 29688 9954 29744
rect 10010 29688 15014 29744
rect 15070 29688 15075 29744
rect 9949 29686 15075 29688
rect 9949 29683 10015 29686
rect 15009 29683 15075 29686
rect 9765 29610 9831 29613
rect 10777 29610 10843 29613
rect 9765 29608 10843 29610
rect 9765 29552 9770 29608
rect 9826 29552 10782 29608
rect 10838 29552 10843 29608
rect 9765 29550 10843 29552
rect 9765 29547 9831 29550
rect 10777 29547 10843 29550
rect 10133 29474 10199 29477
rect 17493 29474 17559 29477
rect 10133 29472 17559 29474
rect 10133 29416 10138 29472
rect 10194 29416 17498 29472
rect 17554 29416 17559 29472
rect 10133 29414 17559 29416
rect 10133 29411 10199 29414
rect 17493 29411 17559 29414
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 3550 29276 3556 29340
rect 3620 29338 3626 29340
rect 8293 29338 8359 29341
rect 3620 29336 8359 29338
rect 3620 29280 8298 29336
rect 8354 29280 8359 29336
rect 3620 29278 8359 29280
rect 3620 29276 3626 29278
rect 8293 29275 8359 29278
rect 8661 29338 8727 29341
rect 8845 29338 8911 29341
rect 13077 29338 13143 29341
rect 8661 29336 13143 29338
rect 8661 29280 8666 29336
rect 8722 29280 8850 29336
rect 8906 29280 13082 29336
rect 13138 29280 13143 29336
rect 8661 29278 13143 29280
rect 8661 29275 8727 29278
rect 8845 29275 8911 29278
rect 13077 29275 13143 29278
rect 38285 29338 38351 29341
rect 39200 29338 39800 29368
rect 38285 29336 39800 29338
rect 38285 29280 38290 29336
rect 38346 29280 39800 29336
rect 38285 29278 39800 29280
rect 38285 29275 38351 29278
rect 39200 29248 39800 29278
rect 7005 29202 7071 29205
rect 7414 29202 7420 29204
rect 7005 29200 7420 29202
rect 7005 29144 7010 29200
rect 7066 29144 7420 29200
rect 7005 29142 7420 29144
rect 7005 29139 7071 29142
rect 7414 29140 7420 29142
rect 7484 29140 7490 29204
rect 12157 29202 12223 29205
rect 15653 29202 15719 29205
rect 12157 29200 15719 29202
rect 12157 29144 12162 29200
rect 12218 29144 15658 29200
rect 15714 29144 15719 29200
rect 12157 29142 15719 29144
rect 12157 29139 12223 29142
rect 15653 29139 15719 29142
rect 1894 29004 1900 29068
rect 1964 29066 1970 29068
rect 2589 29066 2655 29069
rect 1964 29064 2655 29066
rect 1964 29008 2594 29064
rect 2650 29008 2655 29064
rect 1964 29006 2655 29008
rect 1964 29004 1970 29006
rect 2589 29003 2655 29006
rect 6494 29004 6500 29068
rect 6564 29066 6570 29068
rect 7741 29066 7807 29069
rect 6564 29064 7807 29066
rect 6564 29008 7746 29064
rect 7802 29008 7807 29064
rect 6564 29006 7807 29008
rect 6564 29004 6570 29006
rect 7741 29003 7807 29006
rect 11646 29004 11652 29068
rect 11716 29066 11722 29068
rect 15745 29066 15811 29069
rect 11716 29064 15811 29066
rect 11716 29008 15750 29064
rect 15806 29008 15811 29064
rect 11716 29006 15811 29008
rect 11716 29004 11722 29006
rect 15745 29003 15811 29006
rect 19517 28930 19583 28933
rect 21950 28930 21956 28932
rect 19517 28928 21956 28930
rect 19517 28872 19522 28928
rect 19578 28872 21956 28928
rect 19517 28870 21956 28872
rect 19517 28867 19583 28870
rect 21950 28868 21956 28870
rect 22020 28868 22026 28932
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 10501 28794 10567 28797
rect 12525 28794 12591 28797
rect 10501 28792 12591 28794
rect 10501 28736 10506 28792
rect 10562 28736 12530 28792
rect 12586 28736 12591 28792
rect 10501 28734 12591 28736
rect 10501 28731 10567 28734
rect 12525 28731 12591 28734
rect 4613 28658 4679 28661
rect 5206 28658 5212 28660
rect 4613 28656 5212 28658
rect 4613 28600 4618 28656
rect 4674 28600 5212 28656
rect 4613 28598 5212 28600
rect 4613 28595 4679 28598
rect 5206 28596 5212 28598
rect 5276 28596 5282 28660
rect 37181 28658 37247 28661
rect 39200 28658 39800 28688
rect 37181 28656 39800 28658
rect 37181 28600 37186 28656
rect 37242 28600 39800 28656
rect 37181 28598 39800 28600
rect 37181 28595 37247 28598
rect 39200 28568 39800 28598
rect 2681 28522 2747 28525
rect 4654 28522 4660 28524
rect 2681 28520 4660 28522
rect 2681 28464 2686 28520
rect 2742 28464 4660 28520
rect 2681 28462 4660 28464
rect 2681 28459 2747 28462
rect 4654 28460 4660 28462
rect 4724 28460 4730 28524
rect 6678 28460 6684 28524
rect 6748 28522 6754 28524
rect 9397 28522 9463 28525
rect 6748 28520 9463 28522
rect 6748 28464 9402 28520
rect 9458 28464 9463 28520
rect 6748 28462 9463 28464
rect 6748 28460 6754 28462
rect 9397 28459 9463 28462
rect 10777 28522 10843 28525
rect 13353 28522 13419 28525
rect 19149 28522 19215 28525
rect 10777 28520 19215 28522
rect 10777 28464 10782 28520
rect 10838 28464 13358 28520
rect 13414 28464 19154 28520
rect 19210 28464 19215 28520
rect 10777 28462 19215 28464
rect 10777 28459 10843 28462
rect 13353 28459 13419 28462
rect 19149 28459 19215 28462
rect 19793 28522 19859 28525
rect 22093 28522 22159 28525
rect 19793 28520 22159 28522
rect 19793 28464 19798 28520
rect 19854 28464 22098 28520
rect 22154 28464 22159 28520
rect 19793 28462 22159 28464
rect 19793 28459 19859 28462
rect 22093 28459 22159 28462
rect 16982 28324 16988 28388
rect 17052 28386 17058 28388
rect 17401 28386 17467 28389
rect 17052 28384 17467 28386
rect 17052 28328 17406 28384
rect 17462 28328 17467 28384
rect 17052 28326 17467 28328
rect 17052 28324 17058 28326
rect 17401 28323 17467 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 9673 28250 9739 28253
rect 18965 28250 19031 28253
rect 9673 28248 19031 28250
rect 9673 28192 9678 28248
rect 9734 28192 18970 28248
rect 19026 28192 19031 28248
rect 9673 28190 19031 28192
rect 9673 28187 9739 28190
rect 18965 28187 19031 28190
rect 8477 28114 8543 28117
rect 9581 28114 9647 28117
rect 8477 28112 9647 28114
rect 8477 28056 8482 28112
rect 8538 28056 9586 28112
rect 9642 28056 9647 28112
rect 8477 28054 9647 28056
rect 8477 28051 8543 28054
rect 9581 28051 9647 28054
rect 12433 28114 12499 28117
rect 16246 28114 16252 28116
rect 12433 28112 16252 28114
rect 12433 28056 12438 28112
rect 12494 28056 16252 28112
rect 12433 28054 16252 28056
rect 12433 28051 12499 28054
rect 16246 28052 16252 28054
rect 16316 28052 16322 28116
rect 20069 28114 20135 28117
rect 20529 28114 20595 28117
rect 20069 28112 20595 28114
rect 20069 28056 20074 28112
rect 20130 28056 20534 28112
rect 20590 28056 20595 28112
rect 20069 28054 20595 28056
rect 20069 28051 20135 28054
rect 20529 28051 20595 28054
rect 200 27978 800 28008
rect 1761 27978 1827 27981
rect 200 27976 1827 27978
rect 200 27920 1766 27976
rect 1822 27920 1827 27976
rect 200 27918 1827 27920
rect 200 27888 800 27918
rect 1761 27915 1827 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 2814 27644 2820 27708
rect 2884 27706 2890 27708
rect 4061 27706 4127 27709
rect 2884 27704 4127 27706
rect 2884 27648 4066 27704
rect 4122 27648 4127 27704
rect 2884 27646 4127 27648
rect 2884 27644 2890 27646
rect 4061 27643 4127 27646
rect 7005 27708 7071 27709
rect 7005 27704 7052 27708
rect 7116 27706 7122 27708
rect 8753 27706 8819 27709
rect 9581 27706 9647 27709
rect 7005 27648 7010 27704
rect 7005 27644 7052 27648
rect 7116 27646 7162 27706
rect 8753 27704 9647 27706
rect 8753 27648 8758 27704
rect 8814 27648 9586 27704
rect 9642 27648 9647 27704
rect 8753 27646 9647 27648
rect 7116 27644 7122 27646
rect 7005 27643 7071 27644
rect 8753 27643 8819 27646
rect 9581 27643 9647 27646
rect 9806 27644 9812 27708
rect 9876 27706 9882 27708
rect 9949 27706 10015 27709
rect 9876 27704 10015 27706
rect 9876 27648 9954 27704
rect 10010 27648 10015 27704
rect 9876 27646 10015 27648
rect 9876 27644 9882 27646
rect 9949 27643 10015 27646
rect 10685 27708 10751 27709
rect 10685 27704 10732 27708
rect 10796 27706 10802 27708
rect 10685 27648 10690 27704
rect 10685 27644 10732 27648
rect 10796 27646 10842 27706
rect 10796 27644 10802 27646
rect 14958 27644 14964 27708
rect 15028 27706 15034 27708
rect 16941 27706 17007 27709
rect 15028 27704 17007 27706
rect 15028 27648 16946 27704
rect 17002 27648 17007 27704
rect 15028 27646 17007 27648
rect 15028 27644 15034 27646
rect 10685 27643 10751 27644
rect 16941 27643 17007 27646
rect 14549 27570 14615 27573
rect 14774 27570 14780 27572
rect 14549 27568 14780 27570
rect 14549 27512 14554 27568
rect 14610 27512 14780 27568
rect 14549 27510 14780 27512
rect 14549 27507 14615 27510
rect 14774 27508 14780 27510
rect 14844 27508 14850 27572
rect 8385 27436 8451 27437
rect 8334 27434 8340 27436
rect 8294 27374 8340 27434
rect 8404 27432 8451 27436
rect 8446 27376 8451 27432
rect 8334 27372 8340 27374
rect 8404 27372 8451 27376
rect 8385 27371 8451 27372
rect 8753 27434 8819 27437
rect 13077 27434 13143 27437
rect 8753 27432 13143 27434
rect 8753 27376 8758 27432
rect 8814 27376 13082 27432
rect 13138 27376 13143 27432
rect 8753 27374 13143 27376
rect 8753 27371 8819 27374
rect 13077 27371 13143 27374
rect 200 27298 800 27328
rect 1761 27298 1827 27301
rect 200 27296 1827 27298
rect 200 27240 1766 27296
rect 1822 27240 1827 27296
rect 200 27238 1827 27240
rect 200 27208 800 27238
rect 1761 27235 1827 27238
rect 37457 27298 37523 27301
rect 39200 27298 39800 27328
rect 37457 27296 39800 27298
rect 37457 27240 37462 27296
rect 37518 27240 39800 27296
rect 37457 27238 39800 27240
rect 37457 27235 37523 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 3734 27100 3740 27164
rect 3804 27162 3810 27164
rect 5073 27162 5139 27165
rect 3804 27160 5139 27162
rect 3804 27104 5078 27160
rect 5134 27104 5139 27160
rect 3804 27102 5139 27104
rect 3804 27100 3810 27102
rect 5073 27099 5139 27102
rect 4981 27028 5047 27029
rect 4981 27026 5028 27028
rect 4936 27024 5028 27026
rect 4936 26968 4986 27024
rect 4936 26966 5028 26968
rect 4981 26964 5028 26966
rect 5092 26964 5098 27028
rect 13445 27026 13511 27029
rect 16573 27026 16639 27029
rect 13445 27024 16639 27026
rect 13445 26968 13450 27024
rect 13506 26968 16578 27024
rect 16634 26968 16639 27024
rect 13445 26966 16639 26968
rect 4981 26963 5047 26964
rect 13445 26963 13511 26966
rect 16573 26963 16639 26966
rect 5574 26828 5580 26892
rect 5644 26890 5650 26892
rect 5717 26890 5783 26893
rect 5644 26888 5783 26890
rect 5644 26832 5722 26888
rect 5778 26832 5783 26888
rect 5644 26830 5783 26832
rect 5644 26828 5650 26830
rect 5717 26827 5783 26830
rect 6637 26890 6703 26893
rect 8201 26890 8267 26893
rect 10225 26890 10291 26893
rect 6637 26888 8034 26890
rect 6637 26832 6642 26888
rect 6698 26832 8034 26888
rect 6637 26830 8034 26832
rect 6637 26827 6703 26830
rect 5441 26754 5507 26757
rect 6862 26754 6868 26756
rect 5441 26752 6868 26754
rect 5441 26696 5446 26752
rect 5502 26696 6868 26752
rect 5441 26694 6868 26696
rect 5441 26691 5507 26694
rect 6862 26692 6868 26694
rect 6932 26692 6938 26756
rect 7974 26754 8034 26830
rect 8201 26888 10291 26890
rect 8201 26832 8206 26888
rect 8262 26832 10230 26888
rect 10286 26832 10291 26888
rect 8201 26830 10291 26832
rect 8201 26827 8267 26830
rect 10225 26827 10291 26830
rect 13629 26890 13695 26893
rect 16062 26890 16068 26892
rect 13629 26888 16068 26890
rect 13629 26832 13634 26888
rect 13690 26832 16068 26888
rect 13629 26830 16068 26832
rect 13629 26827 13695 26830
rect 16062 26828 16068 26830
rect 16132 26890 16138 26892
rect 17585 26890 17651 26893
rect 16132 26888 17651 26890
rect 16132 26832 17590 26888
rect 17646 26832 17651 26888
rect 16132 26830 17651 26832
rect 16132 26828 16138 26830
rect 17585 26827 17651 26830
rect 19425 26890 19491 26893
rect 25221 26890 25287 26893
rect 19425 26888 25287 26890
rect 19425 26832 19430 26888
rect 19486 26832 25226 26888
rect 25282 26832 25287 26888
rect 19425 26830 25287 26832
rect 19425 26827 19491 26830
rect 25221 26827 25287 26830
rect 8702 26754 8708 26756
rect 7974 26694 8708 26754
rect 8702 26692 8708 26694
rect 8772 26754 8778 26756
rect 8772 26694 9138 26754
rect 8772 26692 8778 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 9078 26618 9138 26694
rect 9254 26692 9260 26756
rect 9324 26754 9330 26756
rect 13537 26754 13603 26757
rect 9324 26752 13603 26754
rect 9324 26696 13542 26752
rect 13598 26696 13603 26752
rect 9324 26694 13603 26696
rect 9324 26692 9330 26694
rect 13537 26691 13603 26694
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 9489 26618 9555 26621
rect 9078 26616 9555 26618
rect 9078 26560 9494 26616
rect 9550 26560 9555 26616
rect 9078 26558 9555 26560
rect 9489 26555 9555 26558
rect 13670 26556 13676 26620
rect 13740 26618 13746 26620
rect 15653 26618 15719 26621
rect 13740 26616 15719 26618
rect 13740 26560 15658 26616
rect 15714 26560 15719 26616
rect 13740 26558 15719 26560
rect 13740 26556 13746 26558
rect 15653 26555 15719 26558
rect 38285 26618 38351 26621
rect 39200 26618 39800 26648
rect 38285 26616 39800 26618
rect 38285 26560 38290 26616
rect 38346 26560 39800 26616
rect 38285 26558 39800 26560
rect 38285 26555 38351 26558
rect 39200 26528 39800 26558
rect 10961 26484 11027 26485
rect 10910 26482 10916 26484
rect 10870 26422 10916 26482
rect 10980 26480 11027 26484
rect 11022 26424 11027 26480
rect 10910 26420 10916 26422
rect 10980 26420 11027 26424
rect 10961 26419 11027 26420
rect 11973 26482 12039 26485
rect 12801 26482 12867 26485
rect 16757 26482 16823 26485
rect 11973 26480 16823 26482
rect 11973 26424 11978 26480
rect 12034 26424 12806 26480
rect 12862 26424 16762 26480
rect 16818 26424 16823 26480
rect 11973 26422 16823 26424
rect 11973 26419 12039 26422
rect 12801 26419 12867 26422
rect 16757 26419 16823 26422
rect 3366 26284 3372 26348
rect 3436 26346 3442 26348
rect 4061 26346 4127 26349
rect 3436 26344 4127 26346
rect 3436 26288 4066 26344
rect 4122 26288 4127 26344
rect 3436 26286 4127 26288
rect 3436 26284 3442 26286
rect 4061 26283 4127 26286
rect 5993 26346 6059 26349
rect 6126 26346 6132 26348
rect 5993 26344 6132 26346
rect 5993 26288 5998 26344
rect 6054 26288 6132 26344
rect 5993 26286 6132 26288
rect 5993 26283 6059 26286
rect 6126 26284 6132 26286
rect 6196 26284 6202 26348
rect 7373 26346 7439 26349
rect 7598 26346 7604 26348
rect 7373 26344 7604 26346
rect 7373 26288 7378 26344
rect 7434 26288 7604 26344
rect 7373 26286 7604 26288
rect 7373 26283 7439 26286
rect 7598 26284 7604 26286
rect 7668 26284 7674 26348
rect 12566 26284 12572 26348
rect 12636 26346 12642 26348
rect 15193 26346 15259 26349
rect 12636 26344 15259 26346
rect 12636 26288 15198 26344
rect 15254 26288 15259 26344
rect 12636 26286 15259 26288
rect 12636 26284 12642 26286
rect 15193 26283 15259 26286
rect 17677 26348 17743 26349
rect 17677 26344 17724 26348
rect 17788 26346 17794 26348
rect 17677 26288 17682 26344
rect 17677 26284 17724 26288
rect 17788 26286 17834 26346
rect 17788 26284 17794 26286
rect 20110 26284 20116 26348
rect 20180 26346 20186 26348
rect 21633 26346 21699 26349
rect 20180 26344 21699 26346
rect 20180 26288 21638 26344
rect 21694 26288 21699 26344
rect 20180 26286 21699 26288
rect 20180 26284 20186 26286
rect 17677 26283 17743 26284
rect 21633 26283 21699 26286
rect 9765 26210 9831 26213
rect 15193 26210 15259 26213
rect 9765 26208 15259 26210
rect 9765 26152 9770 26208
rect 9826 26152 15198 26208
rect 15254 26152 15259 26208
rect 9765 26150 15259 26152
rect 9765 26147 9831 26150
rect 15193 26147 15259 26150
rect 22001 26210 22067 26213
rect 23013 26210 23079 26213
rect 22001 26208 23079 26210
rect 22001 26152 22006 26208
rect 22062 26152 23018 26208
rect 23074 26152 23079 26208
rect 22001 26150 23079 26152
rect 22001 26147 22067 26150
rect 23013 26147 23079 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 3049 26074 3115 26077
rect 1534 26072 3115 26074
rect 1534 26016 3054 26072
rect 3110 26016 3115 26072
rect 1534 26014 3115 26016
rect 200 25938 800 25968
rect 1534 25938 1594 26014
rect 3049 26011 3115 26014
rect 4705 26074 4771 26077
rect 6821 26074 6887 26077
rect 4705 26072 6887 26074
rect 4705 26016 4710 26072
rect 4766 26016 6826 26072
rect 6882 26016 6887 26072
rect 4705 26014 6887 26016
rect 4705 26011 4771 26014
rect 6821 26011 6887 26014
rect 11237 26074 11303 26077
rect 18229 26074 18295 26077
rect 11237 26072 18295 26074
rect 11237 26016 11242 26072
rect 11298 26016 18234 26072
rect 18290 26016 18295 26072
rect 11237 26014 18295 26016
rect 11237 26011 11303 26014
rect 18229 26011 18295 26014
rect 200 25878 1594 25938
rect 2313 25938 2379 25941
rect 23054 25938 23060 25940
rect 2313 25936 23060 25938
rect 2313 25880 2318 25936
rect 2374 25880 23060 25936
rect 2313 25878 23060 25880
rect 200 25848 800 25878
rect 2313 25875 2379 25878
rect 23054 25876 23060 25878
rect 23124 25876 23130 25940
rect 38193 25938 38259 25941
rect 39200 25938 39800 25968
rect 38193 25936 39800 25938
rect 38193 25880 38198 25936
rect 38254 25880 39800 25936
rect 38193 25878 39800 25880
rect 38193 25875 38259 25878
rect 39200 25848 39800 25878
rect 4061 25802 4127 25805
rect 6913 25802 6979 25805
rect 7281 25804 7347 25805
rect 4061 25800 6979 25802
rect 4061 25744 4066 25800
rect 4122 25744 6918 25800
rect 6974 25744 6979 25800
rect 4061 25742 6979 25744
rect 4061 25739 4127 25742
rect 6913 25739 6979 25742
rect 7230 25740 7236 25804
rect 7300 25802 7347 25804
rect 8845 25802 8911 25805
rect 17677 25802 17743 25805
rect 7300 25800 7392 25802
rect 7342 25744 7392 25800
rect 7300 25742 7392 25744
rect 8845 25800 17743 25802
rect 8845 25744 8850 25800
rect 8906 25744 17682 25800
rect 17738 25744 17743 25800
rect 8845 25742 17743 25744
rect 7300 25740 7347 25742
rect 7281 25739 7347 25740
rect 8845 25739 8911 25742
rect 17677 25739 17743 25742
rect 19333 25802 19399 25805
rect 22277 25802 22343 25805
rect 19333 25800 22343 25802
rect 19333 25744 19338 25800
rect 19394 25744 22282 25800
rect 22338 25744 22343 25800
rect 19333 25742 22343 25744
rect 19333 25739 19399 25742
rect 22277 25739 22343 25742
rect 15469 25668 15535 25669
rect 15469 25664 15516 25668
rect 15580 25666 15586 25668
rect 22461 25666 22527 25669
rect 22870 25666 22876 25668
rect 15469 25608 15474 25664
rect 15469 25604 15516 25608
rect 15580 25606 15626 25666
rect 22461 25664 22876 25666
rect 22461 25608 22466 25664
rect 22522 25608 22876 25664
rect 22461 25606 22876 25608
rect 15580 25604 15586 25606
rect 15469 25603 15535 25604
rect 22461 25603 22527 25606
rect 22870 25604 22876 25606
rect 22940 25604 22946 25668
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 11145 25530 11211 25533
rect 16849 25530 16915 25533
rect 11145 25528 16915 25530
rect 11145 25472 11150 25528
rect 11206 25472 16854 25528
rect 16910 25472 16915 25528
rect 11145 25470 16915 25472
rect 11145 25467 11211 25470
rect 16849 25467 16915 25470
rect 6269 25394 6335 25397
rect 7741 25394 7807 25397
rect 15837 25394 15903 25397
rect 6269 25392 7807 25394
rect 6269 25336 6274 25392
rect 6330 25336 7746 25392
rect 7802 25336 7807 25392
rect 6269 25334 7807 25336
rect 6269 25331 6335 25334
rect 7741 25331 7807 25334
rect 9630 25392 15903 25394
rect 9630 25336 15842 25392
rect 15898 25336 15903 25392
rect 9630 25334 15903 25336
rect 200 25258 800 25288
rect 1761 25258 1827 25261
rect 200 25256 1827 25258
rect 200 25200 1766 25256
rect 1822 25200 1827 25256
rect 200 25198 1827 25200
rect 200 25168 800 25198
rect 1761 25195 1827 25198
rect 4429 25258 4495 25261
rect 8109 25258 8175 25261
rect 4429 25256 8175 25258
rect 4429 25200 4434 25256
rect 4490 25200 8114 25256
rect 8170 25200 8175 25256
rect 4429 25198 8175 25200
rect 4429 25195 4495 25198
rect 8109 25195 8175 25198
rect 9630 25125 9690 25334
rect 15837 25331 15903 25334
rect 37641 25258 37707 25261
rect 2037 25122 2103 25125
rect 5993 25122 6059 25125
rect 2037 25120 6059 25122
rect 2037 25064 2042 25120
rect 2098 25064 5998 25120
rect 6054 25064 6059 25120
rect 2037 25062 6059 25064
rect 2037 25059 2103 25062
rect 5993 25059 6059 25062
rect 9581 25120 9690 25125
rect 9581 25064 9586 25120
rect 9642 25064 9690 25120
rect 9581 25062 9690 25064
rect 15334 25256 37707 25258
rect 15334 25200 37646 25256
rect 37702 25200 37707 25256
rect 15334 25198 37707 25200
rect 9581 25059 9647 25062
rect 4981 24986 5047 24989
rect 5901 24988 5967 24989
rect 5206 24986 5212 24988
rect 4981 24984 5212 24986
rect 4981 24928 4986 24984
rect 5042 24928 5212 24984
rect 4981 24926 5212 24928
rect 4981 24923 5047 24926
rect 5206 24924 5212 24926
rect 5276 24924 5282 24988
rect 5901 24984 5948 24988
rect 6012 24986 6018 24988
rect 9121 24986 9187 24989
rect 9857 24986 9923 24989
rect 5901 24928 5906 24984
rect 5901 24924 5948 24928
rect 6012 24926 6058 24986
rect 9121 24984 9923 24986
rect 9121 24928 9126 24984
rect 9182 24928 9862 24984
rect 9918 24928 9923 24984
rect 9121 24926 9923 24928
rect 6012 24924 6018 24926
rect 5901 24923 5967 24924
rect 9121 24923 9187 24926
rect 9857 24923 9923 24926
rect 13854 24924 13860 24988
rect 13924 24986 13930 24988
rect 14549 24986 14615 24989
rect 15334 24986 15394 25198
rect 37641 25195 37707 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 13924 24984 14615 24986
rect 13924 24928 14554 24984
rect 14610 24928 14615 24984
rect 13924 24926 14615 24928
rect 13924 24924 13930 24926
rect 14549 24923 14615 24926
rect 14782 24926 15394 24986
rect 3049 24850 3115 24853
rect 12985 24850 13051 24853
rect 3049 24848 13051 24850
rect 3049 24792 3054 24848
rect 3110 24792 12990 24848
rect 13046 24792 13051 24848
rect 3049 24790 13051 24792
rect 3049 24787 3115 24790
rect 12985 24787 13051 24790
rect 4153 24714 4219 24717
rect 4153 24712 4676 24714
rect 4153 24656 4158 24712
rect 4214 24656 4676 24712
rect 4153 24654 4676 24656
rect 4153 24651 4219 24654
rect 200 24578 800 24608
rect 3417 24578 3483 24581
rect 200 24576 3483 24578
rect 200 24520 3422 24576
rect 3478 24520 3483 24576
rect 200 24518 3483 24520
rect 4616 24578 4676 24654
rect 5574 24652 5580 24716
rect 5644 24714 5650 24716
rect 9121 24714 9187 24717
rect 5644 24712 9187 24714
rect 5644 24656 9126 24712
rect 9182 24656 9187 24712
rect 5644 24654 9187 24656
rect 5644 24652 5650 24654
rect 9121 24651 9187 24654
rect 9990 24652 9996 24716
rect 10060 24714 10066 24716
rect 11053 24714 11119 24717
rect 10060 24712 11119 24714
rect 10060 24656 11058 24712
rect 11114 24656 11119 24712
rect 10060 24654 11119 24656
rect 10060 24652 10066 24654
rect 11053 24651 11119 24654
rect 14641 24714 14707 24717
rect 14782 24714 14842 24926
rect 14641 24712 14842 24714
rect 14641 24656 14646 24712
rect 14702 24656 14842 24712
rect 14641 24654 14842 24656
rect 20161 24714 20227 24717
rect 22277 24714 22343 24717
rect 20161 24712 22343 24714
rect 20161 24656 20166 24712
rect 20222 24656 22282 24712
rect 22338 24656 22343 24712
rect 20161 24654 22343 24656
rect 14641 24651 14707 24654
rect 20161 24651 20227 24654
rect 22277 24651 22343 24654
rect 6729 24578 6795 24581
rect 4616 24576 6795 24578
rect 4616 24520 6734 24576
rect 6790 24520 6795 24576
rect 4616 24518 6795 24520
rect 200 24488 800 24518
rect 3417 24515 3483 24518
rect 6729 24515 6795 24518
rect 11053 24578 11119 24581
rect 18689 24578 18755 24581
rect 11053 24576 18755 24578
rect 11053 24520 11058 24576
rect 11114 24520 18694 24576
rect 18750 24520 18755 24576
rect 11053 24518 18755 24520
rect 11053 24515 11119 24518
rect 18689 24515 18755 24518
rect 38193 24578 38259 24581
rect 39200 24578 39800 24608
rect 38193 24576 39800 24578
rect 38193 24520 38198 24576
rect 38254 24520 39800 24576
rect 38193 24518 39800 24520
rect 38193 24515 38259 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 39800 24518
rect 34930 24447 35246 24448
rect 5073 24442 5139 24445
rect 8109 24442 8175 24445
rect 5073 24440 8175 24442
rect 5073 24384 5078 24440
rect 5134 24384 8114 24440
rect 8170 24384 8175 24440
rect 5073 24382 8175 24384
rect 5073 24379 5139 24382
rect 8109 24379 8175 24382
rect 11697 24442 11763 24445
rect 13905 24442 13971 24445
rect 11697 24440 13971 24442
rect 11697 24384 11702 24440
rect 11758 24384 13910 24440
rect 13966 24384 13971 24440
rect 11697 24382 13971 24384
rect 11697 24379 11763 24382
rect 13905 24379 13971 24382
rect 19701 24442 19767 24445
rect 20110 24442 20116 24444
rect 19701 24440 20116 24442
rect 19701 24384 19706 24440
rect 19762 24384 20116 24440
rect 19701 24382 20116 24384
rect 19701 24379 19767 24382
rect 20110 24380 20116 24382
rect 20180 24380 20186 24444
rect 7741 24306 7807 24309
rect 8477 24306 8543 24309
rect 7741 24304 8543 24306
rect 7741 24248 7746 24304
rect 7802 24248 8482 24304
rect 8538 24248 8543 24304
rect 7741 24246 8543 24248
rect 7741 24243 7807 24246
rect 8477 24243 8543 24246
rect 11278 24244 11284 24308
rect 11348 24306 11354 24308
rect 15837 24306 15903 24309
rect 11348 24304 15903 24306
rect 11348 24248 15842 24304
rect 15898 24248 15903 24304
rect 11348 24246 15903 24248
rect 11348 24244 11354 24246
rect 15837 24243 15903 24246
rect 7097 24170 7163 24173
rect 12750 24170 12756 24172
rect 7097 24168 12756 24170
rect 7097 24112 7102 24168
rect 7158 24112 12756 24168
rect 7097 24110 12756 24112
rect 7097 24107 7163 24110
rect 12750 24108 12756 24110
rect 12820 24108 12826 24172
rect 24485 24170 24551 24173
rect 15334 24168 24551 24170
rect 15334 24112 24490 24168
rect 24546 24112 24551 24168
rect 15334 24110 24551 24112
rect 5901 24034 5967 24037
rect 7557 24034 7623 24037
rect 5901 24032 7623 24034
rect 5901 23976 5906 24032
rect 5962 23976 7562 24032
rect 7618 23976 7623 24032
rect 5901 23974 7623 23976
rect 5901 23971 5967 23974
rect 7557 23971 7623 23974
rect 9673 24034 9739 24037
rect 10225 24034 10291 24037
rect 9673 24032 10291 24034
rect 9673 23976 9678 24032
rect 9734 23976 10230 24032
rect 10286 23976 10291 24032
rect 9673 23974 10291 23976
rect 9673 23971 9739 23974
rect 10225 23971 10291 23974
rect 15101 24034 15167 24037
rect 15334 24034 15394 24110
rect 24485 24107 24551 24110
rect 15101 24032 15394 24034
rect 15101 23976 15106 24032
rect 15162 23976 15394 24032
rect 15101 23974 15394 23976
rect 15101 23971 15167 23974
rect 16798 23972 16804 24036
rect 16868 24034 16874 24036
rect 19425 24034 19491 24037
rect 16868 24032 19491 24034
rect 16868 23976 19430 24032
rect 19486 23976 19491 24032
rect 16868 23974 19491 23976
rect 16868 23972 16874 23974
rect 19425 23971 19491 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4061 23898 4127 23901
rect 6913 23898 6979 23901
rect 8937 23898 9003 23901
rect 4061 23896 6979 23898
rect 4061 23840 4066 23896
rect 4122 23840 6918 23896
rect 6974 23840 6979 23896
rect 4061 23838 6979 23840
rect 4061 23835 4127 23838
rect 6913 23835 6979 23838
rect 7054 23896 9003 23898
rect 7054 23840 8942 23896
rect 8998 23840 9003 23896
rect 7054 23838 9003 23840
rect 3233 23762 3299 23765
rect 7054 23762 7114 23838
rect 8937 23835 9003 23838
rect 10041 23898 10107 23901
rect 13813 23898 13879 23901
rect 16389 23898 16455 23901
rect 17861 23898 17927 23901
rect 10041 23896 13879 23898
rect 10041 23840 10046 23896
rect 10102 23840 13818 23896
rect 13874 23840 13879 23896
rect 10041 23838 13879 23840
rect 10041 23835 10107 23838
rect 13813 23835 13879 23838
rect 15886 23896 17927 23898
rect 15886 23840 16394 23896
rect 16450 23840 17866 23896
rect 17922 23840 17927 23896
rect 15886 23838 17927 23840
rect 3233 23760 7114 23762
rect 3233 23704 3238 23760
rect 3294 23704 7114 23760
rect 3233 23702 7114 23704
rect 7465 23762 7531 23765
rect 9949 23762 10015 23765
rect 15886 23762 15946 23838
rect 16389 23835 16455 23838
rect 17861 23835 17927 23838
rect 37457 23898 37523 23901
rect 39200 23898 39800 23928
rect 37457 23896 39800 23898
rect 37457 23840 37462 23896
rect 37518 23840 39800 23896
rect 37457 23838 39800 23840
rect 37457 23835 37523 23838
rect 39200 23808 39800 23838
rect 7465 23760 10015 23762
rect 7465 23704 7470 23760
rect 7526 23704 9954 23760
rect 10010 23704 10015 23760
rect 7465 23702 10015 23704
rect 3233 23699 3299 23702
rect 7465 23699 7531 23702
rect 9949 23699 10015 23702
rect 12390 23702 15946 23762
rect 16021 23762 16087 23765
rect 22461 23762 22527 23765
rect 16021 23760 22527 23762
rect 16021 23704 16026 23760
rect 16082 23704 22466 23760
rect 22522 23704 22527 23760
rect 16021 23702 22527 23704
rect 12390 23626 12450 23702
rect 16021 23699 16087 23702
rect 22461 23699 22527 23702
rect 8526 23566 12450 23626
rect 13721 23626 13787 23629
rect 17217 23626 17283 23629
rect 17953 23626 18019 23629
rect 13721 23624 18019 23626
rect 13721 23568 13726 23624
rect 13782 23568 17222 23624
rect 17278 23568 17958 23624
rect 18014 23568 18019 23624
rect 13721 23566 18019 23568
rect 105 23490 171 23493
rect 62 23488 171 23490
rect 62 23432 110 23488
rect 166 23432 171 23488
rect 62 23427 171 23432
rect 5257 23490 5323 23493
rect 5574 23490 5580 23492
rect 5257 23488 5580 23490
rect 5257 23432 5262 23488
rect 5318 23432 5580 23488
rect 5257 23430 5580 23432
rect 5257 23427 5323 23430
rect 5574 23428 5580 23430
rect 5644 23428 5650 23492
rect 6545 23490 6611 23493
rect 8109 23490 8175 23493
rect 6545 23488 8175 23490
rect 6545 23432 6550 23488
rect 6606 23432 8114 23488
rect 8170 23432 8175 23488
rect 6545 23430 8175 23432
rect 6545 23427 6611 23430
rect 8109 23427 8175 23430
rect 62 23218 122 23427
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 6729 23354 6795 23357
rect 8526 23354 8586 23566
rect 13721 23563 13787 23566
rect 17217 23563 17283 23566
rect 17953 23563 18019 23566
rect 8845 23492 8911 23493
rect 8845 23488 8892 23492
rect 8956 23490 8962 23492
rect 8845 23432 8850 23488
rect 8845 23428 8892 23432
rect 8956 23430 9002 23490
rect 8956 23428 8962 23430
rect 10542 23428 10548 23492
rect 10612 23490 10618 23492
rect 11053 23490 11119 23493
rect 10612 23488 11119 23490
rect 10612 23432 11058 23488
rect 11114 23432 11119 23488
rect 10612 23430 11119 23432
rect 10612 23428 10618 23430
rect 8845 23427 8911 23428
rect 11053 23427 11119 23430
rect 12157 23490 12223 23493
rect 12617 23490 12683 23493
rect 15285 23490 15351 23493
rect 12157 23488 12683 23490
rect 12157 23432 12162 23488
rect 12218 23432 12622 23488
rect 12678 23432 12683 23488
rect 12157 23430 12683 23432
rect 12157 23427 12223 23430
rect 12617 23427 12683 23430
rect 12758 23488 15351 23490
rect 12758 23432 15290 23488
rect 15346 23432 15351 23488
rect 12758 23430 15351 23432
rect 6729 23352 8586 23354
rect 6729 23296 6734 23352
rect 6790 23296 8586 23352
rect 6729 23294 8586 23296
rect 9305 23354 9371 23357
rect 10777 23354 10843 23357
rect 9305 23352 10843 23354
rect 9305 23296 9310 23352
rect 9366 23296 10782 23352
rect 10838 23296 10843 23352
rect 9305 23294 10843 23296
rect 6729 23291 6795 23294
rect 9305 23291 9371 23294
rect 10777 23291 10843 23294
rect 11237 23354 11303 23357
rect 12758 23354 12818 23430
rect 15285 23427 15351 23430
rect 21766 23428 21772 23492
rect 21836 23490 21842 23492
rect 21909 23490 21975 23493
rect 21836 23488 21975 23490
rect 21836 23432 21914 23488
rect 21970 23432 21975 23488
rect 21836 23430 21975 23432
rect 21836 23428 21842 23430
rect 21909 23427 21975 23430
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 11237 23352 12818 23354
rect 11237 23296 11242 23352
rect 11298 23296 12818 23352
rect 11237 23294 12818 23296
rect 11237 23291 11303 23294
rect 12934 23292 12940 23356
rect 13004 23354 13010 23356
rect 13537 23354 13603 23357
rect 13004 23352 13603 23354
rect 13004 23296 13542 23352
rect 13598 23296 13603 23352
rect 13004 23294 13603 23296
rect 13004 23292 13010 23294
rect 13537 23291 13603 23294
rect 19149 23354 19215 23357
rect 23565 23354 23631 23357
rect 19149 23352 23631 23354
rect 19149 23296 19154 23352
rect 19210 23296 23570 23352
rect 23626 23296 23631 23352
rect 19149 23294 23631 23296
rect 19149 23291 19215 23294
rect 23565 23291 23631 23294
rect 200 23218 800 23248
rect 5073 23220 5139 23221
rect 5022 23218 5028 23220
rect 62 23158 800 23218
rect 4982 23158 5028 23218
rect 5092 23216 5139 23220
rect 5134 23160 5139 23216
rect 200 23128 800 23158
rect 5022 23156 5028 23158
rect 5092 23156 5139 23160
rect 5206 23156 5212 23220
rect 5276 23218 5282 23220
rect 26417 23218 26483 23221
rect 5276 23216 26483 23218
rect 5276 23160 26422 23216
rect 26478 23160 26483 23216
rect 5276 23158 26483 23160
rect 5276 23156 5282 23158
rect 5073 23155 5139 23156
rect 26417 23155 26483 23158
rect 1485 23082 1551 23085
rect 1485 23080 2790 23082
rect 1485 23024 1490 23080
rect 1546 23024 2790 23080
rect 1485 23022 2790 23024
rect 1485 23019 1551 23022
rect 2730 22810 2790 23022
rect 5022 23020 5028 23084
rect 5092 23082 5098 23084
rect 5717 23082 5783 23085
rect 9765 23084 9831 23085
rect 9765 23082 9812 23084
rect 5092 23080 5783 23082
rect 5092 23024 5722 23080
rect 5778 23024 5783 23080
rect 5092 23022 5783 23024
rect 9720 23080 9812 23082
rect 9720 23024 9770 23080
rect 9720 23022 9812 23024
rect 5092 23020 5098 23022
rect 5717 23019 5783 23022
rect 9765 23020 9812 23022
rect 9876 23020 9882 23084
rect 12249 23082 12315 23085
rect 13261 23082 13327 23085
rect 12249 23080 13327 23082
rect 12249 23024 12254 23080
rect 12310 23024 13266 23080
rect 13322 23024 13327 23080
rect 12249 23022 13327 23024
rect 9765 23019 9874 23020
rect 12249 23019 12315 23022
rect 13261 23019 13327 23022
rect 14457 23082 14523 23085
rect 21909 23082 21975 23085
rect 27061 23082 27127 23085
rect 14457 23080 21282 23082
rect 14457 23024 14462 23080
rect 14518 23024 21282 23080
rect 14457 23022 21282 23024
rect 14457 23019 14523 23022
rect 5441 22946 5507 22949
rect 8334 22946 8340 22948
rect 5441 22944 8340 22946
rect 5441 22888 5446 22944
rect 5502 22888 8340 22944
rect 5441 22886 8340 22888
rect 5441 22883 5507 22886
rect 8334 22884 8340 22886
rect 8404 22884 8410 22948
rect 9814 22946 9874 23019
rect 21222 22946 21282 23022
rect 21909 23080 27127 23082
rect 21909 23024 21914 23080
rect 21970 23024 27066 23080
rect 27122 23024 27127 23080
rect 21909 23022 27127 23024
rect 21909 23019 21975 23022
rect 27061 23019 27127 23022
rect 24710 22946 24716 22948
rect 9814 22886 17234 22946
rect 21222 22886 24716 22946
rect 7414 22810 7420 22812
rect 2730 22750 7420 22810
rect 7414 22748 7420 22750
rect 7484 22748 7490 22812
rect 12433 22810 12499 22813
rect 15561 22810 15627 22813
rect 12433 22808 15627 22810
rect 12433 22752 12438 22808
rect 12494 22752 15566 22808
rect 15622 22752 15627 22808
rect 12433 22750 15627 22752
rect 12433 22747 12499 22750
rect 15561 22747 15627 22750
rect 16665 22810 16731 22813
rect 16982 22810 16988 22812
rect 16665 22808 16988 22810
rect 16665 22752 16670 22808
rect 16726 22752 16988 22808
rect 16665 22750 16988 22752
rect 16665 22747 16731 22750
rect 16982 22748 16988 22750
rect 17052 22748 17058 22812
rect 11513 22674 11579 22677
rect 12249 22674 12315 22677
rect 13537 22674 13603 22677
rect 11513 22672 13603 22674
rect 11513 22616 11518 22672
rect 11574 22616 12254 22672
rect 12310 22616 13542 22672
rect 13598 22616 13603 22672
rect 11513 22614 13603 22616
rect 11513 22611 11579 22614
rect 12249 22611 12315 22614
rect 13537 22611 13603 22614
rect 13905 22674 13971 22677
rect 16573 22674 16639 22677
rect 13905 22672 16639 22674
rect 13905 22616 13910 22672
rect 13966 22616 16578 22672
rect 16634 22616 16639 22672
rect 13905 22614 16639 22616
rect 17174 22674 17234 22886
rect 24710 22884 24716 22886
rect 24780 22884 24786 22948
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 20345 22810 20411 22813
rect 22737 22810 22803 22813
rect 20345 22808 22803 22810
rect 20345 22752 20350 22808
rect 20406 22752 22742 22808
rect 22798 22752 22803 22808
rect 20345 22750 22803 22752
rect 20345 22747 20411 22750
rect 22737 22747 22803 22750
rect 21817 22674 21883 22677
rect 17174 22672 21883 22674
rect 17174 22616 21822 22672
rect 21878 22616 21883 22672
rect 17174 22614 21883 22616
rect 13905 22611 13971 22614
rect 16573 22611 16639 22614
rect 21817 22611 21883 22614
rect 200 22538 800 22568
rect 1577 22538 1643 22541
rect 200 22536 1643 22538
rect 200 22480 1582 22536
rect 1638 22480 1643 22536
rect 200 22478 1643 22480
rect 200 22448 800 22478
rect 1577 22475 1643 22478
rect 11237 22538 11303 22541
rect 17953 22538 18019 22541
rect 11237 22536 18019 22538
rect 11237 22480 11242 22536
rect 11298 22480 17958 22536
rect 18014 22480 18019 22536
rect 11237 22478 18019 22480
rect 11237 22475 11303 22478
rect 17953 22475 18019 22478
rect 19517 22538 19583 22541
rect 20713 22538 20779 22541
rect 19517 22536 20779 22538
rect 19517 22480 19522 22536
rect 19578 22480 20718 22536
rect 20774 22480 20779 22536
rect 19517 22478 20779 22480
rect 19517 22475 19583 22478
rect 20713 22475 20779 22478
rect 21265 22538 21331 22541
rect 23289 22538 23355 22541
rect 21265 22536 23355 22538
rect 21265 22480 21270 22536
rect 21326 22480 23294 22536
rect 23350 22480 23355 22536
rect 21265 22478 23355 22480
rect 21265 22475 21331 22478
rect 23289 22475 23355 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 11421 22402 11487 22405
rect 12249 22402 12315 22405
rect 11421 22400 12315 22402
rect 11421 22344 11426 22400
rect 11482 22344 12254 22400
rect 12310 22344 12315 22400
rect 11421 22342 12315 22344
rect 11421 22339 11487 22342
rect 12249 22339 12315 22342
rect 12801 22402 12867 22405
rect 12934 22402 12940 22404
rect 12801 22400 12940 22402
rect 12801 22344 12806 22400
rect 12862 22344 12940 22400
rect 12801 22342 12940 22344
rect 12801 22339 12867 22342
rect 12934 22340 12940 22342
rect 13004 22340 13010 22404
rect 13118 22340 13124 22404
rect 13188 22402 13194 22404
rect 15653 22402 15719 22405
rect 18689 22402 18755 22405
rect 13188 22342 14106 22402
rect 13188 22340 13194 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 5758 22204 5764 22268
rect 5828 22266 5834 22268
rect 5993 22266 6059 22269
rect 5828 22264 6059 22266
rect 5828 22208 5998 22264
rect 6054 22208 6059 22264
rect 5828 22206 6059 22208
rect 5828 22204 5834 22206
rect 5993 22203 6059 22206
rect 8017 22266 8083 22269
rect 12709 22266 12775 22269
rect 14046 22266 14106 22342
rect 15653 22400 18755 22402
rect 15653 22344 15658 22400
rect 15714 22344 18694 22400
rect 18750 22344 18755 22400
rect 15653 22342 18755 22344
rect 15653 22339 15719 22342
rect 18689 22339 18755 22342
rect 23197 22402 23263 22405
rect 24945 22402 25011 22405
rect 29177 22402 29243 22405
rect 23197 22400 29243 22402
rect 23197 22344 23202 22400
rect 23258 22344 24950 22400
rect 25006 22344 29182 22400
rect 29238 22344 29243 22400
rect 23197 22342 29243 22344
rect 23197 22339 23263 22342
rect 24945 22339 25011 22342
rect 29177 22339 29243 22342
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 18873 22266 18939 22269
rect 8017 22264 12634 22266
rect 8017 22208 8022 22264
rect 8078 22208 12634 22264
rect 8017 22206 12634 22208
rect 8017 22203 8083 22206
rect 7557 22130 7623 22133
rect 8017 22130 8083 22133
rect 7557 22128 8083 22130
rect 7557 22072 7562 22128
rect 7618 22072 8022 22128
rect 8078 22072 8083 22128
rect 7557 22070 8083 22072
rect 7557 22067 7623 22070
rect 8017 22067 8083 22070
rect 9438 22068 9444 22132
rect 9508 22130 9514 22132
rect 12382 22130 12388 22132
rect 9508 22070 12388 22130
rect 9508 22068 9514 22070
rect 12382 22068 12388 22070
rect 12452 22068 12458 22132
rect 3693 21994 3759 21997
rect 4797 21994 4863 21997
rect 3693 21992 4863 21994
rect 3693 21936 3698 21992
rect 3754 21936 4802 21992
rect 4858 21936 4863 21992
rect 3693 21934 4863 21936
rect 3693 21931 3759 21934
rect 4797 21931 4863 21934
rect 5758 21932 5764 21996
rect 5828 21994 5834 21996
rect 5993 21994 6059 21997
rect 5828 21992 6059 21994
rect 5828 21936 5998 21992
rect 6054 21936 6059 21992
rect 5828 21934 6059 21936
rect 5828 21932 5834 21934
rect 5993 21931 6059 21934
rect 7281 21994 7347 21997
rect 8661 21994 8727 21997
rect 7281 21992 8727 21994
rect 7281 21936 7286 21992
rect 7342 21936 8666 21992
rect 8722 21936 8727 21992
rect 7281 21934 8727 21936
rect 7281 21931 7347 21934
rect 8661 21931 8727 21934
rect 8845 21994 8911 21997
rect 11053 21994 11119 21997
rect 8845 21992 11119 21994
rect 8845 21936 8850 21992
rect 8906 21936 11058 21992
rect 11114 21936 11119 21992
rect 8845 21934 11119 21936
rect 8845 21931 8911 21934
rect 11053 21931 11119 21934
rect 11329 21994 11395 21997
rect 11881 21994 11947 21997
rect 11329 21992 11947 21994
rect 11329 21936 11334 21992
rect 11390 21936 11886 21992
rect 11942 21936 11947 21992
rect 11329 21934 11947 21936
rect 12574 21994 12634 22206
rect 12709 22264 13922 22266
rect 12709 22208 12714 22264
rect 12770 22208 13922 22264
rect 12709 22206 13922 22208
rect 14046 22264 18939 22266
rect 14046 22208 18878 22264
rect 18934 22208 18939 22264
rect 14046 22206 18939 22208
rect 12709 22203 12775 22206
rect 12750 22068 12756 22132
rect 12820 22130 12826 22132
rect 13169 22130 13235 22133
rect 13862 22130 13922 22206
rect 18873 22203 18939 22206
rect 20069 22266 20135 22269
rect 24853 22266 24919 22269
rect 20069 22264 24919 22266
rect 20069 22208 20074 22264
rect 20130 22208 24858 22264
rect 24914 22208 24919 22264
rect 20069 22206 24919 22208
rect 20069 22203 20135 22206
rect 24853 22203 24919 22206
rect 14457 22130 14523 22133
rect 12820 22128 13738 22130
rect 12820 22072 13174 22128
rect 13230 22072 13738 22128
rect 12820 22070 13738 22072
rect 13862 22128 14523 22130
rect 13862 22072 14462 22128
rect 14518 22072 14523 22128
rect 13862 22070 14523 22072
rect 12820 22068 12826 22070
rect 13169 22067 13235 22070
rect 13486 21994 13492 21996
rect 12574 21934 13492 21994
rect 11329 21931 11395 21934
rect 11881 21931 11947 21934
rect 13486 21932 13492 21934
rect 13556 21932 13562 21996
rect 13678 21994 13738 22070
rect 14457 22067 14523 22070
rect 17953 22130 18019 22133
rect 18781 22130 18847 22133
rect 21633 22130 21699 22133
rect 17953 22128 21699 22130
rect 17953 22072 17958 22128
rect 18014 22072 18786 22128
rect 18842 22072 21638 22128
rect 21694 22072 21699 22128
rect 17953 22070 21699 22072
rect 17953 22067 18019 22070
rect 18781 22067 18847 22070
rect 21633 22067 21699 22070
rect 22686 22068 22692 22132
rect 22756 22130 22762 22132
rect 23289 22130 23355 22133
rect 27797 22130 27863 22133
rect 22756 22128 23355 22130
rect 22756 22072 23294 22128
rect 23350 22072 23355 22128
rect 22756 22070 23355 22072
rect 22756 22068 22762 22070
rect 23289 22067 23355 22070
rect 23430 22128 27863 22130
rect 23430 22072 27802 22128
rect 27858 22072 27863 22128
rect 23430 22070 27863 22072
rect 23013 21994 23079 21997
rect 13678 21992 23079 21994
rect 13678 21936 23018 21992
rect 23074 21936 23079 21992
rect 13678 21934 23079 21936
rect 23013 21931 23079 21934
rect 2405 21858 2471 21861
rect 8569 21858 8635 21861
rect 2405 21856 8635 21858
rect 2405 21800 2410 21856
rect 2466 21800 8574 21856
rect 8630 21800 8635 21856
rect 2405 21798 8635 21800
rect 2405 21795 2471 21798
rect 8569 21795 8635 21798
rect 10501 21858 10567 21861
rect 18045 21858 18111 21861
rect 10501 21856 18111 21858
rect 10501 21800 10506 21856
rect 10562 21800 18050 21856
rect 18106 21800 18111 21856
rect 10501 21798 18111 21800
rect 10501 21795 10567 21798
rect 18045 21795 18111 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4613 21722 4679 21725
rect 4889 21722 4955 21725
rect 4613 21720 4955 21722
rect 4613 21664 4618 21720
rect 4674 21664 4894 21720
rect 4950 21664 4955 21720
rect 4613 21662 4955 21664
rect 4613 21659 4679 21662
rect 4889 21659 4955 21662
rect 7465 21722 7531 21725
rect 7833 21722 7899 21725
rect 7465 21720 7899 21722
rect 7465 21664 7470 21720
rect 7526 21664 7838 21720
rect 7894 21664 7899 21720
rect 7465 21662 7899 21664
rect 7465 21659 7531 21662
rect 7833 21659 7899 21662
rect 10041 21722 10107 21725
rect 15193 21722 15259 21725
rect 10041 21720 15259 21722
rect 10041 21664 10046 21720
rect 10102 21664 15198 21720
rect 15254 21664 15259 21720
rect 10041 21662 15259 21664
rect 10041 21659 10107 21662
rect 15193 21659 15259 21662
rect 15377 21722 15443 21725
rect 16481 21722 16547 21725
rect 15377 21720 16547 21722
rect 15377 21664 15382 21720
rect 15438 21664 16486 21720
rect 16542 21664 16547 21720
rect 15377 21662 16547 21664
rect 15377 21659 15443 21662
rect 16481 21659 16547 21662
rect 17861 21722 17927 21725
rect 19425 21722 19491 21725
rect 17861 21720 19491 21722
rect 17861 21664 17866 21720
rect 17922 21664 19430 21720
rect 19486 21664 19491 21720
rect 17861 21662 19491 21664
rect 17861 21659 17927 21662
rect 19425 21659 19491 21662
rect 21909 21722 21975 21725
rect 22645 21722 22711 21725
rect 21909 21720 22711 21722
rect 21909 21664 21914 21720
rect 21970 21664 22650 21720
rect 22706 21664 22711 21720
rect 21909 21662 22711 21664
rect 21909 21659 21975 21662
rect 22645 21659 22711 21662
rect 23013 21722 23079 21725
rect 23197 21722 23263 21725
rect 23013 21720 23263 21722
rect 23013 21664 23018 21720
rect 23074 21664 23202 21720
rect 23258 21664 23263 21720
rect 23013 21662 23263 21664
rect 23013 21659 23079 21662
rect 23197 21659 23263 21662
rect 1945 21588 2011 21589
rect 1894 21524 1900 21588
rect 1964 21586 2011 21588
rect 1964 21584 2056 21586
rect 2006 21528 2056 21584
rect 1964 21526 2056 21528
rect 1964 21524 2011 21526
rect 9622 21524 9628 21588
rect 9692 21586 9698 21588
rect 10501 21586 10567 21589
rect 9692 21584 10567 21586
rect 9692 21528 10506 21584
rect 10562 21528 10567 21584
rect 9692 21526 10567 21528
rect 9692 21524 9698 21526
rect 1945 21523 2011 21524
rect 10501 21523 10567 21526
rect 10685 21586 10751 21589
rect 13077 21586 13143 21589
rect 10685 21584 13143 21586
rect 10685 21528 10690 21584
rect 10746 21528 13082 21584
rect 13138 21528 13143 21584
rect 10685 21526 13143 21528
rect 10685 21523 10751 21526
rect 13077 21523 13143 21526
rect 13813 21586 13879 21589
rect 22829 21586 22895 21589
rect 23430 21586 23490 22070
rect 27797 22067 27863 22070
rect 26877 21996 26943 21997
rect 26877 21994 26924 21996
rect 26832 21992 26924 21994
rect 26988 21994 26994 21996
rect 29085 21994 29151 21997
rect 26988 21992 29151 21994
rect 26832 21936 26882 21992
rect 26988 21936 29090 21992
rect 29146 21936 29151 21992
rect 26832 21934 26924 21936
rect 26877 21932 26924 21934
rect 26988 21934 29151 21936
rect 26988 21932 26994 21934
rect 26877 21931 26943 21932
rect 29085 21931 29151 21934
rect 38285 21858 38351 21861
rect 39200 21858 39800 21888
rect 38285 21856 39800 21858
rect 38285 21800 38290 21856
rect 38346 21800 39800 21856
rect 38285 21798 39800 21800
rect 38285 21795 38351 21798
rect 39200 21768 39800 21798
rect 38193 21722 38259 21725
rect 13813 21584 23490 21586
rect 13813 21528 13818 21584
rect 13874 21528 22834 21584
rect 22890 21528 23490 21584
rect 13813 21526 23490 21528
rect 31710 21720 38259 21722
rect 31710 21664 38198 21720
rect 38254 21664 38259 21720
rect 31710 21662 38259 21664
rect 13813 21523 13879 21526
rect 22829 21523 22895 21526
rect 6637 21450 6703 21453
rect 9121 21450 9187 21453
rect 6637 21448 9187 21450
rect 6637 21392 6642 21448
rect 6698 21392 9126 21448
rect 9182 21392 9187 21448
rect 6637 21390 9187 21392
rect 6637 21387 6703 21390
rect 9121 21387 9187 21390
rect 10685 21450 10751 21453
rect 10869 21450 10935 21453
rect 10685 21448 10935 21450
rect 10685 21392 10690 21448
rect 10746 21392 10874 21448
rect 10930 21392 10935 21448
rect 10685 21390 10935 21392
rect 10685 21387 10751 21390
rect 10869 21387 10935 21390
rect 11237 21450 11303 21453
rect 11881 21450 11947 21453
rect 13721 21450 13787 21453
rect 11237 21448 13787 21450
rect 11237 21392 11242 21448
rect 11298 21392 11886 21448
rect 11942 21392 13726 21448
rect 13782 21392 13787 21448
rect 11237 21390 13787 21392
rect 11237 21387 11303 21390
rect 11881 21387 11947 21390
rect 13721 21387 13787 21390
rect 14590 21388 14596 21452
rect 14660 21450 14666 21452
rect 17125 21450 17191 21453
rect 14660 21448 17191 21450
rect 14660 21392 17130 21448
rect 17186 21392 17191 21448
rect 14660 21390 17191 21392
rect 14660 21388 14666 21390
rect 17125 21387 17191 21390
rect 18505 21450 18571 21453
rect 18822 21450 18828 21452
rect 18505 21448 18828 21450
rect 18505 21392 18510 21448
rect 18566 21392 18828 21448
rect 18505 21390 18828 21392
rect 18505 21387 18571 21390
rect 18822 21388 18828 21390
rect 18892 21388 18898 21452
rect 19057 21450 19123 21453
rect 22185 21450 22251 21453
rect 19057 21448 22251 21450
rect 19057 21392 19062 21448
rect 19118 21392 22190 21448
rect 22246 21392 22251 21448
rect 19057 21390 22251 21392
rect 19057 21387 19123 21390
rect 22185 21387 22251 21390
rect 23289 21450 23355 21453
rect 31710 21450 31770 21662
rect 38193 21659 38259 21662
rect 23289 21448 31770 21450
rect 23289 21392 23294 21448
rect 23350 21392 31770 21448
rect 23289 21390 31770 21392
rect 23289 21387 23355 21390
rect 3325 21314 3391 21317
rect 3734 21314 3740 21316
rect 3325 21312 3740 21314
rect 3325 21256 3330 21312
rect 3386 21256 3740 21312
rect 3325 21254 3740 21256
rect 3325 21251 3391 21254
rect 3734 21252 3740 21254
rect 3804 21252 3810 21316
rect 5165 21314 5231 21317
rect 5390 21314 5396 21316
rect 5165 21312 5396 21314
rect 5165 21256 5170 21312
rect 5226 21256 5396 21312
rect 5165 21254 5396 21256
rect 5165 21251 5231 21254
rect 5390 21252 5396 21254
rect 5460 21314 5466 21316
rect 7465 21314 7531 21317
rect 5460 21312 7531 21314
rect 5460 21256 7470 21312
rect 7526 21256 7531 21312
rect 5460 21254 7531 21256
rect 5460 21252 5466 21254
rect 7465 21251 7531 21254
rect 9305 21314 9371 21317
rect 12750 21314 12756 21316
rect 9305 21312 12756 21314
rect 9305 21256 9310 21312
rect 9366 21256 12756 21312
rect 9305 21254 12756 21256
rect 9305 21251 9371 21254
rect 12750 21252 12756 21254
rect 12820 21252 12826 21316
rect 12985 21314 13051 21317
rect 19517 21314 19583 21317
rect 21357 21314 21423 21317
rect 12985 21312 19442 21314
rect 12985 21256 12990 21312
rect 13046 21256 19442 21312
rect 12985 21254 19442 21256
rect 12985 21251 13051 21254
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 3969 21178 4035 21181
rect 200 21176 4035 21178
rect 200 21120 3974 21176
rect 4030 21120 4035 21176
rect 200 21118 4035 21120
rect 200 21088 800 21118
rect 3969 21115 4035 21118
rect 5022 21116 5028 21180
rect 5092 21178 5098 21180
rect 5165 21178 5231 21181
rect 5092 21176 5231 21178
rect 5092 21120 5170 21176
rect 5226 21120 5231 21176
rect 5092 21118 5231 21120
rect 5092 21116 5098 21118
rect 5165 21115 5231 21118
rect 8201 21178 8267 21181
rect 19190 21178 19196 21180
rect 8201 21176 19196 21178
rect 8201 21120 8206 21176
rect 8262 21120 19196 21176
rect 8201 21118 19196 21120
rect 8201 21115 8267 21118
rect 19190 21116 19196 21118
rect 19260 21116 19266 21180
rect 19382 21178 19442 21254
rect 19517 21312 21423 21314
rect 19517 21256 19522 21312
rect 19578 21256 21362 21312
rect 21418 21256 21423 21312
rect 19517 21254 21423 21256
rect 19517 21251 19583 21254
rect 21357 21251 21423 21254
rect 22553 21314 22619 21317
rect 28625 21314 28691 21317
rect 22553 21312 28691 21314
rect 22553 21256 22558 21312
rect 22614 21256 28630 21312
rect 28686 21256 28691 21312
rect 22553 21254 28691 21256
rect 22553 21251 22619 21254
rect 28625 21251 28691 21254
rect 22556 21178 22616 21251
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19382 21118 22616 21178
rect 38101 21178 38167 21181
rect 39200 21178 39800 21208
rect 38101 21176 39800 21178
rect 38101 21120 38106 21176
rect 38162 21120 39800 21176
rect 38101 21118 39800 21120
rect 38101 21115 38167 21118
rect 39200 21088 39800 21118
rect 6821 21042 6887 21045
rect 10174 21042 10180 21044
rect 6821 21040 10180 21042
rect 6821 20984 6826 21040
rect 6882 20984 10180 21040
rect 6821 20982 10180 20984
rect 6821 20979 6887 20982
rect 10174 20980 10180 20982
rect 10244 20980 10250 21044
rect 10869 21042 10935 21045
rect 12525 21042 12591 21045
rect 10869 21040 12591 21042
rect 10869 20984 10874 21040
rect 10930 20984 12530 21040
rect 12586 20984 12591 21040
rect 10869 20982 12591 20984
rect 10869 20979 10935 20982
rect 12525 20979 12591 20982
rect 14181 21042 14247 21045
rect 18137 21042 18203 21045
rect 14181 21040 18203 21042
rect 14181 20984 14186 21040
rect 14242 20984 18142 21040
rect 18198 20984 18203 21040
rect 14181 20982 18203 20984
rect 14181 20979 14247 20982
rect 18137 20979 18203 20982
rect 19190 20980 19196 21044
rect 19260 21042 19266 21044
rect 24117 21042 24183 21045
rect 19260 21040 24183 21042
rect 19260 20984 24122 21040
rect 24178 20984 24183 21040
rect 19260 20982 24183 20984
rect 19260 20980 19266 20982
rect 24117 20979 24183 20982
rect 3049 20906 3115 20909
rect 9254 20906 9260 20908
rect 3049 20904 9260 20906
rect 3049 20848 3054 20904
rect 3110 20848 9260 20904
rect 3049 20846 9260 20848
rect 3049 20843 3115 20846
rect 9254 20844 9260 20846
rect 9324 20844 9330 20908
rect 9806 20844 9812 20908
rect 9876 20906 9882 20908
rect 12341 20906 12407 20909
rect 9876 20904 12407 20906
rect 9876 20848 12346 20904
rect 12402 20848 12407 20904
rect 9876 20846 12407 20848
rect 9876 20844 9882 20846
rect 12341 20843 12407 20846
rect 12525 20906 12591 20909
rect 15009 20906 15075 20909
rect 12525 20904 15075 20906
rect 12525 20848 12530 20904
rect 12586 20848 15014 20904
rect 15070 20848 15075 20904
rect 12525 20846 15075 20848
rect 12525 20843 12591 20846
rect 15009 20843 15075 20846
rect 16021 20906 16087 20909
rect 25957 20906 26023 20909
rect 16021 20904 26023 20906
rect 16021 20848 16026 20904
rect 16082 20848 25962 20904
rect 26018 20848 26023 20904
rect 16021 20846 26023 20848
rect 16021 20843 16087 20846
rect 25957 20843 26023 20846
rect 5073 20770 5139 20773
rect 6678 20770 6684 20772
rect 5073 20768 6684 20770
rect 5073 20712 5078 20768
rect 5134 20712 6684 20768
rect 5073 20710 6684 20712
rect 5073 20707 5139 20710
rect 6678 20708 6684 20710
rect 6748 20708 6754 20772
rect 8201 20770 8267 20773
rect 14457 20770 14523 20773
rect 15561 20772 15627 20773
rect 15510 20770 15516 20772
rect 8201 20768 14523 20770
rect 8201 20712 8206 20768
rect 8262 20712 14462 20768
rect 14518 20712 14523 20768
rect 8201 20710 14523 20712
rect 15434 20710 15516 20770
rect 15580 20770 15627 20772
rect 16113 20770 16179 20773
rect 15580 20768 16179 20770
rect 15622 20712 16118 20768
rect 16174 20712 16179 20768
rect 8201 20707 8267 20710
rect 14457 20707 14523 20710
rect 15510 20708 15516 20710
rect 15580 20710 16179 20712
rect 15580 20708 15627 20710
rect 15561 20707 15627 20708
rect 16113 20707 16179 20710
rect 16665 20770 16731 20773
rect 17861 20770 17927 20773
rect 16665 20768 17927 20770
rect 16665 20712 16670 20768
rect 16726 20712 17866 20768
rect 17922 20712 17927 20768
rect 16665 20710 17927 20712
rect 16665 20707 16731 20710
rect 17861 20707 17927 20710
rect 19149 20770 19215 20773
rect 19425 20770 19491 20773
rect 20161 20772 20227 20773
rect 19149 20768 19491 20770
rect 19149 20712 19154 20768
rect 19210 20712 19430 20768
rect 19486 20712 19491 20768
rect 19149 20710 19491 20712
rect 19149 20707 19215 20710
rect 19425 20707 19491 20710
rect 20110 20708 20116 20772
rect 20180 20770 20227 20772
rect 20345 20770 20411 20773
rect 24945 20770 25011 20773
rect 20180 20768 20272 20770
rect 20222 20712 20272 20768
rect 20180 20710 20272 20712
rect 20345 20768 25011 20770
rect 20345 20712 20350 20768
rect 20406 20712 24950 20768
rect 25006 20712 25011 20768
rect 20345 20710 25011 20712
rect 20180 20708 20227 20710
rect 20161 20707 20227 20708
rect 20345 20707 20411 20710
rect 24945 20707 25011 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4797 20634 4863 20637
rect 9029 20634 9095 20637
rect 4797 20632 9095 20634
rect 4797 20576 4802 20632
rect 4858 20576 9034 20632
rect 9090 20576 9095 20632
rect 4797 20574 9095 20576
rect 4797 20571 4863 20574
rect 9029 20571 9095 20574
rect 9213 20634 9279 20637
rect 12198 20634 12204 20636
rect 9213 20632 12204 20634
rect 9213 20576 9218 20632
rect 9274 20576 12204 20632
rect 9213 20574 12204 20576
rect 9213 20571 9279 20574
rect 12198 20572 12204 20574
rect 12268 20572 12274 20636
rect 12382 20572 12388 20636
rect 12452 20634 12458 20636
rect 17953 20634 18019 20637
rect 12452 20632 18019 20634
rect 12452 20576 17958 20632
rect 18014 20576 18019 20632
rect 12452 20574 18019 20576
rect 12452 20572 12458 20574
rect 17953 20571 18019 20574
rect 18505 20634 18571 20637
rect 19425 20634 19491 20637
rect 18505 20632 19491 20634
rect 18505 20576 18510 20632
rect 18566 20576 19430 20632
rect 19486 20576 19491 20632
rect 18505 20574 19491 20576
rect 18505 20571 18571 20574
rect 19425 20571 19491 20574
rect 19977 20634 20043 20637
rect 23933 20634 23999 20637
rect 19977 20632 23999 20634
rect 19977 20576 19982 20632
rect 20038 20576 23938 20632
rect 23994 20576 23999 20632
rect 19977 20574 23999 20576
rect 19977 20571 20043 20574
rect 23933 20571 23999 20574
rect 200 20498 800 20528
rect 4061 20498 4127 20501
rect 200 20496 4127 20498
rect 200 20440 4066 20496
rect 4122 20440 4127 20496
rect 200 20438 4127 20440
rect 200 20408 800 20438
rect 4061 20435 4127 20438
rect 7557 20498 7623 20501
rect 13537 20498 13603 20501
rect 7557 20496 13603 20498
rect 7557 20440 7562 20496
rect 7618 20440 13542 20496
rect 13598 20440 13603 20496
rect 7557 20438 13603 20440
rect 7557 20435 7623 20438
rect 13537 20435 13603 20438
rect 13721 20498 13787 20501
rect 20478 20498 20484 20500
rect 13721 20496 20484 20498
rect 13721 20440 13726 20496
rect 13782 20440 20484 20496
rect 13721 20438 20484 20440
rect 13721 20435 13787 20438
rect 20478 20436 20484 20438
rect 20548 20498 20554 20500
rect 20621 20498 20687 20501
rect 20548 20496 20687 20498
rect 20548 20440 20626 20496
rect 20682 20440 20687 20496
rect 20548 20438 20687 20440
rect 20548 20436 20554 20438
rect 20621 20435 20687 20438
rect 21817 20498 21883 20501
rect 22461 20498 22527 20501
rect 22921 20498 22987 20501
rect 21817 20496 22527 20498
rect 21817 20440 21822 20496
rect 21878 20440 22466 20496
rect 22522 20440 22527 20496
rect 21817 20438 22527 20440
rect 21817 20435 21883 20438
rect 22461 20435 22527 20438
rect 22694 20496 22987 20498
rect 22694 20440 22926 20496
rect 22982 20440 22987 20496
rect 22694 20438 22987 20440
rect 6862 20300 6868 20364
rect 6932 20362 6938 20364
rect 8661 20362 8727 20365
rect 6932 20360 8727 20362
rect 6932 20304 8666 20360
rect 8722 20304 8727 20360
rect 6932 20302 8727 20304
rect 6932 20300 6938 20302
rect 8661 20299 8727 20302
rect 9673 20362 9739 20365
rect 11830 20362 11836 20364
rect 9673 20360 11836 20362
rect 9673 20304 9678 20360
rect 9734 20304 11836 20360
rect 9673 20302 11836 20304
rect 9673 20299 9739 20302
rect 11830 20300 11836 20302
rect 11900 20300 11906 20364
rect 11973 20362 12039 20365
rect 15377 20362 15443 20365
rect 11973 20360 15443 20362
rect 11973 20304 11978 20360
rect 12034 20304 15382 20360
rect 15438 20304 15443 20360
rect 11973 20302 15443 20304
rect 11973 20299 12039 20302
rect 15377 20299 15443 20302
rect 17350 20300 17356 20364
rect 17420 20362 17426 20364
rect 22369 20362 22435 20365
rect 17420 20360 22435 20362
rect 17420 20304 22374 20360
rect 22430 20304 22435 20360
rect 17420 20302 22435 20304
rect 17420 20300 17426 20302
rect 22369 20299 22435 20302
rect 22553 20362 22619 20365
rect 22694 20362 22754 20438
rect 22921 20435 22987 20438
rect 24117 20498 24183 20501
rect 27889 20498 27955 20501
rect 24117 20496 27955 20498
rect 24117 20440 24122 20496
rect 24178 20440 27894 20496
rect 27950 20440 27955 20496
rect 24117 20438 27955 20440
rect 24117 20435 24183 20438
rect 27889 20435 27955 20438
rect 22553 20360 22754 20362
rect 22553 20304 22558 20360
rect 22614 20304 22754 20360
rect 22553 20302 22754 20304
rect 24301 20362 24367 20365
rect 25957 20362 26023 20365
rect 24301 20360 26023 20362
rect 24301 20304 24306 20360
rect 24362 20304 25962 20360
rect 26018 20304 26023 20360
rect 24301 20302 26023 20304
rect 22553 20299 22619 20302
rect 24301 20299 24367 20302
rect 25957 20299 26023 20302
rect 6453 20228 6519 20229
rect 6453 20224 6500 20228
rect 6564 20226 6570 20228
rect 6453 20168 6458 20224
rect 6453 20164 6500 20168
rect 6564 20166 6610 20226
rect 6564 20164 6570 20166
rect 6862 20164 6868 20228
rect 6932 20226 6938 20228
rect 27102 20226 27108 20228
rect 6932 20166 27108 20226
rect 6932 20164 6938 20166
rect 27102 20164 27108 20166
rect 27172 20164 27178 20228
rect 6453 20163 6519 20164
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 6637 20090 6703 20093
rect 20662 20090 20668 20092
rect 6637 20088 20668 20090
rect 6637 20032 6642 20088
rect 6698 20032 20668 20088
rect 6637 20030 20668 20032
rect 6637 20027 6703 20030
rect 20662 20028 20668 20030
rect 20732 20028 20738 20092
rect 21357 20090 21423 20093
rect 26049 20090 26115 20093
rect 21357 20088 26115 20090
rect 21357 20032 21362 20088
rect 21418 20032 26054 20088
rect 26110 20032 26115 20088
rect 21357 20030 26115 20032
rect 21357 20027 21423 20030
rect 26049 20027 26115 20030
rect 3693 19954 3759 19957
rect 9581 19954 9647 19957
rect 3693 19952 9647 19954
rect 3693 19896 3698 19952
rect 3754 19896 9586 19952
rect 9642 19896 9647 19952
rect 3693 19894 9647 19896
rect 3693 19891 3759 19894
rect 9581 19891 9647 19894
rect 10593 19954 10659 19957
rect 13077 19954 13143 19957
rect 10593 19952 13143 19954
rect 10593 19896 10598 19952
rect 10654 19896 13082 19952
rect 13138 19896 13143 19952
rect 10593 19894 13143 19896
rect 10593 19891 10659 19894
rect 13077 19891 13143 19894
rect 13813 19954 13879 19957
rect 16021 19954 16087 19957
rect 18413 19954 18479 19957
rect 13813 19952 16087 19954
rect 13813 19896 13818 19952
rect 13874 19896 16026 19952
rect 16082 19896 16087 19952
rect 13813 19894 16087 19896
rect 13813 19891 13879 19894
rect 16021 19891 16087 19894
rect 16254 19952 18479 19954
rect 16254 19896 18418 19952
rect 18474 19896 18479 19952
rect 16254 19894 18479 19896
rect 13 19818 79 19821
rect 200 19818 800 19848
rect 4889 19820 4955 19821
rect 4838 19818 4844 19820
rect 13 19816 800 19818
rect 13 19760 18 19816
rect 74 19760 800 19816
rect 13 19758 800 19760
rect 4798 19758 4844 19818
rect 4908 19816 4955 19820
rect 4950 19760 4955 19816
rect 13 19755 79 19758
rect 200 19728 800 19758
rect 4838 19756 4844 19758
rect 4908 19756 4955 19760
rect 7782 19756 7788 19820
rect 7852 19818 7858 19820
rect 9489 19818 9555 19821
rect 10225 19820 10291 19821
rect 10174 19818 10180 19820
rect 7852 19816 9555 19818
rect 7852 19760 9494 19816
rect 9550 19760 9555 19816
rect 7852 19758 9555 19760
rect 10134 19758 10180 19818
rect 10244 19816 10291 19820
rect 10286 19760 10291 19816
rect 7852 19756 7858 19758
rect 4889 19755 4955 19756
rect 9489 19755 9555 19758
rect 10174 19756 10180 19758
rect 10244 19756 10291 19760
rect 12382 19756 12388 19820
rect 12452 19818 12458 19820
rect 12525 19818 12591 19821
rect 12452 19816 12591 19818
rect 12452 19760 12530 19816
rect 12586 19760 12591 19816
rect 12452 19758 12591 19760
rect 12452 19756 12458 19758
rect 10225 19755 10291 19756
rect 12525 19755 12591 19758
rect 12893 19818 12959 19821
rect 16254 19818 16314 19894
rect 18413 19891 18479 19894
rect 18822 19892 18828 19956
rect 18892 19954 18898 19956
rect 20437 19954 20503 19957
rect 18892 19952 20503 19954
rect 18892 19896 20442 19952
rect 20498 19896 20503 19952
rect 18892 19894 20503 19896
rect 18892 19892 18898 19894
rect 20437 19891 20503 19894
rect 22369 19954 22435 19957
rect 27705 19954 27771 19957
rect 22369 19952 27771 19954
rect 22369 19896 22374 19952
rect 22430 19896 27710 19952
rect 27766 19896 27771 19952
rect 22369 19894 27771 19896
rect 22369 19891 22435 19894
rect 27705 19891 27771 19894
rect 12893 19816 16314 19818
rect 12893 19760 12898 19816
rect 12954 19760 16314 19816
rect 12893 19758 16314 19760
rect 16389 19818 16455 19821
rect 19241 19818 19307 19821
rect 16389 19816 19307 19818
rect 16389 19760 16394 19816
rect 16450 19760 19246 19816
rect 19302 19760 19307 19816
rect 16389 19758 19307 19760
rect 12893 19755 12959 19758
rect 16389 19755 16455 19758
rect 19241 19755 19307 19758
rect 19701 19818 19767 19821
rect 20161 19820 20227 19821
rect 19701 19816 20040 19818
rect 19701 19760 19706 19816
rect 19762 19760 20040 19816
rect 19701 19758 20040 19760
rect 19701 19755 19767 19758
rect 5349 19682 5415 19685
rect 18229 19682 18295 19685
rect 5349 19680 18295 19682
rect 5349 19624 5354 19680
rect 5410 19624 18234 19680
rect 18290 19624 18295 19680
rect 5349 19622 18295 19624
rect 5349 19619 5415 19622
rect 18229 19619 18295 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 6361 19546 6427 19549
rect 11329 19546 11395 19549
rect 6361 19544 11395 19546
rect 6361 19488 6366 19544
rect 6422 19488 11334 19544
rect 11390 19488 11395 19544
rect 6361 19486 11395 19488
rect 6361 19483 6427 19486
rect 11329 19483 11395 19486
rect 11605 19546 11671 19549
rect 14089 19546 14155 19549
rect 11605 19544 14155 19546
rect 11605 19488 11610 19544
rect 11666 19488 14094 19544
rect 14150 19488 14155 19544
rect 11605 19486 14155 19488
rect 11605 19483 11671 19486
rect 14089 19483 14155 19486
rect 14825 19546 14891 19549
rect 15193 19546 15259 19549
rect 16297 19546 16363 19549
rect 14825 19544 16363 19546
rect 14825 19488 14830 19544
rect 14886 19488 15198 19544
rect 15254 19488 16302 19544
rect 16358 19488 16363 19544
rect 14825 19486 16363 19488
rect 14825 19483 14891 19486
rect 15193 19483 15259 19486
rect 16297 19483 16363 19486
rect 16941 19546 17007 19549
rect 19425 19546 19491 19549
rect 16941 19544 19491 19546
rect 16941 19488 16946 19544
rect 17002 19488 19430 19544
rect 19486 19488 19491 19544
rect 16941 19486 19491 19488
rect 19980 19546 20040 19758
rect 20110 19756 20116 19820
rect 20180 19818 20227 19820
rect 20180 19816 20272 19818
rect 20222 19760 20272 19816
rect 20180 19758 20272 19760
rect 20180 19756 20227 19758
rect 20662 19756 20668 19820
rect 20732 19818 20738 19820
rect 26233 19818 26299 19821
rect 20732 19816 26299 19818
rect 20732 19760 26238 19816
rect 26294 19760 26299 19816
rect 20732 19758 26299 19760
rect 20732 19756 20738 19758
rect 20161 19755 20227 19756
rect 26233 19755 26299 19758
rect 38285 19818 38351 19821
rect 39200 19818 39800 19848
rect 38285 19816 39800 19818
rect 38285 19760 38290 19816
rect 38346 19760 39800 19816
rect 38285 19758 39800 19760
rect 38285 19755 38351 19758
rect 39200 19728 39800 19758
rect 20110 19620 20116 19684
rect 20180 19682 20186 19684
rect 21633 19682 21699 19685
rect 25405 19682 25471 19685
rect 20180 19680 25471 19682
rect 20180 19624 21638 19680
rect 21694 19624 25410 19680
rect 25466 19624 25471 19680
rect 20180 19622 25471 19624
rect 20180 19620 20186 19622
rect 21633 19619 21699 19622
rect 25405 19619 25471 19622
rect 27061 19546 27127 19549
rect 19980 19544 27127 19546
rect 19980 19488 27066 19544
rect 27122 19488 27127 19544
rect 19980 19486 27127 19488
rect 16941 19483 17007 19486
rect 19425 19483 19491 19486
rect 27061 19483 27127 19486
rect 2865 19412 2931 19413
rect 2814 19348 2820 19412
rect 2884 19410 2931 19412
rect 2884 19408 2976 19410
rect 2926 19352 2976 19408
rect 2884 19350 2976 19352
rect 2884 19348 2931 19350
rect 4654 19348 4660 19412
rect 4724 19410 4730 19412
rect 4797 19410 4863 19413
rect 4724 19408 4863 19410
rect 4724 19352 4802 19408
rect 4858 19352 4863 19408
rect 4724 19350 4863 19352
rect 4724 19348 4730 19350
rect 2865 19347 2931 19348
rect 4797 19347 4863 19350
rect 7649 19410 7715 19413
rect 9029 19410 9095 19413
rect 7649 19408 9095 19410
rect 7649 19352 7654 19408
rect 7710 19352 9034 19408
rect 9090 19352 9095 19408
rect 7649 19350 9095 19352
rect 7649 19347 7715 19350
rect 9029 19347 9095 19350
rect 9949 19410 10015 19413
rect 11329 19410 11395 19413
rect 13721 19410 13787 19413
rect 9949 19408 10932 19410
rect 9949 19352 9954 19408
rect 10010 19353 10932 19408
rect 11329 19408 13787 19410
rect 10010 19352 10935 19353
rect 9949 19350 10935 19352
rect 9949 19347 10015 19350
rect 10869 19348 10935 19350
rect 10869 19292 10874 19348
rect 10930 19292 10935 19348
rect 11329 19352 11334 19408
rect 11390 19352 13726 19408
rect 13782 19352 13787 19408
rect 11329 19350 13787 19352
rect 11329 19347 11395 19350
rect 13721 19347 13787 19350
rect 14089 19410 14155 19413
rect 16665 19410 16731 19413
rect 14089 19408 16731 19410
rect 14089 19352 14094 19408
rect 14150 19352 16670 19408
rect 16726 19352 16731 19408
rect 14089 19350 16731 19352
rect 14089 19347 14155 19350
rect 16665 19347 16731 19350
rect 17309 19410 17375 19413
rect 17585 19410 17651 19413
rect 18137 19410 18203 19413
rect 20110 19410 20116 19412
rect 17309 19408 18203 19410
rect 17309 19352 17314 19408
rect 17370 19352 17590 19408
rect 17646 19352 18142 19408
rect 18198 19352 18203 19408
rect 17309 19350 18203 19352
rect 17309 19347 17375 19350
rect 17585 19347 17651 19350
rect 18137 19347 18203 19350
rect 19014 19350 20116 19410
rect 10869 19287 10935 19292
rect 7097 19274 7163 19277
rect 7741 19274 7807 19277
rect 7097 19272 7807 19274
rect 7097 19216 7102 19272
rect 7158 19216 7746 19272
rect 7802 19216 7807 19272
rect 7097 19214 7807 19216
rect 7097 19211 7163 19214
rect 7741 19211 7807 19214
rect 9581 19274 9647 19277
rect 9990 19274 9996 19276
rect 9581 19272 9996 19274
rect 9581 19216 9586 19272
rect 9642 19216 9996 19272
rect 9581 19214 9996 19216
rect 9581 19211 9647 19214
rect 9990 19212 9996 19214
rect 10060 19212 10066 19276
rect 11145 19274 11211 19277
rect 18689 19274 18755 19277
rect 11145 19272 18755 19274
rect 11145 19216 11150 19272
rect 11206 19216 18694 19272
rect 18750 19216 18755 19272
rect 11145 19214 18755 19216
rect 11145 19211 11211 19214
rect 18689 19211 18755 19214
rect 8201 19138 8267 19141
rect 11646 19138 11652 19140
rect 8201 19136 11652 19138
rect 8201 19080 8206 19136
rect 8262 19080 11652 19136
rect 8201 19078 11652 19080
rect 8201 19075 8267 19078
rect 11646 19076 11652 19078
rect 11716 19076 11722 19140
rect 11881 19138 11947 19141
rect 19014 19138 19074 19350
rect 20110 19348 20116 19350
rect 20180 19348 20186 19412
rect 25037 19410 25103 19413
rect 20302 19408 25103 19410
rect 20302 19352 25042 19408
rect 25098 19352 25103 19408
rect 20302 19350 25103 19352
rect 19149 19274 19215 19277
rect 20302 19274 20362 19350
rect 25037 19347 25103 19350
rect 26049 19410 26115 19413
rect 27613 19410 27679 19413
rect 26049 19408 27679 19410
rect 26049 19352 26054 19408
rect 26110 19352 27618 19408
rect 27674 19352 27679 19408
rect 26049 19350 27679 19352
rect 26049 19347 26115 19350
rect 27613 19347 27679 19350
rect 19149 19272 20362 19274
rect 19149 19216 19154 19272
rect 19210 19216 20362 19272
rect 19149 19214 20362 19216
rect 20621 19274 20687 19277
rect 26785 19274 26851 19277
rect 20621 19272 26851 19274
rect 20621 19216 20626 19272
rect 20682 19216 26790 19272
rect 26846 19216 26851 19272
rect 20621 19214 26851 19216
rect 19149 19211 19215 19214
rect 20621 19211 20687 19214
rect 26785 19211 26851 19214
rect 11881 19136 19074 19138
rect 11881 19080 11886 19136
rect 11942 19080 19074 19136
rect 11881 19078 19074 19080
rect 19149 19138 19215 19141
rect 20437 19138 20503 19141
rect 27061 19138 27127 19141
rect 19149 19136 20362 19138
rect 19149 19080 19154 19136
rect 19210 19080 20362 19136
rect 19149 19078 20362 19080
rect 11881 19075 11947 19078
rect 19149 19075 19215 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 9254 18940 9260 19004
rect 9324 19002 9330 19004
rect 9489 19002 9555 19005
rect 9324 19000 9555 19002
rect 9324 18944 9494 19000
rect 9550 18944 9555 19000
rect 9324 18942 9555 18944
rect 9324 18940 9330 18942
rect 9489 18939 9555 18942
rect 10358 18940 10364 19004
rect 10428 19002 10434 19004
rect 10910 19002 10916 19004
rect 10428 18942 10916 19002
rect 10428 18940 10434 18942
rect 10910 18940 10916 18942
rect 10980 18940 10986 19004
rect 11053 19002 11119 19005
rect 18781 19002 18847 19005
rect 11053 19000 18847 19002
rect 11053 18944 11058 19000
rect 11114 18944 18786 19000
rect 18842 18944 18847 19000
rect 11053 18942 18847 18944
rect 11053 18939 11119 18942
rect 18781 18939 18847 18942
rect 19333 19002 19399 19005
rect 20161 19002 20227 19005
rect 19333 19000 20227 19002
rect 19333 18944 19338 19000
rect 19394 18944 20166 19000
rect 20222 18944 20227 19000
rect 19333 18942 20227 18944
rect 20302 19002 20362 19078
rect 20437 19136 27127 19138
rect 20437 19080 20442 19136
rect 20498 19080 27066 19136
rect 27122 19080 27127 19136
rect 20437 19078 27127 19080
rect 20437 19075 20503 19078
rect 27061 19075 27127 19078
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19168
rect 34930 19007 35246 19008
rect 26141 19002 26207 19005
rect 20302 19000 26207 19002
rect 20302 18944 26146 19000
rect 26202 18944 26207 19000
rect 20302 18942 26207 18944
rect 19333 18939 19399 18942
rect 20161 18939 20227 18942
rect 26141 18939 26207 18942
rect 6269 18866 6335 18869
rect 10133 18866 10199 18869
rect 6269 18864 10199 18866
rect 6269 18808 6274 18864
rect 6330 18808 10138 18864
rect 10194 18808 10199 18864
rect 6269 18806 10199 18808
rect 6269 18803 6335 18806
rect 10133 18803 10199 18806
rect 10910 18804 10916 18868
rect 10980 18866 10986 18868
rect 11881 18866 11947 18869
rect 10980 18864 11947 18866
rect 10980 18808 11886 18864
rect 11942 18808 11947 18864
rect 10980 18806 11947 18808
rect 10980 18804 10986 18806
rect 11881 18803 11947 18806
rect 12065 18866 12131 18869
rect 12893 18866 12959 18869
rect 12065 18864 12959 18866
rect 12065 18808 12070 18864
rect 12126 18808 12898 18864
rect 12954 18808 12959 18864
rect 12065 18806 12959 18808
rect 12065 18803 12131 18806
rect 12893 18803 12959 18806
rect 13353 18866 13419 18869
rect 20345 18866 20411 18869
rect 20897 18866 20963 18869
rect 13353 18864 20963 18866
rect 13353 18808 13358 18864
rect 13414 18808 20350 18864
rect 20406 18808 20902 18864
rect 20958 18808 20963 18864
rect 13353 18806 20963 18808
rect 13353 18803 13419 18806
rect 20345 18803 20411 18806
rect 20897 18803 20963 18806
rect 21909 18866 21975 18869
rect 24301 18866 24367 18869
rect 21909 18864 24367 18866
rect 21909 18808 21914 18864
rect 21970 18808 24306 18864
rect 24362 18808 24367 18864
rect 21909 18806 24367 18808
rect 21909 18803 21975 18806
rect 24301 18803 24367 18806
rect 5349 18730 5415 18733
rect 17718 18730 17724 18732
rect 5349 18728 17724 18730
rect 5349 18672 5354 18728
rect 5410 18672 17724 18728
rect 5349 18670 17724 18672
rect 5349 18667 5415 18670
rect 17718 18668 17724 18670
rect 17788 18668 17794 18732
rect 17953 18730 18019 18733
rect 18965 18730 19031 18733
rect 20253 18730 20319 18733
rect 25681 18730 25747 18733
rect 17953 18728 19031 18730
rect 17953 18672 17958 18728
rect 18014 18672 18970 18728
rect 19026 18672 19031 18728
rect 17953 18670 19031 18672
rect 17953 18667 18019 18670
rect 18965 18667 19031 18670
rect 19382 18670 20178 18730
rect 4705 18594 4771 18597
rect 9213 18594 9279 18597
rect 4705 18592 9279 18594
rect 4705 18536 4710 18592
rect 4766 18536 9218 18592
rect 9274 18536 9279 18592
rect 4705 18534 9279 18536
rect 4705 18531 4771 18534
rect 9213 18531 9279 18534
rect 9857 18594 9923 18597
rect 11881 18594 11947 18597
rect 9857 18592 11947 18594
rect 9857 18536 9862 18592
rect 9918 18536 11886 18592
rect 11942 18536 11947 18592
rect 9857 18534 11947 18536
rect 9857 18531 9923 18534
rect 11881 18531 11947 18534
rect 12014 18532 12020 18596
rect 12084 18594 12090 18596
rect 13353 18594 13419 18597
rect 12084 18592 13419 18594
rect 12084 18536 13358 18592
rect 13414 18536 13419 18592
rect 12084 18534 13419 18536
rect 12084 18532 12090 18534
rect 13353 18531 13419 18534
rect 13905 18594 13971 18597
rect 15469 18594 15535 18597
rect 13905 18592 15535 18594
rect 13905 18536 13910 18592
rect 13966 18536 15474 18592
rect 15530 18536 15535 18592
rect 13905 18534 15535 18536
rect 13905 18531 13971 18534
rect 15469 18531 15535 18534
rect 16113 18594 16179 18597
rect 19149 18594 19215 18597
rect 16113 18592 19215 18594
rect 16113 18536 16118 18592
rect 16174 18536 19154 18592
rect 19210 18536 19215 18592
rect 16113 18534 19215 18536
rect 16113 18531 16179 18534
rect 19149 18531 19215 18534
rect 200 18458 800 18488
rect 1761 18458 1827 18461
rect 200 18456 1827 18458
rect 200 18400 1766 18456
rect 1822 18400 1827 18456
rect 200 18398 1827 18400
rect 200 18368 800 18398
rect 1761 18395 1827 18398
rect 8661 18458 8727 18461
rect 12065 18458 12131 18461
rect 8661 18456 12131 18458
rect 8661 18400 8666 18456
rect 8722 18400 12070 18456
rect 12126 18400 12131 18456
rect 8661 18398 12131 18400
rect 8661 18395 8727 18398
rect 12065 18395 12131 18398
rect 12341 18458 12407 18461
rect 14774 18458 14780 18460
rect 12341 18456 14780 18458
rect 12341 18400 12346 18456
rect 12402 18400 14780 18456
rect 12341 18398 14780 18400
rect 12341 18395 12407 18398
rect 14774 18396 14780 18398
rect 14844 18458 14850 18460
rect 19382 18458 19442 18670
rect 20118 18594 20178 18670
rect 20253 18728 25747 18730
rect 20253 18672 20258 18728
rect 20314 18672 25686 18728
rect 25742 18672 25747 18728
rect 20253 18670 25747 18672
rect 20253 18667 20319 18670
rect 25681 18667 25747 18670
rect 23841 18594 23907 18597
rect 20118 18592 23907 18594
rect 20118 18536 23846 18592
rect 23902 18536 23907 18592
rect 20118 18534 23907 18536
rect 23841 18531 23907 18534
rect 24669 18594 24735 18597
rect 26325 18594 26391 18597
rect 24669 18592 26391 18594
rect 24669 18536 24674 18592
rect 24730 18536 26330 18592
rect 26386 18536 26391 18592
rect 24669 18534 26391 18536
rect 24669 18531 24735 18534
rect 26325 18531 26391 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 14844 18398 19442 18458
rect 21633 18458 21699 18461
rect 27337 18458 27403 18461
rect 21633 18456 27403 18458
rect 21633 18400 21638 18456
rect 21694 18400 27342 18456
rect 27398 18400 27403 18456
rect 21633 18398 27403 18400
rect 14844 18396 14850 18398
rect 21633 18395 21699 18398
rect 27337 18395 27403 18398
rect 38285 18458 38351 18461
rect 39200 18458 39800 18488
rect 38285 18456 39800 18458
rect 38285 18400 38290 18456
rect 38346 18400 39800 18456
rect 38285 18398 39800 18400
rect 38285 18395 38351 18398
rect 39200 18368 39800 18398
rect 7414 18260 7420 18324
rect 7484 18322 7490 18324
rect 16389 18322 16455 18325
rect 7484 18320 16455 18322
rect 7484 18264 16394 18320
rect 16450 18264 16455 18320
rect 7484 18262 16455 18264
rect 7484 18260 7490 18262
rect 16389 18259 16455 18262
rect 17953 18322 18019 18325
rect 21030 18322 21036 18324
rect 17953 18320 21036 18322
rect 17953 18264 17958 18320
rect 18014 18264 21036 18320
rect 17953 18262 21036 18264
rect 17953 18259 18019 18262
rect 21030 18260 21036 18262
rect 21100 18260 21106 18324
rect 22134 18260 22140 18324
rect 22204 18322 22210 18324
rect 23565 18322 23631 18325
rect 27061 18322 27127 18325
rect 22204 18320 27127 18322
rect 22204 18264 23570 18320
rect 23626 18264 27066 18320
rect 27122 18264 27127 18320
rect 22204 18262 27127 18264
rect 22204 18260 22210 18262
rect 23565 18259 23631 18262
rect 27061 18259 27127 18262
rect 8569 18186 8635 18189
rect 8569 18184 9276 18186
rect 8569 18128 8574 18184
rect 8630 18128 9276 18184
rect 8569 18126 9276 18128
rect 8569 18123 8635 18126
rect 7833 18050 7899 18053
rect 8569 18050 8635 18053
rect 7833 18048 8635 18050
rect 7833 17992 7838 18048
rect 7894 17992 8574 18048
rect 8630 17992 8635 18048
rect 7833 17990 8635 17992
rect 7833 17987 7899 17990
rect 8569 17987 8635 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 7189 17914 7255 17917
rect 9029 17914 9095 17917
rect 7189 17912 9095 17914
rect 7189 17856 7194 17912
rect 7250 17856 9034 17912
rect 9090 17856 9095 17912
rect 7189 17854 9095 17856
rect 7189 17851 7255 17854
rect 9029 17851 9095 17854
rect 200 17778 800 17808
rect 4061 17778 4127 17781
rect 200 17776 4127 17778
rect 200 17720 4066 17776
rect 4122 17720 4127 17776
rect 200 17718 4127 17720
rect 200 17688 800 17718
rect 4061 17715 4127 17718
rect 6913 17778 6979 17781
rect 9216 17778 9276 18126
rect 9397 18184 9463 18189
rect 9397 18128 9402 18184
rect 9458 18128 9463 18184
rect 9397 18123 9463 18128
rect 10961 18186 11027 18189
rect 27245 18186 27311 18189
rect 29177 18186 29243 18189
rect 10961 18184 27311 18186
rect 10961 18128 10966 18184
rect 11022 18128 27250 18184
rect 27306 18128 27311 18184
rect 10961 18126 27311 18128
rect 10961 18123 11027 18126
rect 27245 18123 27311 18126
rect 29134 18184 29243 18186
rect 29134 18128 29182 18184
rect 29238 18128 29243 18184
rect 29134 18123 29243 18128
rect 29453 18186 29519 18189
rect 31293 18186 31359 18189
rect 29453 18184 31359 18186
rect 29453 18128 29458 18184
rect 29514 18128 31298 18184
rect 31354 18128 31359 18184
rect 29453 18126 31359 18128
rect 29453 18123 29519 18126
rect 31293 18123 31359 18126
rect 9400 18050 9460 18123
rect 13854 18050 13860 18052
rect 9400 17990 13860 18050
rect 13854 17988 13860 17990
rect 13924 17988 13930 18052
rect 14273 18050 14339 18053
rect 16798 18050 16804 18052
rect 14273 18048 16804 18050
rect 14273 17992 14278 18048
rect 14334 17992 16804 18048
rect 14273 17990 16804 17992
rect 14273 17987 14339 17990
rect 16798 17988 16804 17990
rect 16868 17988 16874 18052
rect 17166 17988 17172 18052
rect 17236 18050 17242 18052
rect 17769 18050 17835 18053
rect 17236 18048 17835 18050
rect 17236 17992 17774 18048
rect 17830 17992 17835 18048
rect 17236 17990 17835 17992
rect 17236 17988 17242 17990
rect 17769 17987 17835 17990
rect 18505 18050 18571 18053
rect 28809 18050 28875 18053
rect 18505 18048 28875 18050
rect 18505 17992 18510 18048
rect 18566 17992 28814 18048
rect 28870 17992 28875 18048
rect 18505 17990 28875 17992
rect 18505 17987 18571 17990
rect 28809 17987 28875 17990
rect 29134 17917 29194 18123
rect 29269 18050 29335 18053
rect 30833 18050 30899 18053
rect 29269 18048 30899 18050
rect 29269 17992 29274 18048
rect 29330 17992 30838 18048
rect 30894 17992 30899 18048
rect 29269 17990 30899 17992
rect 29269 17987 29335 17990
rect 30833 17987 30899 17990
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 10542 17852 10548 17916
rect 10612 17914 10618 17916
rect 10869 17914 10935 17917
rect 10612 17912 10935 17914
rect 10612 17856 10874 17912
rect 10930 17856 10935 17912
rect 10612 17854 10935 17856
rect 10612 17852 10618 17854
rect 10869 17851 10935 17854
rect 11237 17914 11303 17917
rect 11697 17914 11763 17917
rect 12433 17914 12499 17917
rect 11237 17912 11763 17914
rect 11237 17856 11242 17912
rect 11298 17856 11702 17912
rect 11758 17856 11763 17912
rect 11237 17854 11763 17856
rect 11237 17851 11303 17854
rect 11697 17851 11763 17854
rect 12390 17912 12499 17914
rect 12390 17856 12438 17912
rect 12494 17856 12499 17912
rect 12390 17851 12499 17856
rect 14089 17914 14155 17917
rect 16062 17914 16068 17916
rect 14089 17912 16068 17914
rect 14089 17856 14094 17912
rect 14150 17856 16068 17912
rect 14089 17854 16068 17856
rect 14089 17851 14155 17854
rect 16062 17852 16068 17854
rect 16132 17914 16138 17916
rect 16132 17854 20408 17914
rect 16132 17852 16138 17854
rect 12390 17778 12450 17851
rect 6913 17776 9138 17778
rect 6913 17720 6918 17776
rect 6974 17720 9138 17776
rect 6913 17718 9138 17720
rect 9216 17718 12450 17778
rect 13353 17778 13419 17781
rect 16113 17778 16179 17781
rect 13353 17776 16179 17778
rect 13353 17720 13358 17776
rect 13414 17720 16118 17776
rect 16174 17720 16179 17776
rect 13353 17718 16179 17720
rect 6913 17715 6979 17718
rect 6913 17642 6979 17645
rect 8886 17642 8892 17644
rect 6913 17640 8892 17642
rect 6913 17584 6918 17640
rect 6974 17584 8892 17640
rect 6913 17582 8892 17584
rect 6913 17579 6979 17582
rect 8886 17580 8892 17582
rect 8956 17580 8962 17644
rect 9078 17642 9138 17718
rect 13353 17715 13419 17718
rect 16113 17715 16179 17718
rect 16573 17778 16639 17781
rect 16982 17778 16988 17780
rect 16573 17776 16988 17778
rect 16573 17720 16578 17776
rect 16634 17720 16988 17776
rect 16573 17718 16988 17720
rect 16573 17715 16639 17718
rect 16982 17716 16988 17718
rect 17052 17716 17058 17780
rect 17125 17778 17191 17781
rect 20110 17778 20116 17780
rect 17125 17776 20116 17778
rect 17125 17720 17130 17776
rect 17186 17720 20116 17776
rect 17125 17718 20116 17720
rect 17125 17715 17191 17718
rect 20110 17716 20116 17718
rect 20180 17716 20186 17780
rect 20348 17778 20408 17854
rect 21214 17852 21220 17916
rect 21284 17914 21290 17916
rect 22829 17914 22895 17917
rect 21284 17912 22895 17914
rect 21284 17856 22834 17912
rect 22890 17856 22895 17912
rect 21284 17854 22895 17856
rect 21284 17852 21290 17854
rect 22829 17851 22895 17854
rect 23013 17914 23079 17917
rect 27245 17914 27311 17917
rect 23013 17912 27311 17914
rect 23013 17856 23018 17912
rect 23074 17856 27250 17912
rect 27306 17856 27311 17912
rect 23013 17854 27311 17856
rect 29134 17912 29243 17917
rect 29134 17856 29182 17912
rect 29238 17856 29243 17912
rect 29134 17854 29243 17856
rect 23013 17851 23079 17854
rect 27245 17851 27311 17854
rect 29177 17851 29243 17854
rect 23841 17778 23907 17781
rect 20348 17776 23907 17778
rect 20348 17720 23846 17776
rect 23902 17720 23907 17776
rect 20348 17718 23907 17720
rect 23841 17715 23907 17718
rect 25405 17778 25471 17781
rect 26366 17778 26372 17780
rect 25405 17776 26372 17778
rect 25405 17720 25410 17776
rect 25466 17720 26372 17776
rect 25405 17718 26372 17720
rect 25405 17715 25471 17718
rect 26366 17716 26372 17718
rect 26436 17716 26442 17780
rect 12157 17642 12223 17645
rect 28717 17642 28783 17645
rect 9078 17582 12082 17642
rect 12022 17509 12082 17582
rect 12157 17640 28783 17642
rect 12157 17584 12162 17640
rect 12218 17584 28722 17640
rect 28778 17584 28783 17640
rect 12157 17582 28783 17584
rect 12157 17579 12223 17582
rect 28717 17579 28783 17582
rect 7598 17444 7604 17508
rect 7668 17506 7674 17508
rect 11697 17506 11763 17509
rect 7668 17504 11763 17506
rect 7668 17448 11702 17504
rect 11758 17448 11763 17504
rect 7668 17446 11763 17448
rect 12022 17504 12131 17509
rect 12022 17448 12070 17504
rect 12126 17448 12131 17504
rect 12022 17446 12131 17448
rect 7668 17444 7674 17446
rect 11697 17443 11763 17446
rect 12065 17443 12131 17446
rect 12893 17506 12959 17509
rect 17125 17506 17191 17509
rect 12893 17504 17191 17506
rect 12893 17448 12898 17504
rect 12954 17448 17130 17504
rect 17186 17448 17191 17504
rect 12893 17446 17191 17448
rect 12893 17443 12959 17446
rect 17125 17443 17191 17446
rect 17534 17444 17540 17508
rect 17604 17506 17610 17508
rect 17953 17506 18019 17509
rect 17604 17504 18019 17506
rect 17604 17448 17958 17504
rect 18014 17448 18019 17504
rect 17604 17446 18019 17448
rect 17604 17444 17610 17446
rect 17953 17443 18019 17446
rect 19977 17506 20043 17509
rect 20161 17506 20227 17509
rect 19977 17504 20227 17506
rect 19977 17448 19982 17504
rect 20038 17448 20166 17504
rect 20222 17448 20227 17504
rect 19977 17446 20227 17448
rect 19977 17443 20043 17446
rect 20161 17443 20227 17446
rect 20437 17506 20503 17509
rect 21214 17506 21220 17508
rect 20437 17504 21220 17506
rect 20437 17448 20442 17504
rect 20498 17448 21220 17504
rect 20437 17446 21220 17448
rect 20437 17443 20503 17446
rect 21214 17444 21220 17446
rect 21284 17444 21290 17508
rect 21357 17506 21423 17509
rect 22134 17506 22140 17508
rect 21357 17504 22140 17506
rect 21357 17448 21362 17504
rect 21418 17448 22140 17504
rect 21357 17446 22140 17448
rect 21357 17443 21423 17446
rect 22134 17444 22140 17446
rect 22204 17444 22210 17508
rect 22318 17444 22324 17508
rect 22388 17506 22394 17508
rect 22553 17506 22619 17509
rect 22388 17504 22619 17506
rect 22388 17448 22558 17504
rect 22614 17448 22619 17504
rect 22388 17446 22619 17448
rect 22388 17444 22394 17446
rect 22553 17443 22619 17446
rect 22829 17506 22895 17509
rect 24945 17506 25011 17509
rect 22829 17504 25011 17506
rect 22829 17448 22834 17504
rect 22890 17448 24950 17504
rect 25006 17448 25011 17504
rect 22829 17446 25011 17448
rect 22829 17443 22895 17446
rect 24945 17443 25011 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 8569 17370 8635 17373
rect 9581 17370 9647 17373
rect 8569 17368 9647 17370
rect 8569 17312 8574 17368
rect 8630 17312 9586 17368
rect 9642 17312 9647 17368
rect 8569 17310 9647 17312
rect 8569 17307 8635 17310
rect 9581 17307 9647 17310
rect 10777 17370 10843 17373
rect 12893 17370 12959 17373
rect 10777 17368 12959 17370
rect 10777 17312 10782 17368
rect 10838 17312 12898 17368
rect 12954 17312 12959 17368
rect 10777 17310 12959 17312
rect 10777 17307 10843 17310
rect 12893 17307 12959 17310
rect 13721 17370 13787 17373
rect 13854 17370 13860 17372
rect 13721 17368 13860 17370
rect 13721 17312 13726 17368
rect 13782 17312 13860 17368
rect 13721 17310 13860 17312
rect 13721 17307 13787 17310
rect 13854 17308 13860 17310
rect 13924 17308 13930 17372
rect 14273 17370 14339 17373
rect 19977 17370 20043 17373
rect 22093 17370 22159 17373
rect 14273 17368 19350 17370
rect 14273 17312 14278 17368
rect 14334 17312 19350 17368
rect 14273 17310 19350 17312
rect 14273 17307 14339 17310
rect 4245 17234 4311 17237
rect 5993 17234 6059 17237
rect 11278 17234 11284 17236
rect 4245 17232 11284 17234
rect 4245 17176 4250 17232
rect 4306 17176 5998 17232
rect 6054 17176 11284 17232
rect 4245 17174 11284 17176
rect 4245 17171 4311 17174
rect 5993 17171 6059 17174
rect 11278 17172 11284 17174
rect 11348 17172 11354 17236
rect 11789 17234 11855 17237
rect 14089 17234 14155 17237
rect 11789 17232 14155 17234
rect 11789 17176 11794 17232
rect 11850 17176 14094 17232
rect 14150 17176 14155 17232
rect 11789 17174 14155 17176
rect 11789 17171 11855 17174
rect 14089 17171 14155 17174
rect 14365 17234 14431 17237
rect 18321 17236 18387 17237
rect 18270 17234 18276 17236
rect 14365 17232 17970 17234
rect 14365 17176 14370 17232
rect 14426 17176 17970 17232
rect 14365 17174 17970 17176
rect 18230 17174 18276 17234
rect 18340 17232 18387 17236
rect 18382 17176 18387 17232
rect 14365 17171 14431 17174
rect 200 17098 800 17128
rect 17910 17101 17970 17174
rect 18270 17172 18276 17174
rect 18340 17172 18387 17176
rect 18822 17172 18828 17236
rect 18892 17234 18898 17236
rect 19149 17234 19215 17237
rect 18892 17232 19215 17234
rect 18892 17176 19154 17232
rect 19210 17176 19215 17232
rect 18892 17174 19215 17176
rect 19290 17234 19350 17310
rect 19977 17368 22159 17370
rect 19977 17312 19982 17368
rect 20038 17312 22098 17368
rect 22154 17312 22159 17368
rect 19977 17310 22159 17312
rect 19977 17307 20043 17310
rect 22093 17307 22159 17310
rect 22277 17370 22343 17373
rect 24853 17370 24919 17373
rect 22277 17368 24919 17370
rect 22277 17312 22282 17368
rect 22338 17312 24858 17368
rect 24914 17312 24919 17368
rect 22277 17310 24919 17312
rect 22277 17307 22343 17310
rect 24853 17307 24919 17310
rect 19609 17234 19675 17237
rect 19290 17232 19675 17234
rect 19290 17176 19614 17232
rect 19670 17176 19675 17232
rect 19290 17174 19675 17176
rect 18892 17172 18898 17174
rect 18321 17171 18387 17172
rect 19149 17171 19215 17174
rect 19609 17171 19675 17174
rect 20345 17234 20411 17237
rect 20713 17234 20779 17237
rect 20345 17232 20779 17234
rect 20345 17176 20350 17232
rect 20406 17176 20718 17232
rect 20774 17176 20779 17232
rect 20345 17174 20779 17176
rect 20345 17171 20411 17174
rect 20713 17171 20779 17174
rect 21081 17234 21147 17237
rect 27705 17234 27771 17237
rect 21081 17232 27771 17234
rect 21081 17176 21086 17232
rect 21142 17176 27710 17232
rect 27766 17176 27771 17232
rect 21081 17174 27771 17176
rect 21081 17171 21147 17174
rect 27705 17171 27771 17174
rect 9857 17098 9923 17101
rect 200 17096 9923 17098
rect 200 17040 9862 17096
rect 9918 17040 9923 17096
rect 200 17038 9923 17040
rect 200 17008 800 17038
rect 9857 17035 9923 17038
rect 13261 17098 13327 17101
rect 17350 17098 17356 17100
rect 13261 17096 17356 17098
rect 13261 17040 13266 17096
rect 13322 17040 17356 17096
rect 13261 17038 17356 17040
rect 13261 17035 13327 17038
rect 17350 17036 17356 17038
rect 17420 17036 17426 17100
rect 17910 17098 18019 17101
rect 19006 17098 19012 17100
rect 17910 17096 19012 17098
rect 17910 17040 17958 17096
rect 18014 17040 19012 17096
rect 17910 17038 19012 17040
rect 17953 17035 18019 17038
rect 19006 17036 19012 17038
rect 19076 17036 19082 17100
rect 19333 17098 19399 17101
rect 21214 17098 21220 17100
rect 19333 17096 21220 17098
rect 19333 17040 19338 17096
rect 19394 17040 21220 17096
rect 19333 17038 21220 17040
rect 19333 17035 19399 17038
rect 21214 17036 21220 17038
rect 21284 17036 21290 17100
rect 21357 17098 21423 17101
rect 23289 17098 23355 17101
rect 21357 17096 23355 17098
rect 21357 17040 21362 17096
rect 21418 17040 23294 17096
rect 23350 17040 23355 17096
rect 21357 17038 23355 17040
rect 21357 17035 21423 17038
rect 23289 17035 23355 17038
rect 24945 17098 25011 17101
rect 27521 17098 27587 17101
rect 24945 17096 27587 17098
rect 24945 17040 24950 17096
rect 25006 17040 27526 17096
rect 27582 17040 27587 17096
rect 24945 17038 27587 17040
rect 24945 17035 25011 17038
rect 27521 17035 27587 17038
rect 37457 17098 37523 17101
rect 39200 17098 39800 17128
rect 37457 17096 39800 17098
rect 37457 17040 37462 17096
rect 37518 17040 39800 17096
rect 37457 17038 39800 17040
rect 37457 17035 37523 17038
rect 39200 17008 39800 17038
rect 12249 16962 12315 16965
rect 5260 16960 12315 16962
rect 5260 16904 12254 16960
rect 12310 16904 12315 16960
rect 5260 16902 12315 16904
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 2405 16690 2471 16693
rect 5260 16690 5320 16902
rect 12249 16899 12315 16902
rect 14181 16962 14247 16965
rect 28441 16962 28507 16965
rect 14181 16960 28507 16962
rect 14181 16904 14186 16960
rect 14242 16904 28446 16960
rect 28502 16904 28507 16960
rect 14181 16902 28507 16904
rect 14181 16899 14247 16902
rect 28441 16899 28507 16902
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 8201 16826 8267 16829
rect 14958 16826 14964 16828
rect 8201 16824 14964 16826
rect 8201 16768 8206 16824
rect 8262 16768 14964 16824
rect 8201 16766 14964 16768
rect 8201 16763 8267 16766
rect 14958 16764 14964 16766
rect 15028 16764 15034 16828
rect 15193 16826 15259 16829
rect 15469 16826 15535 16829
rect 15193 16824 15535 16826
rect 15193 16768 15198 16824
rect 15254 16768 15474 16824
rect 15530 16768 15535 16824
rect 15193 16766 15535 16768
rect 15193 16763 15259 16766
rect 15469 16763 15535 16766
rect 16941 16826 17007 16829
rect 19333 16826 19399 16829
rect 16941 16824 19399 16826
rect 16941 16768 16946 16824
rect 17002 16768 19338 16824
rect 19394 16768 19399 16824
rect 16941 16766 19399 16768
rect 16941 16763 17007 16766
rect 19333 16763 19399 16766
rect 19517 16826 19583 16829
rect 21357 16826 21423 16829
rect 19517 16824 21423 16826
rect 19517 16768 19522 16824
rect 19578 16768 21362 16824
rect 21418 16768 21423 16824
rect 19517 16766 21423 16768
rect 19517 16763 19583 16766
rect 21357 16763 21423 16766
rect 21725 16826 21791 16829
rect 22093 16826 22159 16829
rect 21725 16824 22159 16826
rect 21725 16768 21730 16824
rect 21786 16768 22098 16824
rect 22154 16768 22159 16824
rect 21725 16766 22159 16768
rect 21725 16763 21791 16766
rect 22093 16763 22159 16766
rect 22277 16826 22343 16829
rect 25037 16826 25103 16829
rect 27061 16826 27127 16829
rect 22277 16824 27127 16826
rect 22277 16768 22282 16824
rect 22338 16768 25042 16824
rect 25098 16768 27066 16824
rect 27122 16768 27127 16824
rect 22277 16766 27127 16768
rect 22277 16763 22343 16766
rect 25037 16763 25103 16766
rect 27061 16763 27127 16766
rect 2405 16688 5320 16690
rect 2405 16632 2410 16688
rect 2466 16632 5320 16688
rect 2405 16630 5320 16632
rect 5441 16690 5507 16693
rect 7230 16690 7236 16692
rect 5441 16688 7236 16690
rect 5441 16632 5446 16688
rect 5502 16632 7236 16688
rect 5441 16630 7236 16632
rect 2405 16627 2471 16630
rect 5441 16627 5507 16630
rect 7230 16628 7236 16630
rect 7300 16628 7306 16692
rect 8569 16690 8635 16693
rect 8702 16690 8708 16692
rect 8569 16688 8708 16690
rect 8569 16632 8574 16688
rect 8630 16632 8708 16688
rect 8569 16630 8708 16632
rect 8569 16627 8635 16630
rect 8702 16628 8708 16630
rect 8772 16628 8778 16692
rect 9121 16690 9187 16693
rect 9254 16690 9260 16692
rect 9121 16688 9260 16690
rect 9121 16632 9126 16688
rect 9182 16632 9260 16688
rect 9121 16630 9260 16632
rect 9121 16627 9187 16630
rect 9254 16628 9260 16630
rect 9324 16628 9330 16692
rect 12157 16690 12223 16693
rect 13261 16690 13327 16693
rect 12157 16688 13327 16690
rect 12157 16632 12162 16688
rect 12218 16632 13266 16688
rect 13322 16632 13327 16688
rect 12157 16630 13327 16632
rect 12157 16627 12223 16630
rect 13261 16627 13327 16630
rect 13905 16690 13971 16693
rect 18505 16690 18571 16693
rect 13905 16688 18571 16690
rect 13905 16632 13910 16688
rect 13966 16632 18510 16688
rect 18566 16632 18571 16688
rect 13905 16630 18571 16632
rect 13905 16627 13971 16630
rect 18505 16627 18571 16630
rect 18873 16690 18939 16693
rect 20161 16690 20227 16693
rect 18873 16688 20227 16690
rect 18873 16632 18878 16688
rect 18934 16632 20166 16688
rect 20222 16632 20227 16688
rect 18873 16630 20227 16632
rect 18873 16627 18939 16630
rect 20161 16627 20227 16630
rect 20478 16628 20484 16692
rect 20548 16690 20554 16692
rect 20621 16690 20687 16693
rect 20548 16688 20687 16690
rect 20548 16632 20626 16688
rect 20682 16632 20687 16688
rect 20548 16630 20687 16632
rect 20548 16628 20554 16630
rect 20621 16627 20687 16630
rect 20846 16628 20852 16692
rect 20916 16690 20922 16692
rect 22185 16690 22251 16693
rect 20916 16688 22251 16690
rect 20916 16632 22190 16688
rect 22246 16632 22251 16688
rect 20916 16630 22251 16632
rect 20916 16628 20922 16630
rect 22185 16627 22251 16630
rect 22921 16690 22987 16693
rect 25681 16690 25747 16693
rect 22921 16688 25747 16690
rect 22921 16632 22926 16688
rect 22982 16632 25686 16688
rect 25742 16632 25747 16688
rect 22921 16630 25747 16632
rect 22921 16627 22987 16630
rect 25681 16627 25747 16630
rect 3877 16554 3943 16557
rect 29085 16554 29151 16557
rect 3877 16552 29151 16554
rect 3877 16496 3882 16552
rect 3938 16496 29090 16552
rect 29146 16496 29151 16552
rect 3877 16494 29151 16496
rect 3877 16491 3943 16494
rect 29085 16491 29151 16494
rect 4061 16418 4127 16421
rect 6862 16418 6868 16420
rect 4061 16416 6868 16418
rect 4061 16360 4066 16416
rect 4122 16360 6868 16416
rect 4061 16358 6868 16360
rect 4061 16355 4127 16358
rect 6862 16356 6868 16358
rect 6932 16356 6938 16420
rect 8753 16418 8819 16421
rect 12065 16418 12131 16421
rect 8753 16416 12131 16418
rect 8753 16360 8758 16416
rect 8814 16360 12070 16416
rect 12126 16360 12131 16416
rect 8753 16358 12131 16360
rect 8753 16355 8819 16358
rect 12065 16355 12131 16358
rect 12382 16356 12388 16420
rect 12452 16418 12458 16420
rect 20437 16418 20503 16421
rect 28625 16418 28691 16421
rect 12452 16358 19488 16418
rect 12452 16356 12458 16358
rect 9070 16220 9076 16284
rect 9140 16282 9146 16284
rect 9489 16282 9555 16285
rect 9140 16280 9555 16282
rect 9140 16224 9494 16280
rect 9550 16224 9555 16280
rect 9140 16222 9555 16224
rect 9140 16220 9146 16222
rect 9489 16219 9555 16222
rect 10777 16282 10843 16285
rect 18873 16282 18939 16285
rect 10777 16280 18939 16282
rect 10777 16224 10782 16280
rect 10838 16224 18878 16280
rect 18934 16224 18939 16280
rect 10777 16222 18939 16224
rect 10777 16219 10843 16222
rect 18873 16219 18939 16222
rect 19057 16282 19123 16285
rect 19241 16282 19307 16285
rect 19057 16280 19307 16282
rect 19057 16224 19062 16280
rect 19118 16224 19246 16280
rect 19302 16224 19307 16280
rect 19057 16222 19307 16224
rect 19057 16219 19123 16222
rect 19241 16219 19307 16222
rect 19428 16180 19488 16358
rect 20437 16416 28691 16418
rect 20437 16360 20442 16416
rect 20498 16360 28630 16416
rect 28686 16360 28691 16416
rect 20437 16358 28691 16360
rect 20437 16355 20503 16358
rect 28625 16355 28691 16358
rect 38101 16418 38167 16421
rect 39200 16418 39800 16448
rect 38101 16416 39800 16418
rect 38101 16360 38106 16416
rect 38162 16360 39800 16416
rect 38101 16358 39800 16360
rect 38101 16355 38167 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 39200 16328 39800 16358
rect 19570 16287 19886 16288
rect 24117 16282 24183 16285
rect 19980 16280 24183 16282
rect 19980 16224 24122 16280
rect 24178 16224 24183 16280
rect 19980 16222 24183 16224
rect 19980 16180 20040 16222
rect 24117 16219 24183 16222
rect 6729 16146 6795 16149
rect 17033 16146 17099 16149
rect 6729 16144 17099 16146
rect 6729 16088 6734 16144
rect 6790 16088 17038 16144
rect 17094 16088 17099 16144
rect 6729 16086 17099 16088
rect 6729 16083 6795 16086
rect 17033 16083 17099 16086
rect 17585 16146 17651 16149
rect 17585 16144 19350 16146
rect 17585 16088 17590 16144
rect 17646 16088 19350 16144
rect 19428 16120 20040 16180
rect 20529 16146 20595 16149
rect 20846 16146 20852 16148
rect 20529 16144 20852 16146
rect 17585 16086 19350 16088
rect 17585 16083 17651 16086
rect 5165 16010 5231 16013
rect 19057 16010 19123 16013
rect 5165 16008 19123 16010
rect 5165 15952 5170 16008
rect 5226 15952 19062 16008
rect 19118 15952 19123 16008
rect 5165 15950 19123 15952
rect 19290 16010 19350 16086
rect 20529 16088 20534 16144
rect 20590 16088 20852 16144
rect 20529 16086 20852 16088
rect 20529 16083 20595 16086
rect 20846 16084 20852 16086
rect 20916 16084 20922 16148
rect 20989 16146 21055 16149
rect 21265 16146 21331 16149
rect 21541 16146 21607 16149
rect 26877 16146 26943 16149
rect 27429 16146 27495 16149
rect 20989 16144 21607 16146
rect 20989 16088 20994 16144
rect 21050 16088 21270 16144
rect 21326 16088 21546 16144
rect 21602 16088 21607 16144
rect 20989 16086 21607 16088
rect 20989 16083 21055 16086
rect 21265 16083 21331 16086
rect 21541 16083 21607 16086
rect 22924 16144 27495 16146
rect 22924 16088 26882 16144
rect 26938 16088 27434 16144
rect 27490 16088 27495 16144
rect 22924 16086 27495 16088
rect 22924 16010 22984 16086
rect 26877 16083 26943 16086
rect 27429 16083 27495 16086
rect 19290 15950 22984 16010
rect 23105 16010 23171 16013
rect 26969 16010 27035 16013
rect 23105 16008 27035 16010
rect 23105 15952 23110 16008
rect 23166 15952 26974 16008
rect 27030 15952 27035 16008
rect 23105 15950 27035 15952
rect 5165 15947 5231 15950
rect 19057 15947 19123 15950
rect 23105 15947 23171 15950
rect 26969 15947 27035 15950
rect 8845 15874 8911 15877
rect 12433 15874 12499 15877
rect 8845 15872 12499 15874
rect 8845 15816 8850 15872
rect 8906 15816 12438 15872
rect 12494 15816 12499 15872
rect 8845 15814 12499 15816
rect 8845 15811 8911 15814
rect 12433 15811 12499 15814
rect 12801 15874 12867 15877
rect 12801 15872 13508 15874
rect 12801 15816 12806 15872
rect 12862 15816 13508 15872
rect 12801 15814 13508 15816
rect 12801 15811 12867 15814
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 1669 15738 1735 15741
rect 200 15736 1735 15738
rect 200 15680 1674 15736
rect 1730 15680 1735 15736
rect 200 15678 1735 15680
rect 200 15648 800 15678
rect 1669 15675 1735 15678
rect 3233 15738 3299 15741
rect 3550 15738 3556 15740
rect 3233 15736 3556 15738
rect 3233 15680 3238 15736
rect 3294 15680 3556 15736
rect 3233 15678 3556 15680
rect 3233 15675 3299 15678
rect 3550 15676 3556 15678
rect 3620 15676 3626 15740
rect 11789 15738 11855 15741
rect 13261 15738 13327 15741
rect 11789 15736 13327 15738
rect 11789 15680 11794 15736
rect 11850 15680 13266 15736
rect 13322 15680 13327 15736
rect 11789 15678 13327 15680
rect 13448 15738 13508 15814
rect 13854 15812 13860 15876
rect 13924 15874 13930 15876
rect 14365 15874 14431 15877
rect 14590 15874 14596 15876
rect 13924 15872 14596 15874
rect 13924 15816 14370 15872
rect 14426 15816 14596 15872
rect 13924 15814 14596 15816
rect 13924 15812 13930 15814
rect 14365 15811 14431 15814
rect 14590 15812 14596 15814
rect 14660 15812 14666 15876
rect 15377 15874 15443 15877
rect 27153 15874 27219 15877
rect 15377 15872 27219 15874
rect 15377 15816 15382 15872
rect 15438 15816 27158 15872
rect 27214 15816 27219 15872
rect 15377 15814 27219 15816
rect 15377 15811 15443 15814
rect 27153 15811 27219 15814
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 16481 15738 16547 15741
rect 13448 15736 16547 15738
rect 13448 15680 16486 15736
rect 16542 15680 16547 15736
rect 13448 15678 16547 15680
rect 11789 15675 11855 15678
rect 13261 15675 13327 15678
rect 16481 15675 16547 15678
rect 17033 15738 17099 15741
rect 18137 15740 18203 15741
rect 17902 15738 17908 15740
rect 17033 15736 17908 15738
rect 17033 15680 17038 15736
rect 17094 15680 17908 15736
rect 17033 15678 17908 15680
rect 17033 15675 17099 15678
rect 17902 15676 17908 15678
rect 17972 15676 17978 15740
rect 18086 15676 18092 15740
rect 18156 15738 18203 15740
rect 19057 15738 19123 15741
rect 23105 15738 23171 15741
rect 24853 15740 24919 15741
rect 24853 15738 24900 15740
rect 18156 15736 18248 15738
rect 18198 15680 18248 15736
rect 18156 15678 18248 15680
rect 19057 15736 23171 15738
rect 19057 15680 19062 15736
rect 19118 15680 23110 15736
rect 23166 15680 23171 15736
rect 19057 15678 23171 15680
rect 24808 15736 24900 15738
rect 24808 15680 24858 15736
rect 24808 15678 24900 15680
rect 18156 15676 18203 15678
rect 18137 15675 18203 15676
rect 19057 15675 19123 15678
rect 23105 15675 23171 15678
rect 24853 15676 24900 15678
rect 24964 15676 24970 15740
rect 24853 15675 24919 15676
rect 11421 15602 11487 15605
rect 12801 15602 12867 15605
rect 11421 15600 12867 15602
rect 11421 15544 11426 15600
rect 11482 15544 12806 15600
rect 12862 15544 12867 15600
rect 11421 15542 12867 15544
rect 11421 15539 11487 15542
rect 12801 15539 12867 15542
rect 13169 15602 13235 15605
rect 16757 15602 16823 15605
rect 13169 15600 16823 15602
rect 13169 15544 13174 15600
rect 13230 15544 16762 15600
rect 16818 15544 16823 15600
rect 13169 15542 16823 15544
rect 13169 15539 13235 15542
rect 16757 15539 16823 15542
rect 17309 15602 17375 15605
rect 21541 15602 21607 15605
rect 17309 15600 21607 15602
rect 17309 15544 17314 15600
rect 17370 15544 21546 15600
rect 21602 15544 21607 15600
rect 17309 15542 21607 15544
rect 17309 15539 17375 15542
rect 21541 15539 21607 15542
rect 22737 15602 22803 15605
rect 25497 15602 25563 15605
rect 22737 15600 25563 15602
rect 22737 15544 22742 15600
rect 22798 15544 25502 15600
rect 25558 15544 25563 15600
rect 22737 15542 25563 15544
rect 22737 15539 22803 15542
rect 25497 15539 25563 15542
rect 7925 15466 7991 15469
rect 13077 15466 13143 15469
rect 7925 15464 13143 15466
rect 7925 15408 7930 15464
rect 7986 15408 13082 15464
rect 13138 15408 13143 15464
rect 7925 15406 13143 15408
rect 7925 15403 7991 15406
rect 13077 15403 13143 15406
rect 14774 15404 14780 15468
rect 14844 15466 14850 15468
rect 17350 15466 17356 15468
rect 14844 15406 17356 15466
rect 14844 15404 14850 15406
rect 17350 15404 17356 15406
rect 17420 15466 17426 15468
rect 17769 15466 17835 15469
rect 17420 15464 17835 15466
rect 17420 15408 17774 15464
rect 17830 15408 17835 15464
rect 17420 15406 17835 15408
rect 17420 15404 17426 15406
rect 17769 15403 17835 15406
rect 17902 15404 17908 15468
rect 17972 15466 17978 15468
rect 20621 15466 20687 15469
rect 17972 15464 20687 15466
rect 17972 15408 20626 15464
rect 20682 15408 20687 15464
rect 17972 15406 20687 15408
rect 17972 15404 17978 15406
rect 20621 15403 20687 15406
rect 20805 15466 20871 15469
rect 22461 15466 22527 15469
rect 20805 15464 22527 15466
rect 20805 15408 20810 15464
rect 20866 15408 22466 15464
rect 22522 15408 22527 15464
rect 20805 15406 22527 15408
rect 20805 15403 20871 15406
rect 22461 15403 22527 15406
rect 9673 15330 9739 15333
rect 10041 15330 10107 15333
rect 11697 15330 11763 15333
rect 12014 15330 12020 15332
rect 9673 15328 10107 15330
rect 9673 15272 9678 15328
rect 9734 15272 10046 15328
rect 10102 15272 10107 15328
rect 9673 15270 10107 15272
rect 9673 15267 9739 15270
rect 10041 15267 10107 15270
rect 10182 15328 12020 15330
rect 10182 15272 11702 15328
rect 11758 15272 12020 15328
rect 10182 15270 12020 15272
rect 7833 15196 7899 15197
rect 7782 15194 7788 15196
rect 7742 15134 7788 15194
rect 7852 15192 7899 15196
rect 7894 15136 7899 15192
rect 7782 15132 7788 15134
rect 7852 15132 7899 15136
rect 9438 15132 9444 15196
rect 9508 15194 9514 15196
rect 9581 15194 9647 15197
rect 9508 15192 9647 15194
rect 9508 15136 9586 15192
rect 9642 15136 9647 15192
rect 9508 15134 9647 15136
rect 9508 15132 9514 15134
rect 7833 15131 7899 15132
rect 9581 15131 9647 15134
rect 9857 15194 9923 15197
rect 10182 15194 10242 15270
rect 11697 15267 11763 15270
rect 12014 15268 12020 15270
rect 12084 15268 12090 15332
rect 12157 15330 12223 15333
rect 14641 15330 14707 15333
rect 12157 15328 14707 15330
rect 12157 15272 12162 15328
rect 12218 15272 14646 15328
rect 14702 15272 14707 15328
rect 12157 15270 14707 15272
rect 12157 15267 12223 15270
rect 14641 15267 14707 15270
rect 15009 15330 15075 15333
rect 18454 15330 18460 15332
rect 15009 15328 18460 15330
rect 15009 15272 15014 15328
rect 15070 15272 18460 15328
rect 15009 15270 18460 15272
rect 15009 15267 15075 15270
rect 18454 15268 18460 15270
rect 18524 15268 18530 15332
rect 20161 15330 20227 15333
rect 20897 15332 20963 15333
rect 20846 15330 20852 15332
rect 20161 15328 20362 15330
rect 20161 15272 20166 15328
rect 20222 15272 20362 15328
rect 20161 15270 20362 15272
rect 20806 15270 20852 15330
rect 20916 15328 20963 15332
rect 20958 15272 20963 15328
rect 20161 15267 20227 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 9857 15192 10242 15194
rect 9857 15136 9862 15192
rect 9918 15136 10242 15192
rect 9857 15134 10242 15136
rect 10961 15194 11027 15197
rect 12198 15194 12204 15196
rect 10961 15192 12204 15194
rect 10961 15136 10966 15192
rect 11022 15136 12204 15192
rect 10961 15134 12204 15136
rect 9857 15131 9923 15134
rect 10961 15131 11027 15134
rect 12198 15132 12204 15134
rect 12268 15132 12274 15196
rect 13721 15194 13787 15197
rect 18822 15194 18828 15196
rect 13721 15192 18828 15194
rect 13721 15136 13726 15192
rect 13782 15136 18828 15192
rect 13721 15134 18828 15136
rect 13721 15131 13787 15134
rect 18822 15132 18828 15134
rect 18892 15132 18898 15196
rect 19149 15194 19215 15197
rect 19425 15194 19491 15197
rect 19149 15192 19491 15194
rect 19149 15136 19154 15192
rect 19210 15136 19430 15192
rect 19486 15136 19491 15192
rect 19149 15134 19491 15136
rect 19149 15131 19215 15134
rect 19425 15131 19491 15134
rect 19977 15194 20043 15197
rect 20110 15194 20116 15196
rect 19977 15192 20116 15194
rect 19977 15136 19982 15192
rect 20038 15136 20116 15192
rect 19977 15134 20116 15136
rect 19977 15131 20043 15134
rect 20110 15132 20116 15134
rect 20180 15132 20186 15196
rect 20302 15194 20362 15270
rect 20846 15268 20852 15270
rect 20916 15268 20963 15272
rect 20897 15267 20963 15268
rect 23197 15194 23263 15197
rect 29085 15194 29151 15197
rect 20302 15192 23263 15194
rect 20302 15136 23202 15192
rect 23258 15136 23263 15192
rect 20302 15134 23263 15136
rect 23197 15131 23263 15134
rect 23430 15192 29151 15194
rect 23430 15136 29090 15192
rect 29146 15136 29151 15192
rect 23430 15134 29151 15136
rect 200 15058 800 15088
rect 3918 15058 3924 15060
rect 200 14998 3924 15058
rect 200 14968 800 14998
rect 3918 14996 3924 14998
rect 3988 14996 3994 15060
rect 6361 15058 6427 15061
rect 17309 15058 17375 15061
rect 21357 15058 21423 15061
rect 6361 15056 17234 15058
rect 6361 15000 6366 15056
rect 6422 15000 17234 15056
rect 6361 14998 17234 15000
rect 6361 14995 6427 14998
rect 8017 14922 8083 14925
rect 10726 14922 10732 14924
rect 8017 14920 10732 14922
rect 8017 14864 8022 14920
rect 8078 14864 10732 14920
rect 8017 14862 10732 14864
rect 8017 14859 8083 14862
rect 10726 14860 10732 14862
rect 10796 14860 10802 14924
rect 12065 14922 12131 14925
rect 17174 14922 17234 14998
rect 17309 15056 21423 15058
rect 17309 15000 17314 15056
rect 17370 15000 21362 15056
rect 21418 15000 21423 15056
rect 17309 14998 21423 15000
rect 17309 14995 17375 14998
rect 21357 14995 21423 14998
rect 21909 15058 21975 15061
rect 23430 15058 23490 15134
rect 29085 15131 29151 15134
rect 27337 15060 27403 15061
rect 21909 15056 23490 15058
rect 21909 15000 21914 15056
rect 21970 15000 23490 15056
rect 21909 14998 23490 15000
rect 21909 14995 21975 14998
rect 26182 14996 26188 15060
rect 26252 15058 26258 15060
rect 27286 15058 27292 15060
rect 26252 14998 27292 15058
rect 27356 15058 27403 15060
rect 38193 15058 38259 15061
rect 39200 15058 39800 15088
rect 27356 15056 27448 15058
rect 27398 15000 27448 15056
rect 26252 14996 26258 14998
rect 27286 14996 27292 14998
rect 27356 14998 27448 15000
rect 38193 15056 39800 15058
rect 38193 15000 38198 15056
rect 38254 15000 39800 15056
rect 38193 14998 39800 15000
rect 27356 14996 27403 14998
rect 27337 14995 27403 14996
rect 38193 14995 38259 14998
rect 39200 14968 39800 14998
rect 26049 14922 26115 14925
rect 12065 14920 17050 14922
rect 12065 14864 12070 14920
rect 12126 14864 17050 14920
rect 12065 14862 17050 14864
rect 17174 14920 26115 14922
rect 17174 14864 26054 14920
rect 26110 14864 26115 14920
rect 17174 14862 26115 14864
rect 12065 14859 12131 14862
rect 5073 14786 5139 14789
rect 7557 14786 7623 14789
rect 5073 14784 7623 14786
rect 5073 14728 5078 14784
rect 5134 14728 7562 14784
rect 7618 14728 7623 14784
rect 5073 14726 7623 14728
rect 5073 14723 5139 14726
rect 7557 14723 7623 14726
rect 8201 14786 8267 14789
rect 12709 14786 12775 14789
rect 8201 14784 12775 14786
rect 8201 14728 8206 14784
rect 8262 14728 12714 14784
rect 12770 14728 12775 14784
rect 8201 14726 12775 14728
rect 8201 14723 8267 14726
rect 12709 14723 12775 14726
rect 13997 14786 14063 14789
rect 16297 14786 16363 14789
rect 13997 14784 16363 14786
rect 13997 14728 14002 14784
rect 14058 14728 16302 14784
rect 16358 14728 16363 14784
rect 13997 14726 16363 14728
rect 13997 14723 14063 14726
rect 16297 14723 16363 14726
rect 16481 14786 16547 14789
rect 16665 14786 16731 14789
rect 16481 14784 16731 14786
rect 16481 14728 16486 14784
rect 16542 14728 16670 14784
rect 16726 14728 16731 14784
rect 16481 14726 16731 14728
rect 16990 14786 17050 14862
rect 26049 14859 26115 14862
rect 19190 14786 19196 14788
rect 16990 14726 19196 14786
rect 16481 14723 16547 14726
rect 16665 14723 16731 14726
rect 19190 14724 19196 14726
rect 19260 14786 19266 14788
rect 20897 14786 20963 14789
rect 19260 14784 20963 14786
rect 19260 14728 20902 14784
rect 20958 14728 20963 14784
rect 19260 14726 20963 14728
rect 19260 14724 19266 14726
rect 20897 14723 20963 14726
rect 21030 14724 21036 14788
rect 21100 14786 21106 14788
rect 22277 14786 22343 14789
rect 22502 14786 22508 14788
rect 21100 14726 21972 14786
rect 21100 14724 21106 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 11789 14650 11855 14653
rect 15837 14650 15903 14653
rect 11789 14648 15903 14650
rect 11789 14592 11794 14648
rect 11850 14592 15842 14648
rect 15898 14592 15903 14648
rect 11789 14590 15903 14592
rect 11789 14587 11855 14590
rect 15837 14587 15903 14590
rect 16113 14650 16179 14653
rect 18321 14650 18387 14653
rect 16113 14648 18387 14650
rect 16113 14592 16118 14648
rect 16174 14592 18326 14648
rect 18382 14592 18387 14648
rect 16113 14590 18387 14592
rect 16113 14587 16179 14590
rect 18321 14587 18387 14590
rect 18454 14588 18460 14652
rect 18524 14650 18530 14652
rect 21725 14650 21791 14653
rect 18524 14648 21791 14650
rect 18524 14592 21730 14648
rect 21786 14592 21791 14648
rect 18524 14590 21791 14592
rect 21912 14650 21972 14726
rect 22277 14784 22508 14786
rect 22277 14728 22282 14784
rect 22338 14728 22508 14784
rect 22277 14726 22508 14728
rect 22277 14723 22343 14726
rect 22502 14724 22508 14726
rect 22572 14724 22578 14788
rect 25313 14786 25379 14789
rect 27061 14786 27127 14789
rect 25313 14784 27127 14786
rect 25313 14728 25318 14784
rect 25374 14728 27066 14784
rect 27122 14728 27127 14784
rect 25313 14726 27127 14728
rect 25313 14723 25379 14726
rect 27061 14723 27127 14726
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 26601 14650 26667 14653
rect 21912 14648 26667 14650
rect 21912 14592 26606 14648
rect 26662 14592 26667 14648
rect 21912 14590 26667 14592
rect 18524 14588 18530 14590
rect 21725 14587 21791 14590
rect 26601 14587 26667 14590
rect 10777 14514 10843 14517
rect 12433 14514 12499 14517
rect 10777 14512 12499 14514
rect 10777 14456 10782 14512
rect 10838 14456 12438 14512
rect 12494 14456 12499 14512
rect 10777 14454 12499 14456
rect 10777 14451 10843 14454
rect 12433 14451 12499 14454
rect 14641 14514 14707 14517
rect 14774 14514 14780 14516
rect 14641 14512 14780 14514
rect 14641 14456 14646 14512
rect 14702 14456 14780 14512
rect 14641 14454 14780 14456
rect 14641 14451 14707 14454
rect 14774 14452 14780 14454
rect 14844 14452 14850 14516
rect 15878 14452 15884 14516
rect 15948 14514 15954 14516
rect 16205 14514 16271 14517
rect 15948 14512 16271 14514
rect 15948 14456 16210 14512
rect 16266 14456 16271 14512
rect 15948 14454 16271 14456
rect 15948 14452 15954 14454
rect 16205 14451 16271 14454
rect 16481 14514 16547 14517
rect 20897 14514 20963 14517
rect 21081 14516 21147 14517
rect 16481 14512 20963 14514
rect 16481 14456 16486 14512
rect 16542 14456 20902 14512
rect 20958 14456 20963 14512
rect 16481 14454 20963 14456
rect 16481 14451 16547 14454
rect 20897 14451 20963 14454
rect 21030 14452 21036 14516
rect 21100 14514 21147 14516
rect 21541 14514 21607 14517
rect 23289 14514 23355 14517
rect 21100 14512 21192 14514
rect 21142 14456 21192 14512
rect 21100 14454 21192 14456
rect 21541 14512 23355 14514
rect 21541 14456 21546 14512
rect 21602 14456 23294 14512
rect 23350 14456 23355 14512
rect 21541 14454 23355 14456
rect 21100 14452 21147 14454
rect 21081 14451 21147 14452
rect 21541 14451 21607 14454
rect 23289 14451 23355 14454
rect 25865 14514 25931 14517
rect 28809 14514 28875 14517
rect 25865 14512 28875 14514
rect 25865 14456 25870 14512
rect 25926 14456 28814 14512
rect 28870 14456 28875 14512
rect 25865 14454 28875 14456
rect 25865 14451 25931 14454
rect 28809 14451 28875 14454
rect 6821 14378 6887 14381
rect 25957 14378 26023 14381
rect 6821 14376 26023 14378
rect 6821 14320 6826 14376
rect 6882 14320 25962 14376
rect 26018 14320 26023 14376
rect 6821 14318 26023 14320
rect 6821 14315 6887 14318
rect 25957 14315 26023 14318
rect 27153 14378 27219 14381
rect 28165 14378 28231 14381
rect 27153 14376 28231 14378
rect 27153 14320 27158 14376
rect 27214 14320 28170 14376
rect 28226 14320 28231 14376
rect 27153 14318 28231 14320
rect 27153 14315 27219 14318
rect 28165 14315 28231 14318
rect 38193 14378 38259 14381
rect 39200 14378 39800 14408
rect 38193 14376 39800 14378
rect 38193 14320 38198 14376
rect 38254 14320 39800 14376
rect 38193 14318 39800 14320
rect 38193 14315 38259 14318
rect 39200 14288 39800 14318
rect 6821 14242 6887 14245
rect 16389 14242 16455 14245
rect 18505 14242 18571 14245
rect 19333 14244 19399 14245
rect 6821 14240 16314 14242
rect 6821 14184 6826 14240
rect 6882 14184 16314 14240
rect 6821 14182 16314 14184
rect 6821 14179 6887 14182
rect 4521 14106 4587 14109
rect 5625 14106 5691 14109
rect 6126 14106 6132 14108
rect 4521 14104 6132 14106
rect 4521 14048 4526 14104
rect 4582 14048 5630 14104
rect 5686 14048 6132 14104
rect 4521 14046 6132 14048
rect 4521 14043 4587 14046
rect 5625 14043 5691 14046
rect 6126 14044 6132 14046
rect 6196 14044 6202 14108
rect 10593 14106 10659 14109
rect 14958 14106 14964 14108
rect 10593 14104 14964 14106
rect 10593 14048 10598 14104
rect 10654 14048 14964 14104
rect 10593 14046 14964 14048
rect 10593 14043 10659 14046
rect 14958 14044 14964 14046
rect 15028 14044 15034 14108
rect 16254 14106 16314 14182
rect 16389 14240 18571 14242
rect 16389 14184 16394 14240
rect 16450 14184 18510 14240
rect 18566 14184 18571 14240
rect 16389 14182 18571 14184
rect 16389 14179 16455 14182
rect 18505 14179 18571 14182
rect 18822 14180 18828 14244
rect 18892 14242 18898 14244
rect 19190 14242 19196 14244
rect 18892 14182 19196 14242
rect 18892 14180 18898 14182
rect 19190 14180 19196 14182
rect 19260 14180 19266 14244
rect 19333 14240 19380 14244
rect 19444 14242 19450 14244
rect 20345 14242 20411 14245
rect 22001 14242 22067 14245
rect 25037 14242 25103 14245
rect 26417 14244 26483 14245
rect 19333 14184 19338 14240
rect 19333 14180 19380 14184
rect 19444 14182 19490 14242
rect 20345 14240 22067 14242
rect 20345 14184 20350 14240
rect 20406 14184 22006 14240
rect 22062 14184 22067 14240
rect 20345 14182 22067 14184
rect 19444 14180 19450 14182
rect 19333 14179 19399 14180
rect 20345 14179 20411 14182
rect 22001 14179 22067 14182
rect 22142 14240 25103 14242
rect 22142 14184 25042 14240
rect 25098 14184 25103 14240
rect 22142 14182 25103 14184
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 18454 14106 18460 14108
rect 16254 14046 18460 14106
rect 18454 14044 18460 14046
rect 18524 14044 18530 14108
rect 18822 14044 18828 14108
rect 18892 14106 18898 14108
rect 19425 14106 19491 14109
rect 18892 14104 19491 14106
rect 18892 14048 19430 14104
rect 19486 14048 19491 14104
rect 18892 14046 19491 14048
rect 18892 14044 18898 14046
rect 19425 14043 19491 14046
rect 21817 14106 21883 14109
rect 22142 14106 22202 14182
rect 25037 14179 25103 14182
rect 26366 14180 26372 14244
rect 26436 14242 26483 14244
rect 26601 14242 26667 14245
rect 26436 14240 26667 14242
rect 26478 14184 26606 14240
rect 26662 14184 26667 14240
rect 26436 14182 26667 14184
rect 26436 14180 26483 14182
rect 26417 14179 26483 14180
rect 26601 14179 26667 14182
rect 21817 14104 22202 14106
rect 21817 14048 21822 14104
rect 21878 14048 22202 14104
rect 21817 14046 22202 14048
rect 22277 14106 22343 14109
rect 26601 14106 26667 14109
rect 22277 14104 26667 14106
rect 22277 14048 22282 14104
rect 22338 14048 26606 14104
rect 26662 14048 26667 14104
rect 22277 14046 26667 14048
rect 21817 14043 21883 14046
rect 22277 14043 22343 14046
rect 26601 14043 26667 14046
rect 5942 13908 5948 13972
rect 6012 13970 6018 13972
rect 10041 13970 10107 13973
rect 16481 13970 16547 13973
rect 6012 13968 16547 13970
rect 6012 13912 10046 13968
rect 10102 13912 16486 13968
rect 16542 13912 16547 13968
rect 6012 13910 16547 13912
rect 6012 13908 6018 13910
rect 10041 13907 10107 13910
rect 16481 13907 16547 13910
rect 16614 13908 16620 13972
rect 16684 13970 16690 13972
rect 25998 13970 26004 13972
rect 16684 13910 26004 13970
rect 16684 13908 16690 13910
rect 25998 13908 26004 13910
rect 26068 13908 26074 13972
rect 29085 13970 29151 13973
rect 30373 13970 30439 13973
rect 29085 13968 30439 13970
rect 29085 13912 29090 13968
rect 29146 13912 30378 13968
rect 30434 13912 30439 13968
rect 29085 13910 30439 13912
rect 29085 13907 29151 13910
rect 30373 13907 30439 13910
rect 10501 13834 10567 13837
rect 12249 13834 12315 13837
rect 10501 13832 12315 13834
rect 10501 13776 10506 13832
rect 10562 13776 12254 13832
rect 12310 13776 12315 13832
rect 10501 13774 12315 13776
rect 10501 13771 10567 13774
rect 12249 13771 12315 13774
rect 13813 13834 13879 13837
rect 18505 13834 18571 13837
rect 13813 13832 18571 13834
rect 13813 13776 13818 13832
rect 13874 13776 18510 13832
rect 18566 13776 18571 13832
rect 13813 13774 18571 13776
rect 13813 13771 13879 13774
rect 18505 13771 18571 13774
rect 18689 13834 18755 13837
rect 20621 13834 20687 13837
rect 18689 13832 20687 13834
rect 18689 13776 18694 13832
rect 18750 13776 20626 13832
rect 20682 13776 20687 13832
rect 18689 13774 20687 13776
rect 18689 13771 18755 13774
rect 20621 13771 20687 13774
rect 20897 13834 20963 13837
rect 22369 13834 22435 13837
rect 20897 13832 22435 13834
rect 20897 13776 20902 13832
rect 20958 13776 22374 13832
rect 22430 13776 22435 13832
rect 20897 13774 22435 13776
rect 20897 13771 20963 13774
rect 22369 13771 22435 13774
rect 27102 13772 27108 13836
rect 27172 13834 27178 13836
rect 27245 13834 27311 13837
rect 27172 13832 27311 13834
rect 27172 13776 27250 13832
rect 27306 13776 27311 13832
rect 27172 13774 27311 13776
rect 27172 13772 27178 13774
rect 27245 13771 27311 13774
rect 27613 13836 27679 13837
rect 27613 13832 27660 13836
rect 27724 13834 27730 13836
rect 27613 13776 27618 13832
rect 27613 13772 27660 13776
rect 27724 13774 27770 13834
rect 27724 13772 27730 13774
rect 27613 13771 27679 13772
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 9213 13698 9279 13701
rect 16389 13698 16455 13701
rect 20345 13698 20411 13701
rect 21081 13700 21147 13701
rect 9213 13696 16314 13698
rect 9213 13640 9218 13696
rect 9274 13640 16314 13696
rect 9213 13638 16314 13640
rect 9213 13635 9279 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 6729 13562 6795 13565
rect 10358 13562 10364 13564
rect 6729 13560 10364 13562
rect 6729 13504 6734 13560
rect 6790 13504 10364 13560
rect 6729 13502 10364 13504
rect 6729 13499 6795 13502
rect 10358 13500 10364 13502
rect 10428 13562 10434 13564
rect 13261 13562 13327 13565
rect 10428 13560 13327 13562
rect 10428 13504 13266 13560
rect 13322 13504 13327 13560
rect 10428 13502 13327 13504
rect 10428 13500 10434 13502
rect 13261 13499 13327 13502
rect 13629 13562 13695 13565
rect 14774 13562 14780 13564
rect 13629 13560 14780 13562
rect 13629 13504 13634 13560
rect 13690 13504 14780 13560
rect 13629 13502 14780 13504
rect 13629 13499 13695 13502
rect 14774 13500 14780 13502
rect 14844 13500 14850 13564
rect 16254 13562 16314 13638
rect 16389 13696 20411 13698
rect 16389 13640 16394 13696
rect 16450 13640 20350 13696
rect 20406 13640 20411 13696
rect 16389 13638 20411 13640
rect 16389 13635 16455 13638
rect 20345 13635 20411 13638
rect 21030 13636 21036 13700
rect 21100 13698 21147 13700
rect 21100 13696 21192 13698
rect 21142 13640 21192 13696
rect 21100 13638 21192 13640
rect 21100 13636 21147 13638
rect 21398 13636 21404 13700
rect 21468 13698 21474 13700
rect 21817 13698 21883 13701
rect 21468 13696 21883 13698
rect 21468 13640 21822 13696
rect 21878 13640 21883 13696
rect 21468 13638 21883 13640
rect 21468 13636 21474 13638
rect 21081 13635 21147 13636
rect 21817 13635 21883 13638
rect 22093 13698 22159 13701
rect 22645 13698 22711 13701
rect 22093 13696 22711 13698
rect 22093 13640 22098 13696
rect 22154 13640 22650 13696
rect 22706 13640 22711 13696
rect 22093 13638 22711 13640
rect 22093 13635 22159 13638
rect 22645 13635 22711 13638
rect 38285 13698 38351 13701
rect 39200 13698 39800 13728
rect 38285 13696 39800 13698
rect 38285 13640 38290 13696
rect 38346 13640 39800 13696
rect 38285 13638 39800 13640
rect 38285 13635 38351 13638
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 16941 13562 17007 13565
rect 16254 13560 17007 13562
rect 16254 13504 16946 13560
rect 17002 13504 17007 13560
rect 16254 13502 17007 13504
rect 16941 13499 17007 13502
rect 17217 13562 17283 13565
rect 26601 13562 26667 13565
rect 17217 13560 26667 13562
rect 17217 13504 17222 13560
rect 17278 13504 26606 13560
rect 26662 13504 26667 13560
rect 17217 13502 26667 13504
rect 17217 13499 17283 13502
rect 26601 13499 26667 13502
rect 8569 13426 8635 13429
rect 11605 13426 11671 13429
rect 8569 13424 11671 13426
rect 8569 13368 8574 13424
rect 8630 13368 11610 13424
rect 11666 13368 11671 13424
rect 8569 13366 11671 13368
rect 8569 13363 8635 13366
rect 11605 13363 11671 13366
rect 11881 13426 11947 13429
rect 14222 13426 14228 13428
rect 11881 13424 14228 13426
rect 11881 13368 11886 13424
rect 11942 13368 14228 13424
rect 11881 13366 14228 13368
rect 11881 13363 11947 13366
rect 14222 13364 14228 13366
rect 14292 13364 14298 13428
rect 14457 13426 14523 13429
rect 27981 13426 28047 13429
rect 14457 13424 28047 13426
rect 14457 13368 14462 13424
rect 14518 13368 27986 13424
rect 28042 13368 28047 13424
rect 14457 13366 28047 13368
rect 14457 13363 14523 13366
rect 27981 13363 28047 13366
rect 5349 13290 5415 13293
rect 9213 13290 9279 13293
rect 9489 13290 9555 13293
rect 5349 13288 7850 13290
rect 5349 13232 5354 13288
rect 5410 13232 7850 13288
rect 5349 13230 7850 13232
rect 5349 13227 5415 13230
rect 2221 13154 2287 13157
rect 7790 13154 7850 13230
rect 9213 13288 9555 13290
rect 9213 13232 9218 13288
rect 9274 13232 9494 13288
rect 9550 13232 9555 13288
rect 9213 13230 9555 13232
rect 9213 13227 9279 13230
rect 9489 13227 9555 13230
rect 11421 13290 11487 13293
rect 16113 13290 16179 13293
rect 11421 13288 16179 13290
rect 11421 13232 11426 13288
rect 11482 13232 16118 13288
rect 16174 13232 16179 13288
rect 11421 13230 16179 13232
rect 11421 13227 11487 13230
rect 16113 13227 16179 13230
rect 16849 13290 16915 13293
rect 20621 13290 20687 13293
rect 16849 13288 20687 13290
rect 16849 13232 16854 13288
rect 16910 13232 20626 13288
rect 20682 13232 20687 13288
rect 16849 13230 20687 13232
rect 16849 13227 16915 13230
rect 20621 13227 20687 13230
rect 20897 13290 20963 13293
rect 24669 13290 24735 13293
rect 20897 13288 24735 13290
rect 20897 13232 20902 13288
rect 20958 13232 24674 13288
rect 24730 13232 24735 13288
rect 20897 13230 24735 13232
rect 20897 13227 20963 13230
rect 24669 13227 24735 13230
rect 13118 13154 13124 13156
rect 2221 13152 7666 13154
rect 2221 13096 2226 13152
rect 2282 13096 7666 13152
rect 2221 13094 7666 13096
rect 7790 13094 13124 13154
rect 2221 13091 2287 13094
rect 200 13018 800 13048
rect 3785 13018 3851 13021
rect 200 13016 3851 13018
rect 200 12960 3790 13016
rect 3846 12960 3851 13016
rect 200 12958 3851 12960
rect 200 12928 800 12958
rect 3785 12955 3851 12958
rect 4153 13018 4219 13021
rect 6913 13018 6979 13021
rect 4153 13016 6979 13018
rect 4153 12960 4158 13016
rect 4214 12960 6918 13016
rect 6974 12960 6979 13016
rect 4153 12958 6979 12960
rect 7606 13018 7666 13094
rect 13118 13092 13124 13094
rect 13188 13092 13194 13156
rect 15193 13154 15259 13157
rect 15469 13154 15535 13157
rect 18873 13154 18939 13157
rect 19057 13156 19123 13157
rect 15193 13152 18939 13154
rect 15193 13096 15198 13152
rect 15254 13096 15474 13152
rect 15530 13096 18878 13152
rect 18934 13096 18939 13152
rect 15193 13094 18939 13096
rect 15193 13091 15259 13094
rect 15469 13091 15535 13094
rect 18873 13091 18939 13094
rect 19006 13092 19012 13156
rect 19076 13154 19123 13156
rect 21909 13154 21975 13157
rect 23105 13154 23171 13157
rect 19076 13152 19168 13154
rect 19118 13096 19168 13152
rect 19076 13094 19168 13096
rect 21909 13152 23171 13154
rect 21909 13096 21914 13152
rect 21970 13096 23110 13152
rect 23166 13096 23171 13152
rect 21909 13094 23171 13096
rect 19076 13092 19123 13094
rect 19057 13091 19123 13092
rect 21909 13091 21975 13094
rect 23105 13091 23171 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 15694 13018 15700 13020
rect 7606 12958 15700 13018
rect 4153 12955 4219 12958
rect 6913 12955 6979 12958
rect 15694 12956 15700 12958
rect 15764 12956 15770 13020
rect 16665 13018 16731 13021
rect 16665 13016 19258 13018
rect 16665 12960 16670 13016
rect 16726 12960 19258 13016
rect 16665 12958 19258 12960
rect 16665 12955 16731 12958
rect 5441 12884 5507 12885
rect 3918 12820 3924 12884
rect 3988 12882 3994 12884
rect 5390 12882 5396 12884
rect 3988 12822 5274 12882
rect 5350 12822 5396 12882
rect 5460 12880 5507 12884
rect 5502 12824 5507 12880
rect 3988 12820 3994 12822
rect 4521 12746 4587 12749
rect 5022 12746 5028 12748
rect 4521 12744 5028 12746
rect 4521 12688 4526 12744
rect 4582 12688 5028 12744
rect 4521 12686 5028 12688
rect 4521 12683 4587 12686
rect 5022 12684 5028 12686
rect 5092 12684 5098 12748
rect 5214 12746 5274 12822
rect 5390 12820 5396 12822
rect 5460 12820 5507 12824
rect 5441 12819 5507 12820
rect 9489 12882 9555 12885
rect 11053 12882 11119 12885
rect 9489 12880 11119 12882
rect 9489 12824 9494 12880
rect 9550 12824 11058 12880
rect 11114 12824 11119 12880
rect 9489 12822 11119 12824
rect 9489 12819 9555 12822
rect 11053 12819 11119 12822
rect 11605 12882 11671 12885
rect 19006 12882 19012 12884
rect 11605 12880 19012 12882
rect 11605 12824 11610 12880
rect 11666 12824 19012 12880
rect 11605 12822 19012 12824
rect 11605 12819 11671 12822
rect 19006 12820 19012 12822
rect 19076 12820 19082 12884
rect 19198 12882 19258 12958
rect 20110 12956 20116 13020
rect 20180 13018 20186 13020
rect 22737 13018 22803 13021
rect 20180 13016 22803 13018
rect 20180 12960 22742 13016
rect 22798 12960 22803 13016
rect 20180 12958 22803 12960
rect 20180 12956 20186 12958
rect 22737 12955 22803 12958
rect 22921 13018 22987 13021
rect 30373 13018 30439 13021
rect 22921 13016 30439 13018
rect 22921 12960 22926 13016
rect 22982 12960 30378 13016
rect 30434 12960 30439 13016
rect 22921 12958 30439 12960
rect 22921 12955 22987 12958
rect 30373 12955 30439 12958
rect 21030 12882 21036 12884
rect 19198 12822 21036 12882
rect 21030 12820 21036 12822
rect 21100 12820 21106 12884
rect 21725 12882 21791 12885
rect 22369 12882 22435 12885
rect 21725 12880 22435 12882
rect 21725 12824 21730 12880
rect 21786 12824 22374 12880
rect 22430 12824 22435 12880
rect 21725 12822 22435 12824
rect 21725 12819 21791 12822
rect 22369 12819 22435 12822
rect 22553 12882 22619 12885
rect 23013 12882 23079 12885
rect 22553 12880 23079 12882
rect 22553 12824 22558 12880
rect 22614 12824 23018 12880
rect 23074 12824 23079 12880
rect 22553 12822 23079 12824
rect 22553 12819 22619 12822
rect 23013 12819 23079 12822
rect 16665 12746 16731 12749
rect 5214 12744 16731 12746
rect 5214 12688 16670 12744
rect 16726 12688 16731 12744
rect 5214 12686 16731 12688
rect 16665 12683 16731 12686
rect 16798 12684 16804 12748
rect 16868 12746 16874 12748
rect 17585 12746 17651 12749
rect 16868 12744 17651 12746
rect 16868 12688 17590 12744
rect 17646 12688 17651 12744
rect 16868 12686 17651 12688
rect 16868 12684 16874 12686
rect 17585 12683 17651 12686
rect 17953 12746 18019 12749
rect 18086 12746 18092 12748
rect 17953 12744 18092 12746
rect 17953 12688 17958 12744
rect 18014 12688 18092 12744
rect 17953 12686 18092 12688
rect 17953 12683 18019 12686
rect 18086 12684 18092 12686
rect 18156 12684 18162 12748
rect 18321 12746 18387 12749
rect 26509 12746 26575 12749
rect 27337 12746 27403 12749
rect 18321 12744 27403 12746
rect 18321 12688 18326 12744
rect 18382 12688 26514 12744
rect 26570 12688 27342 12744
rect 27398 12688 27403 12744
rect 18321 12686 27403 12688
rect 18321 12683 18387 12686
rect 26509 12683 26575 12686
rect 27337 12683 27403 12686
rect 8109 12610 8175 12613
rect 28901 12610 28967 12613
rect 8109 12608 28967 12610
rect 8109 12552 8114 12608
rect 8170 12552 28906 12608
rect 28962 12552 28967 12608
rect 8109 12550 28967 12552
rect 8109 12547 8175 12550
rect 28901 12547 28967 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 5073 12474 5139 12477
rect 9622 12474 9628 12476
rect 5073 12472 9628 12474
rect 5073 12416 5078 12472
rect 5134 12416 9628 12472
rect 5073 12414 9628 12416
rect 5073 12411 5139 12414
rect 9622 12412 9628 12414
rect 9692 12412 9698 12476
rect 10777 12472 10843 12477
rect 10777 12416 10782 12472
rect 10838 12416 10843 12472
rect 10777 12411 10843 12416
rect 11462 12412 11468 12476
rect 11532 12474 11538 12476
rect 12801 12474 12867 12477
rect 11532 12472 12867 12474
rect 11532 12416 12806 12472
rect 12862 12416 12867 12472
rect 11532 12414 12867 12416
rect 11532 12412 11538 12414
rect 12801 12411 12867 12414
rect 14457 12474 14523 12477
rect 14733 12474 14799 12477
rect 14457 12472 14799 12474
rect 14457 12416 14462 12472
rect 14518 12416 14738 12472
rect 14794 12416 14799 12472
rect 14457 12414 14799 12416
rect 14457 12411 14523 12414
rect 14733 12411 14799 12414
rect 15929 12474 15995 12477
rect 16614 12474 16620 12476
rect 15929 12472 16620 12474
rect 15929 12416 15934 12472
rect 15990 12416 16620 12472
rect 15929 12414 16620 12416
rect 15929 12411 15995 12414
rect 16614 12412 16620 12414
rect 16684 12412 16690 12476
rect 16757 12474 16823 12477
rect 23013 12474 23079 12477
rect 16757 12472 23079 12474
rect 16757 12416 16762 12472
rect 16818 12416 23018 12472
rect 23074 12416 23079 12472
rect 16757 12414 23079 12416
rect 16757 12411 16823 12414
rect 23013 12411 23079 12414
rect 200 12338 800 12368
rect 3877 12338 3943 12341
rect 8569 12340 8635 12341
rect 200 12336 3943 12338
rect 200 12280 3882 12336
rect 3938 12280 3943 12336
rect 200 12278 3943 12280
rect 200 12248 800 12278
rect 3877 12275 3943 12278
rect 8518 12276 8524 12340
rect 8588 12338 8635 12340
rect 10780 12338 10840 12411
rect 11094 12338 11100 12340
rect 8588 12336 8680 12338
rect 8630 12280 8680 12336
rect 8588 12278 8680 12280
rect 10780 12278 11100 12338
rect 8588 12276 8635 12278
rect 11094 12276 11100 12278
rect 11164 12276 11170 12340
rect 12433 12338 12499 12341
rect 13261 12338 13327 12341
rect 20110 12338 20116 12340
rect 12433 12336 20116 12338
rect 12433 12280 12438 12336
rect 12494 12280 13266 12336
rect 13322 12280 20116 12336
rect 12433 12278 20116 12280
rect 8569 12275 8635 12276
rect 12433 12275 12499 12278
rect 13261 12275 13327 12278
rect 20110 12276 20116 12278
rect 20180 12276 20186 12340
rect 20345 12338 20411 12341
rect 20805 12338 20871 12341
rect 20345 12336 20871 12338
rect 20345 12280 20350 12336
rect 20406 12280 20810 12336
rect 20866 12280 20871 12336
rect 20345 12278 20871 12280
rect 20345 12275 20411 12278
rect 20805 12275 20871 12278
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 3693 12202 3759 12205
rect 7005 12202 7071 12205
rect 3693 12200 7071 12202
rect 3693 12144 3698 12200
rect 3754 12144 7010 12200
rect 7066 12144 7071 12200
rect 3693 12142 7071 12144
rect 3693 12139 3759 12142
rect 7005 12139 7071 12142
rect 8385 12202 8451 12205
rect 13813 12202 13879 12205
rect 8385 12200 13879 12202
rect 8385 12144 8390 12200
rect 8446 12144 13818 12200
rect 13874 12144 13879 12200
rect 8385 12142 13879 12144
rect 8385 12139 8451 12142
rect 13813 12139 13879 12142
rect 14549 12202 14615 12205
rect 23933 12202 23999 12205
rect 14549 12200 23999 12202
rect 14549 12144 14554 12200
rect 14610 12144 23938 12200
rect 23994 12144 23999 12200
rect 14549 12142 23999 12144
rect 14549 12139 14615 12142
rect 23933 12139 23999 12142
rect 25129 12202 25195 12205
rect 28257 12202 28323 12205
rect 25129 12200 28323 12202
rect 25129 12144 25134 12200
rect 25190 12144 28262 12200
rect 28318 12144 28323 12200
rect 25129 12142 28323 12144
rect 25129 12139 25195 12142
rect 28257 12139 28323 12142
rect 3969 12066 4035 12069
rect 7373 12066 7439 12069
rect 3969 12064 7439 12066
rect 3969 12008 3974 12064
rect 4030 12008 7378 12064
rect 7434 12008 7439 12064
rect 3969 12006 7439 12008
rect 3969 12003 4035 12006
rect 7373 12003 7439 12006
rect 7925 12066 7991 12069
rect 8569 12066 8635 12069
rect 19149 12066 19215 12069
rect 7925 12064 19215 12066
rect 7925 12008 7930 12064
rect 7986 12008 8574 12064
rect 8630 12008 19154 12064
rect 19210 12008 19215 12064
rect 7925 12006 19215 12008
rect 7925 12003 7991 12006
rect 8569 12003 8635 12006
rect 19149 12003 19215 12006
rect 19977 12066 20043 12069
rect 20621 12068 20687 12069
rect 20621 12066 20668 12068
rect 19977 12064 20668 12066
rect 20732 12066 20738 12068
rect 20897 12066 20963 12069
rect 22318 12066 22324 12068
rect 19977 12008 19982 12064
rect 20038 12008 20626 12064
rect 19977 12006 20668 12008
rect 19977 12003 20043 12006
rect 20621 12004 20668 12006
rect 20732 12006 20814 12066
rect 20897 12064 22324 12066
rect 20897 12008 20902 12064
rect 20958 12008 22324 12064
rect 20897 12006 22324 12008
rect 20732 12004 20738 12006
rect 20621 12003 20687 12004
rect 20897 12003 20963 12006
rect 22318 12004 22324 12006
rect 22388 12004 22394 12068
rect 23197 12066 23263 12069
rect 26049 12066 26115 12069
rect 23197 12064 26115 12066
rect 23197 12008 23202 12064
rect 23258 12008 26054 12064
rect 26110 12008 26115 12064
rect 23197 12006 26115 12008
rect 23197 12003 23263 12006
rect 26049 12003 26115 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 2497 11930 2563 11933
rect 7741 11930 7807 11933
rect 10777 11930 10843 11933
rect 2497 11928 19304 11930
rect 2497 11872 2502 11928
rect 2558 11872 7746 11928
rect 7802 11872 10782 11928
rect 10838 11872 19304 11928
rect 2497 11870 19304 11872
rect 2497 11867 2563 11870
rect 7741 11867 7807 11870
rect 10777 11867 10843 11870
rect 7741 11794 7807 11797
rect 19057 11794 19123 11797
rect 7741 11792 19123 11794
rect 7741 11736 7746 11792
rect 7802 11736 19062 11792
rect 19118 11736 19123 11792
rect 7741 11734 19123 11736
rect 7741 11731 7807 11734
rect 19057 11731 19123 11734
rect 8385 11660 8451 11661
rect 8334 11596 8340 11660
rect 8404 11658 8451 11660
rect 10133 11658 10199 11661
rect 11462 11658 11468 11660
rect 8404 11656 8496 11658
rect 8446 11600 8496 11656
rect 8404 11598 8496 11600
rect 10133 11656 11468 11658
rect 10133 11600 10138 11656
rect 10194 11600 11468 11656
rect 10133 11598 11468 11600
rect 8404 11596 8451 11598
rect 8385 11595 8451 11596
rect 10133 11595 10199 11598
rect 11462 11596 11468 11598
rect 11532 11596 11538 11660
rect 11697 11658 11763 11661
rect 12382 11658 12388 11660
rect 11697 11656 12388 11658
rect 11697 11600 11702 11656
rect 11758 11600 12388 11656
rect 11697 11598 12388 11600
rect 11697 11595 11763 11598
rect 12382 11596 12388 11598
rect 12452 11596 12458 11660
rect 13537 11658 13603 11661
rect 15469 11658 15535 11661
rect 13537 11656 15535 11658
rect 13537 11600 13542 11656
rect 13598 11600 15474 11656
rect 15530 11600 15535 11656
rect 13537 11598 15535 11600
rect 13537 11595 13603 11598
rect 15469 11595 15535 11598
rect 16205 11658 16271 11661
rect 18229 11660 18295 11661
rect 17718 11658 17724 11660
rect 16205 11656 17724 11658
rect 16205 11600 16210 11656
rect 16266 11600 17724 11656
rect 16205 11598 17724 11600
rect 16205 11595 16271 11598
rect 17718 11596 17724 11598
rect 17788 11596 17794 11660
rect 18229 11658 18276 11660
rect 18184 11656 18276 11658
rect 18184 11600 18234 11656
rect 18184 11598 18276 11600
rect 18229 11596 18276 11598
rect 18340 11596 18346 11660
rect 18413 11658 18479 11661
rect 19057 11658 19123 11661
rect 18413 11656 19123 11658
rect 18413 11600 18418 11656
rect 18474 11600 19062 11656
rect 19118 11600 19123 11656
rect 18413 11598 19123 11600
rect 19244 11658 19304 11870
rect 19374 11868 19380 11932
rect 19444 11868 19450 11932
rect 20110 11868 20116 11932
rect 20180 11930 20186 11932
rect 22870 11930 22876 11932
rect 20180 11870 22876 11930
rect 20180 11868 20186 11870
rect 22870 11868 22876 11870
rect 22940 11930 22946 11932
rect 24577 11930 24643 11933
rect 22940 11928 24643 11930
rect 22940 11872 24582 11928
rect 24638 11872 24643 11928
rect 22940 11870 24643 11872
rect 22940 11868 22946 11870
rect 19382 11794 19442 11868
rect 24577 11867 24643 11870
rect 25313 11928 25379 11933
rect 25313 11872 25318 11928
rect 25374 11872 25379 11928
rect 25313 11867 25379 11872
rect 20897 11794 20963 11797
rect 19382 11792 20963 11794
rect 19382 11736 20902 11792
rect 20958 11736 20963 11792
rect 19382 11734 20963 11736
rect 20897 11731 20963 11734
rect 21582 11732 21588 11796
rect 21652 11794 21658 11796
rect 21909 11794 21975 11797
rect 21652 11792 21975 11794
rect 21652 11736 21914 11792
rect 21970 11736 21975 11792
rect 21652 11734 21975 11736
rect 21652 11732 21658 11734
rect 21909 11731 21975 11734
rect 22921 11794 22987 11797
rect 25129 11794 25195 11797
rect 22921 11792 25195 11794
rect 22921 11736 22926 11792
rect 22982 11736 25134 11792
rect 25190 11736 25195 11792
rect 22921 11734 25195 11736
rect 22921 11731 22987 11734
rect 25129 11731 25195 11734
rect 21357 11658 21423 11661
rect 19244 11656 21423 11658
rect 19244 11600 21362 11656
rect 21418 11600 21423 11656
rect 19244 11598 21423 11600
rect 18229 11595 18295 11596
rect 18413 11595 18479 11598
rect 19057 11595 19123 11598
rect 21357 11595 21423 11598
rect 21725 11658 21791 11661
rect 25316 11658 25376 11867
rect 21725 11656 25376 11658
rect 21725 11600 21730 11656
rect 21786 11600 25376 11656
rect 21725 11598 25376 11600
rect 37457 11658 37523 11661
rect 39200 11658 39800 11688
rect 37457 11656 39800 11658
rect 37457 11600 37462 11656
rect 37518 11600 39800 11656
rect 37457 11598 39800 11600
rect 21725 11595 21791 11598
rect 37457 11595 37523 11598
rect 39200 11568 39800 11598
rect 5441 11524 5507 11525
rect 5390 11522 5396 11524
rect 5350 11462 5396 11522
rect 5460 11520 5507 11524
rect 5502 11464 5507 11520
rect 5390 11460 5396 11462
rect 5460 11460 5507 11464
rect 5441 11459 5507 11460
rect 8201 11522 8267 11525
rect 19972 11522 19978 11524
rect 8201 11520 19978 11522
rect 8201 11464 8206 11520
rect 8262 11464 19978 11520
rect 8201 11462 19978 11464
rect 8201 11459 8267 11462
rect 19972 11460 19978 11462
rect 20042 11460 20048 11524
rect 21398 11522 21404 11524
rect 20118 11462 21404 11522
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 11053 11386 11119 11389
rect 12433 11386 12499 11389
rect 11053 11384 12499 11386
rect 11053 11328 11058 11384
rect 11114 11328 12438 11384
rect 12494 11328 12499 11384
rect 11053 11326 12499 11328
rect 11053 11323 11119 11326
rect 12433 11323 12499 11326
rect 13118 11324 13124 11388
rect 13188 11386 13194 11388
rect 13813 11386 13879 11389
rect 13188 11384 13879 11386
rect 13188 11328 13818 11384
rect 13874 11328 13879 11384
rect 13188 11326 13879 11328
rect 13188 11324 13194 11326
rect 13813 11323 13879 11326
rect 14549 11386 14615 11389
rect 17534 11386 17540 11388
rect 14549 11384 17540 11386
rect 14549 11328 14554 11384
rect 14610 11328 17540 11384
rect 14549 11326 17540 11328
rect 14549 11323 14615 11326
rect 17534 11324 17540 11326
rect 17604 11324 17610 11388
rect 17718 11324 17724 11388
rect 17788 11386 17794 11388
rect 20118 11386 20178 11462
rect 21398 11460 21404 11462
rect 21468 11460 21474 11524
rect 22001 11522 22067 11525
rect 22318 11522 22324 11524
rect 22001 11520 22324 11522
rect 22001 11464 22006 11520
rect 22062 11464 22324 11520
rect 22001 11462 22324 11464
rect 22001 11459 22067 11462
rect 22318 11460 22324 11462
rect 22388 11522 22394 11524
rect 24577 11522 24643 11525
rect 22388 11520 24643 11522
rect 22388 11464 24582 11520
rect 24638 11464 24643 11520
rect 22388 11462 24643 11464
rect 22388 11460 22394 11462
rect 24577 11459 24643 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 17788 11326 20178 11386
rect 20253 11386 20319 11389
rect 20478 11386 20484 11388
rect 20253 11384 20484 11386
rect 20253 11328 20258 11384
rect 20314 11328 20484 11384
rect 20253 11326 20484 11328
rect 17788 11324 17794 11326
rect 20253 11323 20319 11326
rect 20478 11324 20484 11326
rect 20548 11324 20554 11388
rect 20713 11386 20779 11389
rect 25589 11386 25655 11389
rect 20713 11384 25655 11386
rect 20713 11328 20718 11384
rect 20774 11328 25594 11384
rect 25650 11328 25655 11384
rect 20713 11326 25655 11328
rect 20713 11323 20779 11326
rect 25589 11323 25655 11326
rect 3417 11250 3483 11253
rect 6729 11250 6795 11253
rect 29269 11250 29335 11253
rect 3417 11248 29335 11250
rect 3417 11192 3422 11248
rect 3478 11192 6734 11248
rect 6790 11192 29274 11248
rect 29330 11192 29335 11248
rect 3417 11190 29335 11192
rect 3417 11187 3483 11190
rect 6729 11187 6795 11190
rect 29269 11187 29335 11190
rect 3877 11114 3943 11117
rect 7925 11114 7991 11117
rect 13537 11114 13603 11117
rect 3877 11112 4170 11114
rect 3877 11056 3882 11112
rect 3938 11056 4170 11112
rect 3877 11054 4170 11056
rect 3877 11051 3943 11054
rect 200 10978 800 11008
rect 3877 10978 3943 10981
rect 200 10976 3943 10978
rect 200 10920 3882 10976
rect 3938 10920 3943 10976
rect 200 10918 3943 10920
rect 200 10888 800 10918
rect 3877 10915 3943 10918
rect 4110 10842 4170 11054
rect 7925 11112 13603 11114
rect 7925 11056 7930 11112
rect 7986 11056 13542 11112
rect 13598 11056 13603 11112
rect 7925 11054 13603 11056
rect 7925 11051 7991 11054
rect 13537 11051 13603 11054
rect 13997 11114 14063 11117
rect 17401 11114 17467 11117
rect 18638 11114 18644 11116
rect 13997 11112 17467 11114
rect 13997 11056 14002 11112
rect 14058 11056 17406 11112
rect 17462 11056 17467 11112
rect 13997 11054 17467 11056
rect 13997 11051 14063 11054
rect 17401 11051 17467 11054
rect 17542 11054 18644 11114
rect 4797 10978 4863 10981
rect 8661 10978 8727 10981
rect 4797 10976 8727 10978
rect 4797 10920 4802 10976
rect 4858 10920 8666 10976
rect 8722 10920 8727 10976
rect 4797 10918 8727 10920
rect 4797 10915 4863 10918
rect 8661 10915 8727 10918
rect 9254 10916 9260 10980
rect 9324 10978 9330 10980
rect 10777 10978 10843 10981
rect 12893 10978 12959 10981
rect 13997 10978 14063 10981
rect 14457 10980 14523 10981
rect 14406 10978 14412 10980
rect 9324 10976 10843 10978
rect 9324 10920 10782 10976
rect 10838 10920 10843 10976
rect 9324 10918 10843 10920
rect 9324 10916 9330 10918
rect 10777 10915 10843 10918
rect 11332 10918 12496 10978
rect 10726 10842 10732 10844
rect 4110 10782 10732 10842
rect 10726 10780 10732 10782
rect 10796 10780 10802 10844
rect 11332 10842 11392 10918
rect 10964 10782 11392 10842
rect 11697 10842 11763 10845
rect 12249 10842 12315 10845
rect 11697 10840 12315 10842
rect 11697 10784 11702 10840
rect 11758 10784 12254 10840
rect 12310 10784 12315 10840
rect 11697 10782 12315 10784
rect 12436 10842 12496 10918
rect 12893 10976 14063 10978
rect 12893 10920 12898 10976
rect 12954 10920 14002 10976
rect 14058 10920 14063 10976
rect 12893 10918 14063 10920
rect 14330 10918 14412 10978
rect 14476 10978 14523 10980
rect 16665 10978 16731 10981
rect 17542 10978 17602 11054
rect 18638 11052 18644 11054
rect 18708 11052 18714 11116
rect 18781 11114 18847 11117
rect 23933 11114 23999 11117
rect 18781 11112 23999 11114
rect 18781 11056 18786 11112
rect 18842 11056 23938 11112
rect 23994 11056 23999 11112
rect 18781 11054 23999 11056
rect 18781 11051 18847 11054
rect 23933 11051 23999 11054
rect 14476 10976 17602 10978
rect 14518 10920 16670 10976
rect 16726 10920 17602 10976
rect 12893 10915 12959 10918
rect 13997 10915 14063 10918
rect 14406 10916 14412 10918
rect 14476 10918 17602 10920
rect 17677 10978 17743 10981
rect 17902 10978 17908 10980
rect 17677 10976 17908 10978
rect 17677 10920 17682 10976
rect 17738 10920 17908 10976
rect 17677 10918 17908 10920
rect 14476 10916 14523 10918
rect 14457 10915 14523 10916
rect 16665 10915 16731 10918
rect 17677 10915 17743 10918
rect 17902 10916 17908 10918
rect 17972 10916 17978 10980
rect 18229 10978 18295 10981
rect 19241 10980 19307 10981
rect 18638 10978 18644 10980
rect 18229 10976 18644 10978
rect 18229 10920 18234 10976
rect 18290 10920 18644 10976
rect 18229 10918 18644 10920
rect 18229 10915 18295 10918
rect 18638 10916 18644 10918
rect 18708 10916 18714 10980
rect 19190 10978 19196 10980
rect 19150 10918 19196 10978
rect 19260 10976 19307 10980
rect 19302 10920 19307 10976
rect 19190 10916 19196 10918
rect 19260 10916 19307 10920
rect 19241 10915 19307 10916
rect 20345 10978 20411 10981
rect 26785 10978 26851 10981
rect 20345 10976 26851 10978
rect 20345 10920 20350 10976
rect 20406 10920 26790 10976
rect 26846 10920 26851 10976
rect 20345 10918 26851 10920
rect 20345 10915 20411 10918
rect 26785 10915 26851 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 12934 10842 12940 10844
rect 12436 10782 12940 10842
rect 6637 10706 6703 10709
rect 8293 10706 8359 10709
rect 6637 10704 8359 10706
rect 6637 10648 6642 10704
rect 6698 10648 8298 10704
rect 8354 10648 8359 10704
rect 6637 10646 8359 10648
rect 6637 10643 6703 10646
rect 8293 10643 8359 10646
rect 10501 10706 10567 10709
rect 10964 10706 11024 10782
rect 11697 10779 11763 10782
rect 12249 10779 12315 10782
rect 12934 10780 12940 10782
rect 13004 10780 13010 10844
rect 13486 10780 13492 10844
rect 13556 10842 13562 10844
rect 13721 10842 13787 10845
rect 19374 10842 19380 10844
rect 13556 10840 19380 10842
rect 13556 10784 13726 10840
rect 13782 10784 19380 10840
rect 13556 10782 19380 10784
rect 13556 10780 13562 10782
rect 13721 10779 13787 10782
rect 19374 10780 19380 10782
rect 19444 10780 19450 10844
rect 20110 10780 20116 10844
rect 20180 10842 20186 10844
rect 26141 10842 26207 10845
rect 20180 10840 26207 10842
rect 20180 10784 26146 10840
rect 26202 10784 26207 10840
rect 20180 10782 26207 10784
rect 20180 10780 20186 10782
rect 26141 10779 26207 10782
rect 10501 10704 11024 10706
rect 10501 10648 10506 10704
rect 10562 10648 11024 10704
rect 10501 10646 11024 10648
rect 11145 10706 11211 10709
rect 14222 10706 14228 10708
rect 11145 10704 14228 10706
rect 11145 10648 11150 10704
rect 11206 10648 14228 10704
rect 11145 10646 14228 10648
rect 10501 10643 10567 10646
rect 11145 10643 11211 10646
rect 14222 10644 14228 10646
rect 14292 10644 14298 10708
rect 14457 10706 14523 10709
rect 23657 10706 23723 10709
rect 14457 10704 23723 10706
rect 14457 10648 14462 10704
rect 14518 10648 23662 10704
rect 23718 10648 23723 10704
rect 14457 10646 23723 10648
rect 14457 10643 14523 10646
rect 23657 10643 23723 10646
rect 9673 10570 9739 10573
rect 10777 10570 10843 10573
rect 9673 10568 10843 10570
rect 9673 10512 9678 10568
rect 9734 10512 10782 10568
rect 10838 10512 10843 10568
rect 9673 10510 10843 10512
rect 9673 10507 9739 10510
rect 10777 10507 10843 10510
rect 11145 10570 11211 10573
rect 11513 10570 11579 10573
rect 11145 10568 11579 10570
rect 11145 10512 11150 10568
rect 11206 10512 11518 10568
rect 11574 10512 11579 10568
rect 11145 10510 11579 10512
rect 11145 10507 11211 10510
rect 11513 10507 11579 10510
rect 11881 10570 11947 10573
rect 14181 10570 14247 10573
rect 11881 10568 14247 10570
rect 11881 10512 11886 10568
rect 11942 10512 14186 10568
rect 14242 10512 14247 10568
rect 11881 10510 14247 10512
rect 11881 10507 11947 10510
rect 14181 10507 14247 10510
rect 14825 10570 14891 10573
rect 17718 10570 17724 10572
rect 14825 10568 17724 10570
rect 14825 10512 14830 10568
rect 14886 10512 17724 10568
rect 14825 10510 17724 10512
rect 14825 10507 14891 10510
rect 17718 10508 17724 10510
rect 17788 10508 17794 10572
rect 17902 10508 17908 10572
rect 17972 10570 17978 10572
rect 26877 10570 26943 10573
rect 17972 10568 26943 10570
rect 17972 10512 26882 10568
rect 26938 10512 26943 10568
rect 17972 10510 26943 10512
rect 17972 10508 17978 10510
rect 26877 10507 26943 10510
rect 5901 10434 5967 10437
rect 11329 10434 11395 10437
rect 14457 10434 14523 10437
rect 5901 10432 6010 10434
rect 5901 10376 5906 10432
rect 5962 10376 6010 10432
rect 5901 10371 6010 10376
rect 11329 10432 14523 10434
rect 11329 10376 11334 10432
rect 11390 10376 14462 10432
rect 14518 10376 14523 10432
rect 11329 10374 14523 10376
rect 11329 10371 11395 10374
rect 14457 10371 14523 10374
rect 14958 10372 14964 10436
rect 15028 10434 15034 10436
rect 15745 10434 15811 10437
rect 15028 10432 15811 10434
rect 15028 10376 15750 10432
rect 15806 10376 15811 10432
rect 15028 10374 15811 10376
rect 15028 10372 15034 10374
rect 15745 10371 15811 10374
rect 16430 10372 16436 10436
rect 16500 10434 16506 10436
rect 20621 10434 20687 10437
rect 16500 10432 20687 10434
rect 16500 10376 20626 10432
rect 20682 10376 20687 10432
rect 16500 10374 20687 10376
rect 16500 10372 16506 10374
rect 20621 10371 20687 10374
rect 20989 10434 21055 10437
rect 22277 10434 22343 10437
rect 20989 10432 22343 10434
rect 20989 10376 20994 10432
rect 21050 10376 22282 10432
rect 22338 10376 22343 10432
rect 20989 10374 22343 10376
rect 20989 10371 21055 10374
rect 22277 10371 22343 10374
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 2865 10298 2931 10301
rect 200 10296 2931 10298
rect 200 10240 2870 10296
rect 2926 10240 2931 10296
rect 200 10238 2931 10240
rect 200 10208 800 10238
rect 2865 10235 2931 10238
rect 5950 10165 6010 10371
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 11094 10236 11100 10300
rect 11164 10298 11170 10300
rect 11329 10298 11395 10301
rect 11164 10296 11395 10298
rect 11164 10240 11334 10296
rect 11390 10240 11395 10296
rect 11164 10238 11395 10240
rect 11164 10236 11170 10238
rect 11329 10235 11395 10238
rect 11513 10298 11579 10301
rect 14181 10298 14247 10301
rect 11513 10296 14247 10298
rect 11513 10240 11518 10296
rect 11574 10240 14186 10296
rect 14242 10240 14247 10296
rect 11513 10238 14247 10240
rect 11513 10235 11579 10238
rect 14181 10235 14247 10238
rect 15101 10298 15167 10301
rect 20805 10298 20871 10301
rect 23749 10298 23815 10301
rect 15101 10296 23815 10298
rect 15101 10240 15106 10296
rect 15162 10240 20810 10296
rect 20866 10240 23754 10296
rect 23810 10240 23815 10296
rect 15101 10238 23815 10240
rect 15101 10235 15167 10238
rect 20805 10235 20871 10238
rect 23749 10235 23815 10238
rect 38101 10298 38167 10301
rect 39200 10298 39800 10328
rect 38101 10296 39800 10298
rect 38101 10240 38106 10296
rect 38162 10240 39800 10296
rect 38101 10238 39800 10240
rect 38101 10235 38167 10238
rect 39200 10208 39800 10238
rect 3233 10162 3299 10165
rect 3366 10162 3372 10164
rect 3233 10160 3372 10162
rect 3233 10104 3238 10160
rect 3294 10104 3372 10160
rect 3233 10102 3372 10104
rect 3233 10099 3299 10102
rect 3366 10100 3372 10102
rect 3436 10100 3442 10164
rect 5901 10160 6010 10165
rect 5901 10104 5906 10160
rect 5962 10104 6010 10160
rect 5901 10102 6010 10104
rect 8937 10162 9003 10165
rect 12525 10162 12591 10165
rect 8937 10160 12591 10162
rect 8937 10104 8942 10160
rect 8998 10104 12530 10160
rect 12586 10104 12591 10160
rect 8937 10102 12591 10104
rect 5901 10099 5967 10102
rect 8937 10099 9003 10102
rect 12525 10099 12591 10102
rect 12801 10162 12867 10165
rect 13445 10162 13511 10165
rect 12801 10160 13511 10162
rect 12801 10104 12806 10160
rect 12862 10104 13450 10160
rect 13506 10104 13511 10160
rect 12801 10102 13511 10104
rect 12801 10099 12867 10102
rect 13445 10099 13511 10102
rect 13854 10100 13860 10164
rect 13924 10162 13930 10164
rect 16205 10162 16271 10165
rect 13924 10160 16271 10162
rect 13924 10104 16210 10160
rect 16266 10104 16271 10160
rect 13924 10102 16271 10104
rect 13924 10100 13930 10102
rect 16205 10099 16271 10102
rect 16757 10162 16823 10165
rect 17534 10162 17540 10164
rect 16757 10160 17540 10162
rect 16757 10104 16762 10160
rect 16818 10104 17540 10160
rect 16757 10102 17540 10104
rect 16757 10099 16823 10102
rect 17534 10100 17540 10102
rect 17604 10100 17610 10164
rect 18045 10162 18111 10165
rect 20110 10162 20116 10164
rect 18045 10160 20116 10162
rect 18045 10104 18050 10160
rect 18106 10104 20116 10160
rect 18045 10102 20116 10104
rect 18045 10099 18111 10102
rect 20110 10100 20116 10102
rect 20180 10100 20186 10164
rect 20846 10100 20852 10164
rect 20916 10162 20922 10164
rect 21081 10162 21147 10165
rect 25681 10162 25747 10165
rect 20916 10160 25747 10162
rect 20916 10104 21086 10160
rect 21142 10104 25686 10160
rect 25742 10104 25747 10160
rect 20916 10102 25747 10104
rect 20916 10100 20922 10102
rect 21081 10099 21147 10102
rect 25681 10099 25747 10102
rect 7373 10026 7439 10029
rect 12801 10026 12867 10029
rect 7373 10024 12867 10026
rect 7373 9968 7378 10024
rect 7434 9968 12806 10024
rect 12862 9968 12867 10024
rect 7373 9966 12867 9968
rect 7373 9963 7439 9966
rect 12801 9963 12867 9966
rect 12934 9964 12940 10028
rect 13004 10026 13010 10028
rect 13813 10026 13879 10029
rect 13004 10024 13879 10026
rect 13004 9968 13818 10024
rect 13874 9968 13879 10024
rect 13004 9966 13879 9968
rect 13004 9964 13010 9966
rect 13813 9963 13879 9966
rect 16297 10026 16363 10029
rect 16614 10026 16620 10028
rect 16297 10024 16620 10026
rect 16297 9968 16302 10024
rect 16358 9968 16620 10024
rect 16297 9966 16620 9968
rect 16297 9963 16363 9966
rect 16614 9964 16620 9966
rect 16684 9964 16690 10028
rect 16757 10026 16823 10029
rect 24577 10026 24643 10029
rect 16757 10024 24643 10026
rect 16757 9968 16762 10024
rect 16818 9968 24582 10024
rect 24638 9968 24643 10024
rect 16757 9966 24643 9968
rect 16757 9963 16823 9966
rect 24577 9963 24643 9966
rect 4429 9890 4495 9893
rect 8569 9890 8635 9893
rect 4429 9888 8635 9890
rect 4429 9832 4434 9888
rect 4490 9832 8574 9888
rect 8630 9832 8635 9888
rect 4429 9830 8635 9832
rect 4429 9827 4495 9830
rect 8569 9827 8635 9830
rect 10910 9828 10916 9892
rect 10980 9890 10986 9892
rect 11053 9890 11119 9893
rect 10980 9888 11119 9890
rect 10980 9832 11058 9888
rect 11114 9832 11119 9888
rect 10980 9830 11119 9832
rect 10980 9828 10986 9830
rect 11053 9827 11119 9830
rect 11462 9828 11468 9892
rect 11532 9890 11538 9892
rect 13997 9890 14063 9893
rect 11532 9888 14063 9890
rect 11532 9832 14002 9888
rect 14058 9832 14063 9888
rect 11532 9830 14063 9832
rect 11532 9828 11538 9830
rect 13997 9827 14063 9830
rect 15837 9890 15903 9893
rect 18873 9890 18939 9893
rect 19333 9890 19399 9893
rect 15837 9888 19399 9890
rect 15837 9832 15842 9888
rect 15898 9832 18878 9888
rect 18934 9832 19338 9888
rect 19394 9832 19399 9888
rect 15837 9830 19399 9832
rect 15837 9827 15903 9830
rect 18873 9827 18939 9830
rect 19333 9827 19399 9830
rect 20437 9890 20503 9893
rect 20621 9890 20687 9893
rect 20437 9888 20687 9890
rect 20437 9832 20442 9888
rect 20498 9832 20626 9888
rect 20682 9832 20687 9888
rect 20437 9830 20687 9832
rect 20437 9827 20503 9830
rect 20621 9827 20687 9830
rect 21081 9890 21147 9893
rect 21909 9890 21975 9893
rect 27337 9890 27403 9893
rect 21081 9888 21975 9890
rect 21081 9832 21086 9888
rect 21142 9832 21914 9888
rect 21970 9832 21975 9888
rect 21081 9830 21975 9832
rect 21081 9827 21147 9830
rect 21909 9827 21975 9830
rect 26190 9888 27403 9890
rect 26190 9832 27342 9888
rect 27398 9832 27403 9888
rect 26190 9830 27403 9832
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 5625 9754 5691 9757
rect 8753 9754 8819 9757
rect 5625 9752 8819 9754
rect 5625 9696 5630 9752
rect 5686 9696 8758 9752
rect 8814 9696 8819 9752
rect 5625 9694 8819 9696
rect 5625 9691 5691 9694
rect 8753 9691 8819 9694
rect 8937 9754 9003 9757
rect 14406 9754 14412 9756
rect 8937 9752 14412 9754
rect 8937 9696 8942 9752
rect 8998 9696 14412 9752
rect 8937 9694 14412 9696
rect 8937 9691 9003 9694
rect 14406 9692 14412 9694
rect 14476 9692 14482 9756
rect 15510 9692 15516 9756
rect 15580 9754 15586 9756
rect 15653 9754 15719 9757
rect 15580 9752 15719 9754
rect 15580 9696 15658 9752
rect 15714 9696 15719 9752
rect 15580 9694 15719 9696
rect 15580 9692 15586 9694
rect 15653 9691 15719 9694
rect 16021 9754 16087 9757
rect 16757 9754 16823 9757
rect 16021 9752 16823 9754
rect 16021 9696 16026 9752
rect 16082 9696 16762 9752
rect 16818 9696 16823 9752
rect 16021 9694 16823 9696
rect 16021 9691 16087 9694
rect 16757 9691 16823 9694
rect 17217 9754 17283 9757
rect 17217 9752 18108 9754
rect 17217 9696 17222 9752
rect 17278 9696 18108 9752
rect 17217 9694 18108 9696
rect 17217 9691 17283 9694
rect 1158 9556 1164 9620
rect 1228 9618 1234 9620
rect 1393 9618 1459 9621
rect 1228 9616 1459 9618
rect 1228 9560 1398 9616
rect 1454 9560 1459 9616
rect 1228 9558 1459 9560
rect 1228 9556 1234 9558
rect 1393 9555 1459 9558
rect 3969 9618 4035 9621
rect 17677 9618 17743 9621
rect 3969 9616 17743 9618
rect 3969 9560 3974 9616
rect 4030 9560 17682 9616
rect 17738 9560 17743 9616
rect 3969 9558 17743 9560
rect 18048 9618 18108 9694
rect 18638 9692 18644 9756
rect 18708 9754 18714 9756
rect 19374 9754 19380 9756
rect 18708 9694 19380 9754
rect 18708 9692 18714 9694
rect 19374 9692 19380 9694
rect 19444 9692 19450 9756
rect 22134 9754 22140 9756
rect 19980 9694 22140 9754
rect 19980 9618 20040 9694
rect 22134 9692 22140 9694
rect 22204 9754 22210 9756
rect 26190 9754 26250 9830
rect 27337 9827 27403 9830
rect 22204 9694 26250 9754
rect 22204 9692 22210 9694
rect 18048 9558 20040 9618
rect 20161 9618 20227 9621
rect 21541 9618 21607 9621
rect 20161 9616 21607 9618
rect 20161 9560 20166 9616
rect 20222 9560 21546 9616
rect 21602 9560 21607 9616
rect 20161 9558 21607 9560
rect 3969 9555 4035 9558
rect 17677 9555 17743 9558
rect 20161 9555 20227 9558
rect 21541 9555 21607 9558
rect 37181 9618 37247 9621
rect 39200 9618 39800 9648
rect 37181 9616 39800 9618
rect 37181 9560 37186 9616
rect 37242 9560 39800 9616
rect 37181 9558 39800 9560
rect 37181 9555 37247 9558
rect 39200 9528 39800 9558
rect 6269 9482 6335 9485
rect 8477 9482 8543 9485
rect 6269 9480 8543 9482
rect 6269 9424 6274 9480
rect 6330 9424 8482 9480
rect 8538 9424 8543 9480
rect 6269 9422 8543 9424
rect 6269 9419 6335 9422
rect 8477 9419 8543 9422
rect 9070 9420 9076 9484
rect 9140 9482 9146 9484
rect 9305 9482 9371 9485
rect 9140 9480 9371 9482
rect 9140 9424 9310 9480
rect 9366 9424 9371 9480
rect 9140 9422 9371 9424
rect 9140 9420 9146 9422
rect 9305 9419 9371 9422
rect 10041 9482 10107 9485
rect 20478 9482 20484 9484
rect 10041 9480 20484 9482
rect 10041 9424 10046 9480
rect 10102 9424 20484 9480
rect 10041 9422 20484 9424
rect 10041 9419 10107 9422
rect 20478 9420 20484 9422
rect 20548 9420 20554 9484
rect 20897 9482 20963 9485
rect 22645 9482 22711 9485
rect 20897 9480 22711 9482
rect 20897 9424 20902 9480
rect 20958 9424 22650 9480
rect 22706 9424 22711 9480
rect 20897 9422 22711 9424
rect 20897 9419 20963 9422
rect 22645 9419 22711 9422
rect 6821 9346 6887 9349
rect 16062 9346 16068 9348
rect 6821 9344 16068 9346
rect 6821 9288 6826 9344
rect 6882 9288 16068 9344
rect 6821 9286 16068 9288
rect 6821 9283 6887 9286
rect 16062 9284 16068 9286
rect 16132 9284 16138 9348
rect 16205 9346 16271 9349
rect 20989 9346 21055 9349
rect 16205 9344 21055 9346
rect 16205 9288 16210 9344
rect 16266 9288 20994 9344
rect 21050 9288 21055 9344
rect 16205 9286 21055 9288
rect 16205 9283 16271 9286
rect 20989 9283 21055 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 7557 9210 7623 9213
rect 20713 9210 20779 9213
rect 7557 9208 20779 9210
rect 7557 9152 7562 9208
rect 7618 9152 20718 9208
rect 20774 9152 20779 9208
rect 7557 9150 20779 9152
rect 7557 9147 7623 9150
rect 20713 9147 20779 9150
rect 21173 9210 21239 9213
rect 24669 9210 24735 9213
rect 21173 9208 24735 9210
rect 21173 9152 21178 9208
rect 21234 9152 24674 9208
rect 24730 9152 24735 9208
rect 21173 9150 24735 9152
rect 21173 9147 21239 9150
rect 24669 9147 24735 9150
rect 6821 9074 6887 9077
rect 10869 9074 10935 9077
rect 6821 9072 10935 9074
rect 6821 9016 6826 9072
rect 6882 9016 10874 9072
rect 10930 9016 10935 9072
rect 6821 9014 10935 9016
rect 6821 9011 6887 9014
rect 10869 9011 10935 9014
rect 11237 9074 11303 9077
rect 11697 9074 11763 9077
rect 11237 9072 11763 9074
rect 11237 9016 11242 9072
rect 11298 9016 11702 9072
rect 11758 9016 11763 9072
rect 11237 9014 11763 9016
rect 11237 9011 11303 9014
rect 11697 9011 11763 9014
rect 11881 9074 11947 9077
rect 12014 9074 12020 9076
rect 11881 9072 12020 9074
rect 11881 9016 11886 9072
rect 11942 9016 12020 9072
rect 11881 9014 12020 9016
rect 11881 9011 11947 9014
rect 12014 9012 12020 9014
rect 12084 9012 12090 9076
rect 12198 9012 12204 9076
rect 12268 9074 12274 9076
rect 13721 9074 13787 9077
rect 12268 9072 13787 9074
rect 12268 9016 13726 9072
rect 13782 9016 13787 9072
rect 12268 9014 13787 9016
rect 12268 9012 12274 9014
rect 13721 9011 13787 9014
rect 14365 9074 14431 9077
rect 16481 9074 16547 9077
rect 14365 9072 16547 9074
rect 14365 9016 14370 9072
rect 14426 9016 16486 9072
rect 16542 9016 16547 9072
rect 14365 9014 16547 9016
rect 14365 9011 14431 9014
rect 16481 9011 16547 9014
rect 16941 9074 17007 9077
rect 17534 9074 17540 9076
rect 16941 9072 17540 9074
rect 16941 9016 16946 9072
rect 17002 9016 17540 9072
rect 16941 9014 17540 9016
rect 16941 9011 17007 9014
rect 17534 9012 17540 9014
rect 17604 9012 17610 9076
rect 18086 9012 18092 9076
rect 18156 9074 18162 9076
rect 18229 9074 18295 9077
rect 18156 9072 18295 9074
rect 18156 9016 18234 9072
rect 18290 9016 18295 9072
rect 18156 9014 18295 9016
rect 18156 9012 18162 9014
rect 18229 9011 18295 9014
rect 19701 9074 19767 9077
rect 21541 9074 21607 9077
rect 24894 9074 24900 9076
rect 19701 9072 21466 9074
rect 19701 9016 19706 9072
rect 19762 9016 21466 9072
rect 19701 9014 21466 9016
rect 19701 9011 19767 9014
rect 200 8938 800 8968
rect 4337 8938 4403 8941
rect 5441 8938 5507 8941
rect 21081 8938 21147 8941
rect 200 8878 2790 8938
rect 200 8848 800 8878
rect 2730 8530 2790 8878
rect 4337 8936 21147 8938
rect 4337 8880 4342 8936
rect 4398 8880 5446 8936
rect 5502 8880 21086 8936
rect 21142 8880 21147 8936
rect 4337 8878 21147 8880
rect 21406 8938 21466 9014
rect 21541 9072 24900 9074
rect 21541 9016 21546 9072
rect 21602 9016 24900 9072
rect 21541 9014 24900 9016
rect 21541 9011 21607 9014
rect 24894 9012 24900 9014
rect 24964 9074 24970 9076
rect 25037 9074 25103 9077
rect 24964 9072 25103 9074
rect 24964 9016 25042 9072
rect 25098 9016 25103 9072
rect 24964 9014 25103 9016
rect 24964 9012 24970 9014
rect 25037 9011 25103 9014
rect 22001 8938 22067 8941
rect 21406 8936 22067 8938
rect 21406 8880 22006 8936
rect 22062 8880 22067 8936
rect 21406 8878 22067 8880
rect 4337 8875 4403 8878
rect 5441 8875 5507 8878
rect 21081 8875 21147 8878
rect 22001 8875 22067 8878
rect 22185 8938 22251 8941
rect 22461 8938 22527 8941
rect 22185 8936 22527 8938
rect 22185 8880 22190 8936
rect 22246 8880 22466 8936
rect 22522 8880 22527 8936
rect 22185 8878 22527 8880
rect 22185 8875 22251 8878
rect 22461 8875 22527 8878
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 2957 8802 3023 8805
rect 16430 8802 16436 8804
rect 2957 8800 16436 8802
rect 2957 8744 2962 8800
rect 3018 8744 16436 8800
rect 2957 8742 16436 8744
rect 2957 8739 3023 8742
rect 16430 8740 16436 8742
rect 16500 8740 16506 8804
rect 16941 8802 17007 8805
rect 16622 8800 17007 8802
rect 16622 8744 16946 8800
rect 17002 8744 17007 8800
rect 16622 8742 17007 8744
rect 7189 8666 7255 8669
rect 7833 8666 7899 8669
rect 7189 8664 7899 8666
rect 7189 8608 7194 8664
rect 7250 8608 7838 8664
rect 7894 8608 7899 8664
rect 7189 8606 7899 8608
rect 7189 8603 7255 8606
rect 7833 8603 7899 8606
rect 8753 8666 8819 8669
rect 10593 8666 10659 8669
rect 8753 8664 10659 8666
rect 8753 8608 8758 8664
rect 8814 8608 10598 8664
rect 10654 8608 10659 8664
rect 8753 8606 10659 8608
rect 8753 8603 8819 8606
rect 10593 8603 10659 8606
rect 10869 8666 10935 8669
rect 11462 8666 11468 8668
rect 10869 8664 11468 8666
rect 10869 8608 10874 8664
rect 10930 8608 11468 8664
rect 10869 8606 11468 8608
rect 10869 8603 10935 8606
rect 11462 8604 11468 8606
rect 11532 8604 11538 8668
rect 11881 8666 11947 8669
rect 16205 8666 16271 8669
rect 11881 8664 16271 8666
rect 11881 8608 11886 8664
rect 11942 8608 16210 8664
rect 16266 8608 16271 8664
rect 11881 8606 16271 8608
rect 11881 8603 11947 8606
rect 16205 8603 16271 8606
rect 16481 8666 16547 8669
rect 16622 8666 16682 8742
rect 16941 8739 17007 8742
rect 17125 8802 17191 8805
rect 17401 8802 17467 8805
rect 17125 8800 17467 8802
rect 17125 8744 17130 8800
rect 17186 8744 17406 8800
rect 17462 8744 17467 8800
rect 17125 8742 17467 8744
rect 17125 8739 17191 8742
rect 17401 8739 17467 8742
rect 18597 8802 18663 8805
rect 19190 8802 19196 8804
rect 18597 8800 19196 8802
rect 18597 8744 18602 8800
rect 18658 8744 19196 8800
rect 18597 8742 19196 8744
rect 18597 8739 18663 8742
rect 19190 8740 19196 8742
rect 19260 8740 19266 8804
rect 20478 8740 20484 8804
rect 20548 8802 20554 8804
rect 20897 8802 20963 8805
rect 20548 8800 20963 8802
rect 20548 8744 20902 8800
rect 20958 8744 20963 8800
rect 20548 8742 20963 8744
rect 20548 8740 20554 8742
rect 20897 8739 20963 8742
rect 21909 8802 21975 8805
rect 26141 8802 26207 8805
rect 21909 8800 26207 8802
rect 21909 8744 21914 8800
rect 21970 8744 26146 8800
rect 26202 8744 26207 8800
rect 21909 8742 26207 8744
rect 21909 8739 21975 8742
rect 26141 8739 26207 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 16481 8664 16682 8666
rect 16481 8608 16486 8664
rect 16542 8608 16682 8664
rect 16481 8606 16682 8608
rect 16757 8666 16823 8669
rect 17350 8666 17356 8668
rect 16757 8664 17356 8666
rect 16757 8608 16762 8664
rect 16818 8608 17356 8664
rect 16757 8606 17356 8608
rect 16481 8603 16547 8606
rect 16757 8603 16823 8606
rect 17350 8604 17356 8606
rect 17420 8666 17426 8668
rect 23381 8666 23447 8669
rect 17420 8606 19488 8666
rect 17420 8604 17426 8606
rect 19428 8564 19488 8606
rect 19980 8664 23447 8666
rect 19980 8608 23386 8664
rect 23442 8608 23447 8664
rect 19980 8606 23447 8608
rect 19980 8564 20040 8606
rect 23381 8603 23447 8606
rect 23565 8666 23631 8669
rect 24577 8666 24643 8669
rect 23565 8664 24643 8666
rect 23565 8608 23570 8664
rect 23626 8608 24582 8664
rect 24638 8608 24643 8664
rect 23565 8606 24643 8608
rect 23565 8603 23631 8606
rect 24577 8603 24643 8606
rect 2730 8470 19304 8530
rect 19428 8504 20040 8564
rect 25497 8530 25563 8533
rect 20118 8528 25563 8530
rect 19244 8428 19304 8470
rect 20118 8472 25502 8528
rect 25558 8472 25563 8528
rect 20118 8470 25563 8472
rect 20118 8428 20178 8470
rect 25497 8467 25563 8470
rect 3969 8394 4035 8397
rect 9438 8394 9444 8396
rect 3969 8392 9444 8394
rect 3969 8336 3974 8392
rect 4030 8336 9444 8392
rect 3969 8334 9444 8336
rect 3969 8331 4035 8334
rect 9438 8332 9444 8334
rect 9508 8332 9514 8396
rect 11329 8394 11395 8397
rect 14038 8394 14044 8396
rect 11329 8392 14044 8394
rect 11329 8336 11334 8392
rect 11390 8336 14044 8392
rect 11329 8334 14044 8336
rect 11329 8331 11395 8334
rect 14038 8332 14044 8334
rect 14108 8394 14114 8396
rect 14181 8394 14247 8397
rect 14108 8392 14247 8394
rect 14108 8336 14186 8392
rect 14242 8336 14247 8392
rect 14108 8334 14247 8336
rect 14108 8332 14114 8334
rect 14181 8331 14247 8334
rect 14590 8332 14596 8396
rect 14660 8394 14666 8396
rect 15193 8394 15259 8397
rect 14660 8392 15259 8394
rect 14660 8336 15198 8392
rect 15254 8336 15259 8392
rect 14660 8334 15259 8336
rect 14660 8332 14666 8334
rect 15193 8331 15259 8334
rect 15878 8332 15884 8396
rect 15948 8394 15954 8396
rect 16389 8394 16455 8397
rect 16849 8394 16915 8397
rect 15948 8392 16915 8394
rect 15948 8336 16394 8392
rect 16450 8336 16854 8392
rect 16910 8336 16915 8392
rect 15948 8334 16915 8336
rect 15948 8332 15954 8334
rect 16389 8331 16455 8334
rect 16849 8331 16915 8334
rect 17953 8394 18019 8397
rect 18597 8394 18663 8397
rect 17953 8392 18663 8394
rect 17953 8336 17958 8392
rect 18014 8336 18602 8392
rect 18658 8336 18663 8392
rect 17953 8334 18663 8336
rect 17953 8331 18019 8334
rect 18597 8331 18663 8334
rect 18873 8394 18939 8397
rect 19057 8394 19123 8397
rect 18873 8392 19123 8394
rect 18873 8336 18878 8392
rect 18934 8336 19062 8392
rect 19118 8336 19123 8392
rect 19244 8368 20178 8428
rect 21817 8394 21883 8397
rect 20256 8392 21883 8394
rect 18873 8334 19123 8336
rect 18873 8331 18939 8334
rect 19057 8331 19123 8334
rect 20256 8336 21822 8392
rect 21878 8336 21883 8392
rect 20256 8334 21883 8336
rect 200 8258 800 8288
rect 3877 8258 3943 8261
rect 200 8256 3943 8258
rect 200 8200 3882 8256
rect 3938 8200 3943 8256
rect 200 8198 3943 8200
rect 200 8168 800 8198
rect 3877 8195 3943 8198
rect 5993 8258 6059 8261
rect 13261 8258 13327 8261
rect 5993 8256 13327 8258
rect 5993 8200 5998 8256
rect 6054 8200 13266 8256
rect 13322 8200 13327 8256
rect 5993 8198 13327 8200
rect 5993 8195 6059 8198
rect 13261 8195 13327 8198
rect 13629 8260 13695 8261
rect 13629 8256 13676 8260
rect 13740 8258 13746 8260
rect 13997 8258 14063 8261
rect 18873 8258 18939 8261
rect 13629 8200 13634 8256
rect 13629 8196 13676 8200
rect 13740 8198 13786 8258
rect 13997 8256 18939 8258
rect 13997 8200 14002 8256
rect 14058 8200 18878 8256
rect 18934 8200 18939 8256
rect 13997 8198 18939 8200
rect 13740 8196 13746 8198
rect 13629 8195 13695 8196
rect 13997 8195 14063 8198
rect 18873 8195 18939 8198
rect 19006 8196 19012 8260
rect 19076 8258 19082 8260
rect 19977 8258 20043 8261
rect 19076 8256 20043 8258
rect 19076 8200 19982 8256
rect 20038 8200 20043 8256
rect 19076 8198 20043 8200
rect 19076 8196 19082 8198
rect 19977 8195 20043 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 5349 8122 5415 8125
rect 7046 8122 7052 8124
rect 5349 8120 7052 8122
rect 5349 8064 5354 8120
rect 5410 8064 7052 8120
rect 5349 8062 7052 8064
rect 5349 8059 5415 8062
rect 7046 8060 7052 8062
rect 7116 8060 7122 8124
rect 9673 8122 9739 8125
rect 9857 8122 9923 8125
rect 17309 8124 17375 8125
rect 9673 8120 9923 8122
rect 9673 8064 9678 8120
rect 9734 8064 9862 8120
rect 9918 8064 9923 8120
rect 9673 8062 9923 8064
rect 9673 8059 9739 8062
rect 9857 8059 9923 8062
rect 9998 8062 17234 8122
rect 5809 7986 5875 7989
rect 9998 7986 10058 8062
rect 5809 7984 10058 7986
rect 5809 7928 5814 7984
rect 5870 7928 10058 7984
rect 5809 7926 10058 7928
rect 5809 7923 5875 7926
rect 12198 7924 12204 7988
rect 12268 7986 12274 7988
rect 12893 7986 12959 7989
rect 12268 7984 12959 7986
rect 12268 7928 12898 7984
rect 12954 7928 12959 7984
rect 12268 7926 12959 7928
rect 12268 7924 12274 7926
rect 12893 7923 12959 7926
rect 13261 7986 13327 7989
rect 16798 7986 16804 7988
rect 13261 7984 16804 7986
rect 13261 7928 13266 7984
rect 13322 7928 16804 7984
rect 13261 7926 16804 7928
rect 13261 7923 13327 7926
rect 16798 7924 16804 7926
rect 16868 7924 16874 7988
rect 17174 7986 17234 8062
rect 17309 8120 17356 8124
rect 17420 8122 17426 8124
rect 17769 8122 17835 8125
rect 20256 8122 20316 8334
rect 21817 8331 21883 8334
rect 22001 8394 22067 8397
rect 25681 8394 25747 8397
rect 22001 8392 25747 8394
rect 22001 8336 22006 8392
rect 22062 8336 25686 8392
rect 25742 8336 25747 8392
rect 22001 8334 25747 8336
rect 22001 8331 22067 8334
rect 25681 8331 25747 8334
rect 20713 8258 20779 8261
rect 23749 8258 23815 8261
rect 20713 8256 23815 8258
rect 20713 8200 20718 8256
rect 20774 8200 23754 8256
rect 23810 8200 23815 8256
rect 20713 8198 23815 8200
rect 20713 8195 20779 8198
rect 23749 8195 23815 8198
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 17309 8064 17314 8120
rect 17309 8060 17356 8064
rect 17420 8062 17466 8122
rect 17769 8120 20316 8122
rect 17769 8064 17774 8120
rect 17830 8064 20316 8120
rect 17769 8062 20316 8064
rect 17420 8060 17426 8062
rect 17309 8059 17375 8060
rect 17769 8059 17835 8062
rect 20662 8060 20668 8124
rect 20732 8122 20738 8124
rect 21173 8122 21239 8125
rect 21357 8122 21423 8125
rect 20732 8120 21423 8122
rect 20732 8064 21178 8120
rect 21234 8064 21362 8120
rect 21418 8064 21423 8120
rect 20732 8062 21423 8064
rect 20732 8060 20738 8062
rect 21173 8059 21239 8062
rect 21357 8059 21423 8062
rect 21541 8122 21607 8125
rect 24853 8122 24919 8125
rect 21541 8120 24919 8122
rect 21541 8064 21546 8120
rect 21602 8064 24858 8120
rect 24914 8064 24919 8120
rect 21541 8062 24919 8064
rect 21541 8059 21607 8062
rect 24853 8059 24919 8062
rect 22093 7986 22159 7989
rect 17174 7984 22159 7986
rect 17174 7928 22098 7984
rect 22154 7928 22159 7984
rect 17174 7926 22159 7928
rect 22093 7923 22159 7926
rect 22461 7986 22527 7989
rect 22829 7986 22895 7989
rect 22461 7984 22895 7986
rect 22461 7928 22466 7984
rect 22522 7928 22834 7984
rect 22890 7928 22895 7984
rect 22461 7926 22895 7928
rect 22461 7923 22527 7926
rect 22829 7923 22895 7926
rect 8661 7850 8727 7853
rect 9806 7850 9812 7852
rect 8661 7848 9812 7850
rect 8661 7792 8666 7848
rect 8722 7792 9812 7848
rect 8661 7790 9812 7792
rect 8661 7787 8727 7790
rect 9806 7788 9812 7790
rect 9876 7788 9882 7852
rect 10593 7850 10659 7853
rect 11278 7850 11284 7852
rect 10593 7848 11284 7850
rect 10593 7792 10598 7848
rect 10654 7792 11284 7848
rect 10593 7790 11284 7792
rect 10593 7787 10659 7790
rect 11278 7788 11284 7790
rect 11348 7850 11354 7852
rect 19057 7850 19123 7853
rect 11348 7848 19123 7850
rect 11348 7792 19062 7848
rect 19118 7792 19123 7848
rect 11348 7790 19123 7792
rect 11348 7788 11354 7790
rect 19057 7787 19123 7790
rect 19374 7788 19380 7852
rect 19444 7850 19450 7852
rect 20989 7850 21055 7853
rect 19444 7848 21055 7850
rect 19444 7792 20994 7848
rect 21050 7792 21055 7848
rect 19444 7790 21055 7792
rect 19444 7788 19450 7790
rect 20989 7787 21055 7790
rect 21398 7788 21404 7852
rect 21468 7850 21474 7852
rect 21909 7850 21975 7853
rect 21468 7848 21975 7850
rect 21468 7792 21914 7848
rect 21970 7792 21975 7848
rect 21468 7790 21975 7792
rect 21468 7788 21474 7790
rect 21909 7787 21975 7790
rect 8201 7714 8267 7717
rect 13813 7714 13879 7717
rect 8201 7712 13879 7714
rect 8201 7656 8206 7712
rect 8262 7656 13818 7712
rect 13874 7656 13879 7712
rect 8201 7654 13879 7656
rect 8201 7651 8267 7654
rect 13813 7651 13879 7654
rect 14457 7714 14523 7717
rect 16021 7714 16087 7717
rect 14457 7712 16087 7714
rect 14457 7656 14462 7712
rect 14518 7656 16026 7712
rect 16082 7656 16087 7712
rect 14457 7654 16087 7656
rect 14457 7651 14523 7654
rect 16021 7651 16087 7654
rect 16798 7652 16804 7716
rect 16868 7714 16874 7716
rect 17166 7714 17172 7716
rect 16868 7654 17172 7714
rect 16868 7652 16874 7654
rect 17166 7652 17172 7654
rect 17236 7652 17242 7716
rect 17718 7652 17724 7716
rect 17788 7714 17794 7716
rect 18321 7714 18387 7717
rect 17788 7712 18387 7714
rect 17788 7656 18326 7712
rect 18382 7656 18387 7712
rect 17788 7654 18387 7656
rect 17788 7652 17794 7654
rect 200 7578 800 7608
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 8753 7578 8819 7581
rect 8886 7578 8892 7580
rect 8753 7576 8892 7578
rect 8753 7520 8758 7576
rect 8814 7520 8892 7576
rect 8753 7518 8892 7520
rect 8753 7515 8819 7518
rect 8886 7516 8892 7518
rect 8956 7516 8962 7580
rect 9029 7578 9095 7581
rect 15561 7578 15627 7581
rect 9029 7576 15627 7578
rect 9029 7520 9034 7576
rect 9090 7520 15566 7576
rect 15622 7520 15627 7576
rect 9029 7518 15627 7520
rect 9029 7515 9095 7518
rect 15561 7515 15627 7518
rect 16614 7516 16620 7580
rect 16684 7578 16690 7580
rect 17033 7578 17099 7581
rect 16684 7576 17099 7578
rect 16684 7520 17038 7576
rect 17094 7520 17099 7576
rect 16684 7518 17099 7520
rect 17174 7578 17234 7652
rect 18321 7651 18387 7654
rect 18505 7714 18571 7717
rect 19425 7714 19491 7717
rect 18505 7712 19491 7714
rect 18505 7656 18510 7712
rect 18566 7656 19430 7712
rect 19486 7656 19491 7712
rect 18505 7654 19491 7656
rect 18505 7651 18571 7654
rect 19425 7651 19491 7654
rect 20713 7714 20779 7717
rect 24301 7714 24367 7717
rect 20713 7712 24367 7714
rect 20713 7656 20718 7712
rect 20774 7656 24306 7712
rect 24362 7656 24367 7712
rect 20713 7654 24367 7656
rect 20713 7651 20779 7654
rect 24301 7651 24367 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 19190 7578 19196 7580
rect 17174 7518 19196 7578
rect 16684 7516 16690 7518
rect 17033 7515 17099 7518
rect 19190 7516 19196 7518
rect 19260 7516 19266 7580
rect 20294 7516 20300 7580
rect 20364 7578 20370 7580
rect 24853 7578 24919 7581
rect 20364 7576 24919 7578
rect 20364 7520 24858 7576
rect 24914 7520 24919 7576
rect 20364 7518 24919 7520
rect 20364 7516 20370 7518
rect 24853 7515 24919 7518
rect 38285 7578 38351 7581
rect 39200 7578 39800 7608
rect 38285 7576 39800 7578
rect 38285 7520 38290 7576
rect 38346 7520 39800 7576
rect 38285 7518 39800 7520
rect 38285 7515 38351 7518
rect 39200 7488 39800 7518
rect 6453 7442 6519 7445
rect 7741 7442 7807 7445
rect 6453 7440 7807 7442
rect 6453 7384 6458 7440
rect 6514 7384 7746 7440
rect 7802 7384 7807 7440
rect 6453 7382 7807 7384
rect 6453 7379 6519 7382
rect 7741 7379 7807 7382
rect 7925 7442 7991 7445
rect 22645 7442 22711 7445
rect 7925 7440 22711 7442
rect 7925 7384 7930 7440
rect 7986 7384 22650 7440
rect 22706 7384 22711 7440
rect 7925 7382 22711 7384
rect 7925 7379 7991 7382
rect 22645 7379 22711 7382
rect 4061 7306 4127 7309
rect 17309 7306 17375 7309
rect 21725 7306 21791 7309
rect 4061 7304 17375 7306
rect 4061 7248 4066 7304
rect 4122 7248 17314 7304
rect 17370 7248 17375 7304
rect 4061 7246 17375 7248
rect 4061 7243 4127 7246
rect 17309 7243 17375 7246
rect 17496 7304 21791 7306
rect 17496 7248 21730 7304
rect 21786 7248 21791 7304
rect 17496 7246 21791 7248
rect 9673 7170 9739 7173
rect 13813 7170 13879 7173
rect 9673 7168 13879 7170
rect 9673 7112 9678 7168
rect 9734 7112 13818 7168
rect 13874 7112 13879 7168
rect 9673 7110 13879 7112
rect 9673 7107 9739 7110
rect 13813 7107 13879 7110
rect 14181 7170 14247 7173
rect 14825 7170 14891 7173
rect 14181 7168 14891 7170
rect 14181 7112 14186 7168
rect 14242 7112 14830 7168
rect 14886 7112 14891 7168
rect 14181 7110 14891 7112
rect 14181 7107 14247 7110
rect 14825 7107 14891 7110
rect 15193 7170 15259 7173
rect 17496 7170 17556 7246
rect 21725 7243 21791 7246
rect 22134 7244 22140 7308
rect 22204 7306 22210 7308
rect 22277 7306 22343 7309
rect 22204 7304 22343 7306
rect 22204 7248 22282 7304
rect 22338 7248 22343 7304
rect 22204 7246 22343 7248
rect 22204 7244 22210 7246
rect 22277 7243 22343 7246
rect 15193 7168 17556 7170
rect 15193 7112 15198 7168
rect 15254 7112 17556 7168
rect 15193 7110 17556 7112
rect 17953 7170 18019 7173
rect 22502 7170 22508 7172
rect 17953 7168 22508 7170
rect 17953 7112 17958 7168
rect 18014 7112 22508 7168
rect 17953 7110 22508 7112
rect 15193 7107 15259 7110
rect 17953 7107 18019 7110
rect 22502 7108 22508 7110
rect 22572 7170 22578 7172
rect 24669 7170 24735 7173
rect 22572 7168 24735 7170
rect 22572 7112 24674 7168
rect 24730 7112 24735 7168
rect 22572 7110 24735 7112
rect 22572 7108 22578 7110
rect 24669 7107 24735 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 7465 7034 7531 7037
rect 10409 7036 10475 7037
rect 9806 7034 9812 7036
rect 7465 7032 9812 7034
rect 7465 6976 7470 7032
rect 7526 6976 9812 7032
rect 7465 6974 9812 6976
rect 7465 6971 7531 6974
rect 9806 6972 9812 6974
rect 9876 6972 9882 7036
rect 10358 7034 10364 7036
rect 10318 6974 10364 7034
rect 10428 7032 10475 7036
rect 10869 7036 10935 7037
rect 10869 7034 10916 7036
rect 10470 6976 10475 7032
rect 10358 6972 10364 6974
rect 10428 6972 10475 6976
rect 10824 7032 10916 7034
rect 10824 6976 10874 7032
rect 10824 6974 10916 6976
rect 10409 6971 10475 6972
rect 10869 6972 10916 6974
rect 10980 6972 10986 7036
rect 11053 7034 11119 7037
rect 11646 7034 11652 7036
rect 11053 7032 11652 7034
rect 11053 6976 11058 7032
rect 11114 6976 11652 7032
rect 11053 6974 11652 6976
rect 10869 6971 10935 6972
rect 11053 6971 11119 6974
rect 11646 6972 11652 6974
rect 11716 6972 11722 7036
rect 11881 7034 11947 7037
rect 15469 7034 15535 7037
rect 11881 7032 15535 7034
rect 11881 6976 11886 7032
rect 11942 6976 15474 7032
rect 15530 6976 15535 7032
rect 11881 6974 15535 6976
rect 11881 6971 11947 6974
rect 15469 6971 15535 6974
rect 15653 7034 15719 7037
rect 18597 7036 18663 7037
rect 18454 7034 18460 7036
rect 15653 7032 18460 7034
rect 15653 6976 15658 7032
rect 15714 6976 18460 7032
rect 15653 6974 18460 6976
rect 15653 6971 15719 6974
rect 18454 6972 18460 6974
rect 18524 6972 18530 7036
rect 18597 7032 18644 7036
rect 18708 7034 18714 7036
rect 18597 6976 18602 7032
rect 18597 6972 18644 6976
rect 18708 6974 18754 7034
rect 18708 6972 18714 6974
rect 19190 6972 19196 7036
rect 19260 7034 19266 7036
rect 19977 7034 20043 7037
rect 19260 7032 20043 7034
rect 19260 6976 19982 7032
rect 20038 6976 20043 7032
rect 19260 6974 20043 6976
rect 19260 6972 19266 6974
rect 18597 6971 18663 6972
rect 19977 6971 20043 6974
rect 20294 6972 20300 7036
rect 20364 7034 20370 7036
rect 22093 7034 22159 7037
rect 20364 7032 22159 7034
rect 20364 6976 22098 7032
rect 22154 6976 22159 7032
rect 20364 6974 22159 6976
rect 20364 6972 20370 6974
rect 22093 6971 22159 6974
rect 12617 6898 12683 6901
rect 6502 6896 12683 6898
rect 6502 6840 12622 6896
rect 12678 6840 12683 6896
rect 6502 6838 12683 6840
rect 2313 6490 2379 6493
rect 5574 6490 5580 6492
rect 2313 6488 5580 6490
rect 2313 6432 2318 6488
rect 2374 6432 5580 6488
rect 2313 6430 5580 6432
rect 2313 6427 2379 6430
rect 5574 6428 5580 6430
rect 5644 6428 5650 6492
rect 2313 6354 2379 6357
rect 6502 6354 6562 6838
rect 12617 6835 12683 6838
rect 12801 6898 12867 6901
rect 15193 6898 15259 6901
rect 12801 6896 15259 6898
rect 12801 6840 12806 6896
rect 12862 6840 15198 6896
rect 15254 6840 15259 6896
rect 12801 6838 15259 6840
rect 12801 6835 12867 6838
rect 15193 6835 15259 6838
rect 15694 6836 15700 6900
rect 15764 6898 15770 6900
rect 22001 6898 22067 6901
rect 15764 6896 22067 6898
rect 15764 6840 22006 6896
rect 22062 6840 22067 6896
rect 15764 6838 22067 6840
rect 15764 6836 15770 6838
rect 22001 6835 22067 6838
rect 23054 6836 23060 6900
rect 23124 6898 23130 6900
rect 23381 6898 23447 6901
rect 24669 6900 24735 6901
rect 24669 6898 24716 6900
rect 23124 6896 23447 6898
rect 23124 6840 23386 6896
rect 23442 6840 23447 6896
rect 23124 6838 23447 6840
rect 24624 6896 24716 6898
rect 24624 6840 24674 6896
rect 24624 6838 24716 6840
rect 23124 6836 23130 6838
rect 23381 6835 23447 6838
rect 24669 6836 24716 6838
rect 24780 6836 24786 6900
rect 38101 6898 38167 6901
rect 39200 6898 39800 6928
rect 38101 6896 39800 6898
rect 38101 6840 38106 6896
rect 38162 6840 39800 6896
rect 38101 6838 39800 6840
rect 24669 6835 24735 6836
rect 38101 6835 38167 6838
rect 39200 6808 39800 6838
rect 9029 6762 9095 6765
rect 9029 6760 10840 6762
rect 9029 6704 9034 6760
rect 9090 6728 10840 6760
rect 9090 6704 11116 6728
rect 9029 6702 11116 6704
rect 9029 6699 9095 6702
rect 10780 6668 11116 6702
rect 12198 6700 12204 6764
rect 12268 6762 12274 6764
rect 17861 6762 17927 6765
rect 12268 6760 17927 6762
rect 12268 6704 17866 6760
rect 17922 6704 17927 6760
rect 12268 6702 17927 6704
rect 12268 6700 12274 6702
rect 17861 6699 17927 6702
rect 18270 6700 18276 6764
rect 18340 6762 18346 6764
rect 18413 6762 18479 6765
rect 18340 6760 18479 6762
rect 18340 6704 18418 6760
rect 18474 6704 18479 6760
rect 18340 6702 18479 6704
rect 18340 6700 18346 6702
rect 18413 6699 18479 6702
rect 18638 6700 18644 6764
rect 18708 6762 18714 6764
rect 20846 6762 20852 6764
rect 18708 6702 20852 6762
rect 18708 6700 18714 6702
rect 9121 6626 9187 6629
rect 9489 6626 9555 6629
rect 9121 6624 9555 6626
rect 9121 6568 9126 6624
rect 9182 6568 9494 6624
rect 9550 6568 9555 6624
rect 9121 6566 9555 6568
rect 9121 6563 9187 6566
rect 9489 6563 9555 6566
rect 10041 6626 10107 6629
rect 10409 6626 10475 6629
rect 10041 6624 10475 6626
rect 10041 6568 10046 6624
rect 10102 6568 10414 6624
rect 10470 6568 10475 6624
rect 10041 6566 10475 6568
rect 11056 6626 11116 6668
rect 19060 6629 19120 6702
rect 20846 6700 20852 6702
rect 20916 6700 20922 6764
rect 21081 6762 21147 6765
rect 22318 6762 22324 6764
rect 21081 6760 22324 6762
rect 21081 6704 21086 6760
rect 21142 6704 22324 6760
rect 21081 6702 22324 6704
rect 21081 6699 21147 6702
rect 22318 6700 22324 6702
rect 22388 6700 22394 6764
rect 12157 6626 12223 6629
rect 11056 6624 12223 6626
rect 11056 6568 12162 6624
rect 12218 6568 12223 6624
rect 11056 6566 12223 6568
rect 10041 6563 10107 6566
rect 10409 6563 10475 6566
rect 12157 6563 12223 6566
rect 12382 6564 12388 6628
rect 12452 6626 12458 6628
rect 15193 6626 15259 6629
rect 12452 6624 15259 6626
rect 12452 6568 15198 6624
rect 15254 6568 15259 6624
rect 12452 6566 15259 6568
rect 12452 6564 12458 6566
rect 15193 6563 15259 6566
rect 15469 6626 15535 6629
rect 16573 6626 16639 6629
rect 15469 6624 16639 6626
rect 15469 6568 15474 6624
rect 15530 6568 16578 6624
rect 16634 6568 16639 6624
rect 15469 6566 16639 6568
rect 15469 6563 15535 6566
rect 16573 6563 16639 6566
rect 16757 6626 16823 6629
rect 17493 6626 17559 6629
rect 16757 6624 17559 6626
rect 16757 6568 16762 6624
rect 16818 6568 17498 6624
rect 17554 6568 17559 6624
rect 16757 6566 17559 6568
rect 16757 6563 16823 6566
rect 17493 6563 17559 6566
rect 17718 6564 17724 6628
rect 17788 6626 17794 6628
rect 18597 6626 18663 6629
rect 17788 6624 18663 6626
rect 17788 6568 18602 6624
rect 18658 6568 18663 6624
rect 17788 6566 18663 6568
rect 17788 6564 17794 6566
rect 18597 6563 18663 6566
rect 19057 6624 19123 6629
rect 19057 6568 19062 6624
rect 19118 6568 19123 6624
rect 19057 6563 19123 6568
rect 20110 6564 20116 6628
rect 20180 6626 20186 6628
rect 20621 6626 20687 6629
rect 20180 6624 20687 6626
rect 20180 6568 20626 6624
rect 20682 6568 20687 6624
rect 20180 6566 20687 6568
rect 20180 6564 20186 6566
rect 20621 6563 20687 6566
rect 21214 6564 21220 6628
rect 21284 6626 21290 6628
rect 23565 6626 23631 6629
rect 21284 6624 23631 6626
rect 21284 6568 23570 6624
rect 23626 6568 23631 6624
rect 21284 6566 23631 6568
rect 21284 6564 21290 6566
rect 23565 6563 23631 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 6821 6490 6887 6493
rect 17953 6490 18019 6493
rect 6821 6488 18019 6490
rect 6821 6432 6826 6488
rect 6882 6432 17958 6488
rect 18014 6432 18019 6488
rect 6821 6430 18019 6432
rect 6821 6427 6887 6430
rect 17953 6427 18019 6430
rect 18781 6490 18847 6493
rect 19006 6490 19012 6492
rect 18781 6488 19012 6490
rect 18781 6432 18786 6488
rect 18842 6432 19012 6488
rect 18781 6430 19012 6432
rect 18781 6427 18847 6430
rect 19006 6428 19012 6430
rect 19076 6428 19082 6492
rect 20805 6490 20871 6493
rect 19980 6488 20871 6490
rect 19980 6432 20810 6488
rect 20866 6432 20871 6488
rect 19980 6430 20871 6432
rect 2313 6352 6562 6354
rect 2313 6296 2318 6352
rect 2374 6296 6562 6352
rect 2313 6294 6562 6296
rect 9305 6354 9371 6357
rect 9990 6354 9996 6356
rect 9305 6352 9996 6354
rect 9305 6296 9310 6352
rect 9366 6296 9996 6352
rect 9305 6294 9996 6296
rect 2313 6291 2379 6294
rect 9305 6291 9371 6294
rect 9990 6292 9996 6294
rect 10060 6292 10066 6356
rect 10358 6292 10364 6356
rect 10428 6354 10434 6356
rect 10593 6354 10659 6357
rect 10428 6352 10659 6354
rect 10428 6296 10598 6352
rect 10654 6296 10659 6352
rect 10428 6294 10659 6296
rect 10428 6292 10434 6294
rect 10593 6291 10659 6294
rect 10777 6354 10843 6357
rect 13997 6354 14063 6357
rect 10777 6352 14063 6354
rect 10777 6296 10782 6352
rect 10838 6296 14002 6352
rect 14058 6296 14063 6352
rect 10777 6294 14063 6296
rect 10777 6291 10843 6294
rect 13997 6291 14063 6294
rect 14641 6354 14707 6357
rect 15653 6354 15719 6357
rect 14641 6352 15719 6354
rect 14641 6296 14646 6352
rect 14702 6296 15658 6352
rect 15714 6296 15719 6352
rect 14641 6294 15719 6296
rect 14641 6291 14707 6294
rect 15653 6291 15719 6294
rect 16849 6354 16915 6357
rect 17493 6354 17559 6357
rect 16849 6352 17559 6354
rect 16849 6296 16854 6352
rect 16910 6296 17498 6352
rect 17554 6296 17559 6352
rect 16849 6294 17559 6296
rect 16849 6291 16915 6294
rect 17493 6291 17559 6294
rect 17902 6292 17908 6356
rect 17972 6354 17978 6356
rect 19609 6354 19675 6357
rect 17972 6352 19675 6354
rect 17972 6296 19614 6352
rect 19670 6296 19675 6352
rect 17972 6294 19675 6296
rect 17972 6292 17978 6294
rect 19609 6291 19675 6294
rect 19793 6354 19859 6357
rect 19980 6354 20040 6430
rect 20805 6427 20871 6430
rect 21030 6428 21036 6492
rect 21100 6490 21106 6492
rect 22277 6490 22343 6493
rect 21100 6488 22343 6490
rect 21100 6432 22282 6488
rect 22338 6432 22343 6488
rect 21100 6430 22343 6432
rect 21100 6428 21106 6430
rect 22277 6427 22343 6430
rect 19793 6352 20040 6354
rect 19793 6296 19798 6352
rect 19854 6296 20040 6352
rect 19793 6294 20040 6296
rect 20253 6354 20319 6357
rect 22921 6354 22987 6357
rect 20253 6352 22987 6354
rect 20253 6296 20258 6352
rect 20314 6296 22926 6352
rect 22982 6296 22987 6352
rect 20253 6294 22987 6296
rect 19793 6291 19859 6294
rect 20253 6291 20319 6294
rect 22921 6291 22987 6294
rect 200 6218 800 6248
rect 3693 6218 3759 6221
rect 200 6216 3759 6218
rect 200 6160 3698 6216
rect 3754 6160 3759 6216
rect 200 6158 3759 6160
rect 200 6128 800 6158
rect 3693 6155 3759 6158
rect 5717 6218 5783 6221
rect 10358 6218 10364 6220
rect 5717 6216 10364 6218
rect 5717 6160 5722 6216
rect 5778 6160 10364 6216
rect 5717 6158 10364 6160
rect 5717 6155 5783 6158
rect 10358 6156 10364 6158
rect 10428 6156 10434 6220
rect 10542 6156 10548 6220
rect 10612 6218 10618 6220
rect 21357 6218 21423 6221
rect 22369 6218 22435 6221
rect 10612 6216 21423 6218
rect 10612 6160 21362 6216
rect 21418 6160 21423 6216
rect 10612 6158 21423 6160
rect 10612 6156 10618 6158
rect 21357 6155 21423 6158
rect 21590 6216 22435 6218
rect 21590 6160 22374 6216
rect 22430 6160 22435 6216
rect 21590 6158 22435 6160
rect 4797 6082 4863 6085
rect 15510 6082 15516 6084
rect 4797 6080 15516 6082
rect 4797 6024 4802 6080
rect 4858 6024 15516 6080
rect 4797 6022 15516 6024
rect 4797 6019 4863 6022
rect 15510 6020 15516 6022
rect 15580 6020 15586 6084
rect 21590 6082 21650 6158
rect 22369 6155 22435 6158
rect 16806 6022 21650 6082
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4705 5946 4771 5949
rect 12198 5946 12204 5948
rect 4705 5944 12204 5946
rect 4705 5888 4710 5944
rect 4766 5888 12204 5944
rect 4705 5886 12204 5888
rect 4705 5883 4771 5886
rect 12198 5884 12204 5886
rect 12268 5884 12274 5948
rect 12382 5884 12388 5948
rect 12452 5946 12458 5948
rect 16806 5946 16866 6022
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 17033 5948 17099 5949
rect 12452 5886 16866 5946
rect 12452 5884 12458 5886
rect 16982 5884 16988 5948
rect 17052 5946 17099 5948
rect 18045 5946 18111 5949
rect 24025 5946 24091 5949
rect 17052 5944 17144 5946
rect 17094 5888 17144 5944
rect 17052 5886 17144 5888
rect 18045 5944 24091 5946
rect 18045 5888 18050 5944
rect 18106 5888 24030 5944
rect 24086 5888 24091 5944
rect 18045 5886 24091 5888
rect 17052 5884 17099 5886
rect 17033 5883 17099 5884
rect 18045 5883 18111 5886
rect 24025 5883 24091 5886
rect 8661 5810 8727 5813
rect 13077 5810 13143 5813
rect 8661 5808 13143 5810
rect 8661 5752 8666 5808
rect 8722 5752 13082 5808
rect 13138 5752 13143 5808
rect 8661 5750 13143 5752
rect 8661 5747 8727 5750
rect 13077 5747 13143 5750
rect 13353 5810 13419 5813
rect 17493 5810 17559 5813
rect 13353 5808 17559 5810
rect 13353 5752 13358 5808
rect 13414 5752 17498 5808
rect 17554 5752 17559 5808
rect 13353 5750 17559 5752
rect 13353 5747 13419 5750
rect 17493 5747 17559 5750
rect 18229 5810 18295 5813
rect 19425 5810 19491 5813
rect 18229 5808 19491 5810
rect 18229 5752 18234 5808
rect 18290 5752 19430 5808
rect 19486 5752 19491 5808
rect 18229 5750 19491 5752
rect 18229 5747 18295 5750
rect 19425 5747 19491 5750
rect 19977 5810 20043 5813
rect 20989 5810 21055 5813
rect 19977 5808 21055 5810
rect 19977 5752 19982 5808
rect 20038 5752 20994 5808
rect 21050 5752 21055 5808
rect 19977 5750 21055 5752
rect 19977 5747 20043 5750
rect 20989 5747 21055 5750
rect 21173 5810 21239 5813
rect 22461 5810 22527 5813
rect 21173 5808 22527 5810
rect 21173 5752 21178 5808
rect 21234 5752 22466 5808
rect 22522 5752 22527 5808
rect 21173 5750 22527 5752
rect 21173 5747 21239 5750
rect 22461 5747 22527 5750
rect 6453 5674 6519 5677
rect 6913 5674 6979 5677
rect 6453 5672 6979 5674
rect 6453 5616 6458 5672
rect 6514 5616 6918 5672
rect 6974 5616 6979 5672
rect 6453 5614 6979 5616
rect 6453 5611 6519 5614
rect 6913 5611 6979 5614
rect 8109 5674 8175 5677
rect 11237 5674 11303 5677
rect 12198 5674 12204 5676
rect 8109 5672 11303 5674
rect 8109 5616 8114 5672
rect 8170 5616 11242 5672
rect 11298 5616 11303 5672
rect 8109 5614 11303 5616
rect 8109 5611 8175 5614
rect 11237 5611 11303 5614
rect 11470 5614 12204 5674
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 5073 5538 5139 5541
rect 10174 5538 10180 5540
rect 5073 5536 10180 5538
rect 5073 5480 5078 5536
rect 5134 5480 10180 5536
rect 5073 5478 10180 5480
rect 5073 5475 5139 5478
rect 10174 5476 10180 5478
rect 10244 5476 10250 5540
rect 10317 5538 10383 5541
rect 10542 5538 10548 5540
rect 10317 5536 10548 5538
rect 10317 5480 10322 5536
rect 10378 5480 10548 5536
rect 10317 5478 10548 5480
rect 10317 5475 10383 5478
rect 10542 5476 10548 5478
rect 10612 5476 10618 5540
rect 11470 5538 11530 5614
rect 12198 5612 12204 5614
rect 12268 5612 12274 5676
rect 12341 5674 12407 5677
rect 12525 5674 12591 5677
rect 12341 5672 12591 5674
rect 12341 5616 12346 5672
rect 12402 5616 12530 5672
rect 12586 5616 12591 5672
rect 12341 5614 12591 5616
rect 12341 5611 12407 5614
rect 12525 5611 12591 5614
rect 12750 5612 12756 5676
rect 12820 5674 12826 5676
rect 15377 5674 15443 5677
rect 12820 5672 15443 5674
rect 12820 5616 15382 5672
rect 15438 5616 15443 5672
rect 12820 5614 15443 5616
rect 12820 5612 12826 5614
rect 15377 5611 15443 5614
rect 16389 5674 16455 5677
rect 17718 5674 17724 5676
rect 16389 5672 17724 5674
rect 16389 5616 16394 5672
rect 16450 5616 17724 5672
rect 16389 5614 17724 5616
rect 16389 5611 16455 5614
rect 17718 5612 17724 5614
rect 17788 5612 17794 5676
rect 18086 5612 18092 5676
rect 18156 5674 18162 5676
rect 20805 5674 20871 5677
rect 27654 5674 27660 5676
rect 18156 5672 20871 5674
rect 18156 5616 20810 5672
rect 20866 5616 20871 5672
rect 18156 5614 20871 5616
rect 18156 5612 18162 5614
rect 20805 5611 20871 5614
rect 22050 5614 27660 5674
rect 10734 5478 11530 5538
rect 11605 5538 11671 5541
rect 13077 5538 13143 5541
rect 13997 5540 14063 5541
rect 13854 5538 13860 5540
rect 11605 5536 13002 5538
rect 11605 5480 11610 5536
rect 11666 5480 13002 5536
rect 11605 5478 13002 5480
rect 6085 5402 6151 5405
rect 7097 5402 7163 5405
rect 8477 5404 8543 5405
rect 8477 5402 8524 5404
rect 6085 5400 7163 5402
rect 6085 5344 6090 5400
rect 6146 5344 7102 5400
rect 7158 5344 7163 5400
rect 6085 5342 7163 5344
rect 8432 5400 8524 5402
rect 8432 5344 8482 5400
rect 8432 5342 8524 5344
rect 6085 5339 6151 5342
rect 7097 5339 7163 5342
rect 8477 5340 8524 5342
rect 8588 5340 8594 5404
rect 8661 5402 8727 5405
rect 10041 5402 10107 5405
rect 8661 5400 10107 5402
rect 8661 5344 8666 5400
rect 8722 5344 10046 5400
rect 10102 5344 10107 5400
rect 8661 5342 10107 5344
rect 8477 5339 8543 5340
rect 8661 5339 8727 5342
rect 10041 5339 10107 5342
rect 10358 5340 10364 5404
rect 10428 5402 10434 5404
rect 10734 5402 10794 5478
rect 11605 5475 11671 5478
rect 12525 5402 12591 5405
rect 10428 5342 10794 5402
rect 10872 5400 12591 5402
rect 10872 5344 12530 5400
rect 12586 5344 12591 5400
rect 10872 5342 12591 5344
rect 12942 5402 13002 5478
rect 13077 5536 13860 5538
rect 13077 5480 13082 5536
rect 13138 5480 13860 5536
rect 13077 5478 13860 5480
rect 13077 5475 13143 5478
rect 13854 5476 13860 5478
rect 13924 5476 13930 5540
rect 13997 5536 14044 5540
rect 14108 5538 14114 5540
rect 15193 5538 15259 5541
rect 15653 5538 15719 5541
rect 16113 5538 16179 5541
rect 13997 5480 14002 5536
rect 13997 5476 14044 5480
rect 14108 5478 14154 5538
rect 15193 5536 15394 5538
rect 15193 5480 15198 5536
rect 15254 5480 15394 5536
rect 15193 5478 15394 5480
rect 14108 5476 14114 5478
rect 13997 5475 14063 5476
rect 15193 5475 15259 5478
rect 15193 5402 15259 5405
rect 12942 5400 15259 5402
rect 12942 5344 15198 5400
rect 15254 5344 15259 5400
rect 12942 5342 15259 5344
rect 15334 5402 15394 5478
rect 15653 5536 16179 5538
rect 15653 5480 15658 5536
rect 15714 5480 16118 5536
rect 16174 5480 16179 5536
rect 15653 5478 16179 5480
rect 15653 5475 15719 5478
rect 16113 5475 16179 5478
rect 16481 5538 16547 5541
rect 19057 5538 19123 5541
rect 16481 5536 19123 5538
rect 16481 5480 16486 5536
rect 16542 5480 19062 5536
rect 19118 5480 19123 5536
rect 16481 5478 19123 5480
rect 16481 5475 16547 5478
rect 19057 5475 19123 5478
rect 20713 5538 20779 5541
rect 22050 5538 22110 5614
rect 27654 5612 27660 5614
rect 27724 5612 27730 5676
rect 20713 5536 22110 5538
rect 20713 5480 20718 5536
rect 20774 5480 22110 5536
rect 20713 5478 22110 5480
rect 24853 5538 24919 5541
rect 26918 5538 26924 5540
rect 24853 5536 26924 5538
rect 24853 5480 24858 5536
rect 24914 5480 26924 5536
rect 24853 5478 26924 5480
rect 20713 5475 20779 5478
rect 24853 5475 24919 5478
rect 26918 5476 26924 5478
rect 26988 5476 26994 5540
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 17493 5402 17559 5405
rect 18689 5402 18755 5405
rect 18822 5402 18828 5404
rect 15334 5342 17050 5402
rect 10428 5340 10434 5342
rect 7281 5266 7347 5269
rect 10872 5266 10932 5342
rect 12525 5339 12591 5342
rect 15193 5339 15259 5342
rect 7281 5264 10932 5266
rect 7281 5208 7286 5264
rect 7342 5208 10932 5264
rect 7281 5206 10932 5208
rect 11237 5266 11303 5269
rect 16757 5266 16823 5269
rect 11237 5264 16823 5266
rect 11237 5208 11242 5264
rect 11298 5208 16762 5264
rect 16818 5208 16823 5264
rect 11237 5206 16823 5208
rect 16990 5266 17050 5342
rect 17493 5400 18828 5402
rect 17493 5344 17498 5400
rect 17554 5344 18694 5400
rect 18750 5344 18828 5400
rect 17493 5342 18828 5344
rect 17493 5339 17559 5342
rect 18689 5339 18755 5342
rect 18822 5340 18828 5342
rect 18892 5340 18898 5404
rect 19977 5402 20043 5405
rect 20897 5402 20963 5405
rect 19977 5400 20963 5402
rect 19977 5344 19982 5400
rect 20038 5344 20902 5400
rect 20958 5344 20963 5400
rect 19977 5342 20963 5344
rect 19977 5339 20043 5342
rect 20897 5339 20963 5342
rect 20805 5266 20871 5269
rect 16990 5264 20871 5266
rect 16990 5208 20810 5264
rect 20866 5208 20871 5264
rect 16990 5206 20871 5208
rect 7281 5203 7347 5206
rect 11237 5203 11303 5206
rect 16757 5203 16823 5206
rect 20805 5203 20871 5206
rect 3877 5130 3943 5133
rect 11697 5130 11763 5133
rect 18137 5130 18203 5133
rect 3877 5128 11763 5130
rect 3877 5072 3882 5128
rect 3938 5072 11702 5128
rect 11758 5072 11763 5128
rect 3877 5070 11763 5072
rect 3877 5067 3943 5070
rect 11697 5067 11763 5070
rect 11838 5128 18203 5130
rect 11838 5072 18142 5128
rect 18198 5072 18203 5128
rect 11838 5070 18203 5072
rect 7046 4932 7052 4996
rect 7116 4994 7122 4996
rect 8845 4994 8911 4997
rect 9765 4994 9831 4997
rect 7116 4992 8911 4994
rect 7116 4936 8850 4992
rect 8906 4936 8911 4992
rect 7116 4934 8911 4936
rect 7116 4932 7122 4934
rect 8845 4931 8911 4934
rect 9032 4992 9831 4994
rect 9032 4936 9770 4992
rect 9826 4936 9831 4992
rect 9032 4934 9831 4936
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 8293 4858 8359 4861
rect 9032 4858 9092 4934
rect 9765 4931 9831 4934
rect 10174 4932 10180 4996
rect 10244 4994 10250 4996
rect 11838 4994 11898 5070
rect 18137 5067 18203 5070
rect 18270 5068 18276 5132
rect 18340 5130 18346 5132
rect 23105 5130 23171 5133
rect 18340 5128 23171 5130
rect 18340 5072 23110 5128
rect 23166 5072 23171 5128
rect 18340 5070 23171 5072
rect 18340 5068 18346 5070
rect 23105 5067 23171 5070
rect 10244 4934 11898 4994
rect 10244 4932 10250 4934
rect 12014 4932 12020 4996
rect 12084 4994 12090 4996
rect 17493 4994 17559 4997
rect 22277 4994 22343 4997
rect 12084 4992 17559 4994
rect 12084 4936 17498 4992
rect 17554 4936 17559 4992
rect 12084 4934 17559 4936
rect 12084 4932 12090 4934
rect 17493 4931 17559 4934
rect 17726 4992 22343 4994
rect 17726 4936 22282 4992
rect 22338 4936 22343 4992
rect 17726 4934 22343 4936
rect 8293 4856 9092 4858
rect 8293 4800 8298 4856
rect 8354 4800 9092 4856
rect 8293 4798 9092 4800
rect 8293 4795 8359 4798
rect 9254 4796 9260 4860
rect 9324 4858 9330 4860
rect 9673 4858 9739 4861
rect 9324 4856 9739 4858
rect 9324 4800 9678 4856
rect 9734 4800 9739 4856
rect 9324 4798 9739 4800
rect 9324 4796 9330 4798
rect 9673 4795 9739 4798
rect 9990 4796 9996 4860
rect 10060 4858 10066 4860
rect 12525 4858 12591 4861
rect 13118 4858 13124 4860
rect 10060 4856 13124 4858
rect 10060 4800 12530 4856
rect 12586 4800 13124 4856
rect 10060 4798 13124 4800
rect 10060 4796 10066 4798
rect 12525 4795 12591 4798
rect 13118 4796 13124 4798
rect 13188 4796 13194 4860
rect 13445 4858 13511 4861
rect 13264 4856 13511 4858
rect 13264 4800 13450 4856
rect 13506 4800 13511 4856
rect 13264 4798 13511 4800
rect 2078 4660 2084 4724
rect 2148 4722 2154 4724
rect 4705 4722 4771 4725
rect 2148 4720 4771 4722
rect 2148 4664 4710 4720
rect 4766 4664 4771 4720
rect 2148 4662 4771 4664
rect 2148 4660 2154 4662
rect 4705 4659 4771 4662
rect 7741 4722 7807 4725
rect 12065 4722 12131 4725
rect 7741 4720 12131 4722
rect 7741 4664 7746 4720
rect 7802 4664 12070 4720
rect 12126 4664 12131 4720
rect 7741 4662 12131 4664
rect 7741 4659 7807 4662
rect 12065 4659 12131 4662
rect 12341 4724 12407 4725
rect 12341 4720 12388 4724
rect 12452 4722 12458 4724
rect 12341 4664 12346 4720
rect 12341 4660 12388 4664
rect 12452 4662 12498 4722
rect 12452 4660 12458 4662
rect 12566 4660 12572 4724
rect 12636 4722 12642 4724
rect 13264 4722 13324 4798
rect 13445 4795 13511 4798
rect 13721 4858 13787 4861
rect 14181 4858 14247 4861
rect 13721 4856 14247 4858
rect 13721 4800 13726 4856
rect 13782 4800 14186 4856
rect 14242 4800 14247 4856
rect 13721 4798 14247 4800
rect 13721 4795 13787 4798
rect 14181 4795 14247 4798
rect 14641 4858 14707 4861
rect 14774 4858 14780 4860
rect 14641 4856 14780 4858
rect 14641 4800 14646 4856
rect 14702 4800 14780 4856
rect 14641 4798 14780 4800
rect 14641 4795 14707 4798
rect 14774 4796 14780 4798
rect 14844 4796 14850 4860
rect 15193 4858 15259 4861
rect 17726 4858 17786 4934
rect 22277 4931 22343 4934
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 15193 4856 17786 4858
rect 15193 4800 15198 4856
rect 15254 4800 17786 4856
rect 15193 4798 17786 4800
rect 17953 4858 18019 4861
rect 22093 4858 22159 4861
rect 17953 4856 22159 4858
rect 17953 4800 17958 4856
rect 18014 4800 22098 4856
rect 22154 4800 22159 4856
rect 17953 4798 22159 4800
rect 15193 4795 15259 4798
rect 17953 4795 18019 4798
rect 22093 4795 22159 4798
rect 38193 4858 38259 4861
rect 39200 4858 39800 4888
rect 38193 4856 39800 4858
rect 38193 4800 38198 4856
rect 38254 4800 39800 4856
rect 38193 4798 39800 4800
rect 38193 4795 38259 4798
rect 39200 4768 39800 4798
rect 12636 4662 13324 4722
rect 12636 4660 12642 4662
rect 13486 4660 13492 4724
rect 13556 4722 13562 4724
rect 15285 4722 15351 4725
rect 13556 4720 15351 4722
rect 13556 4664 15290 4720
rect 15346 4664 15351 4720
rect 13556 4662 15351 4664
rect 13556 4660 13562 4662
rect 12341 4659 12407 4660
rect 15285 4659 15351 4662
rect 15694 4660 15700 4724
rect 15764 4722 15770 4724
rect 16665 4722 16731 4725
rect 15764 4720 16731 4722
rect 15764 4664 16670 4720
rect 16726 4664 16731 4720
rect 15764 4662 16731 4664
rect 15764 4660 15770 4662
rect 16665 4659 16731 4662
rect 17350 4660 17356 4724
rect 17420 4722 17426 4724
rect 21357 4722 21423 4725
rect 17420 4720 21423 4722
rect 17420 4664 21362 4720
rect 21418 4664 21423 4720
rect 17420 4662 21423 4664
rect 17420 4660 17426 4662
rect 21357 4659 21423 4662
rect 7281 4586 7347 4589
rect 20713 4586 20779 4589
rect 7281 4584 20779 4586
rect 7281 4528 7286 4584
rect 7342 4528 20718 4584
rect 20774 4528 20779 4584
rect 7281 4526 20779 4528
rect 7281 4523 7347 4526
rect 20713 4523 20779 4526
rect 7005 4450 7071 4453
rect 13721 4450 13787 4453
rect 7005 4448 13787 4450
rect 7005 4392 7010 4448
rect 7066 4392 13726 4448
rect 13782 4392 13787 4448
rect 7005 4390 13787 4392
rect 7005 4387 7071 4390
rect 13721 4387 13787 4390
rect 15101 4450 15167 4453
rect 15694 4450 15700 4452
rect 15101 4448 15700 4450
rect 15101 4392 15106 4448
rect 15162 4392 15700 4448
rect 15101 4390 15700 4392
rect 15101 4387 15167 4390
rect 15694 4388 15700 4390
rect 15764 4388 15770 4452
rect 15837 4450 15903 4453
rect 19149 4450 19215 4453
rect 15837 4448 19215 4450
rect 15837 4392 15842 4448
rect 15898 4392 19154 4448
rect 19210 4392 19215 4448
rect 15837 4390 19215 4392
rect 15837 4387 15903 4390
rect 19149 4387 19215 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 2405 4314 2471 4317
rect 2957 4314 3023 4317
rect 2405 4312 3023 4314
rect 2405 4256 2410 4312
rect 2466 4256 2962 4312
rect 3018 4256 3023 4312
rect 2405 4254 3023 4256
rect 2405 4251 2471 4254
rect 2957 4251 3023 4254
rect 8201 4314 8267 4317
rect 18086 4314 18092 4316
rect 8201 4312 18092 4314
rect 8201 4256 8206 4312
rect 8262 4256 18092 4312
rect 8201 4254 18092 4256
rect 8201 4251 8267 4254
rect 18086 4252 18092 4254
rect 18156 4252 18162 4316
rect 200 4178 800 4208
rect 3969 4178 4035 4181
rect 200 4176 4035 4178
rect 200 4120 3974 4176
rect 4030 4120 4035 4176
rect 200 4118 4035 4120
rect 200 4088 800 4118
rect 3969 4115 4035 4118
rect 5993 4178 6059 4181
rect 12014 4178 12020 4180
rect 5993 4176 12020 4178
rect 5993 4120 5998 4176
rect 6054 4120 12020 4176
rect 5993 4118 12020 4120
rect 5993 4115 6059 4118
rect 12014 4116 12020 4118
rect 12084 4116 12090 4180
rect 12157 4176 12223 4181
rect 12157 4120 12162 4176
rect 12218 4120 12223 4176
rect 12157 4115 12223 4120
rect 12801 4178 12867 4181
rect 16389 4178 16455 4181
rect 12801 4176 16455 4178
rect 12801 4120 12806 4176
rect 12862 4120 16394 4176
rect 16450 4120 16455 4176
rect 12801 4118 16455 4120
rect 12801 4115 12867 4118
rect 16389 4115 16455 4118
rect 17033 4178 17099 4181
rect 20621 4178 20687 4181
rect 17033 4176 20687 4178
rect 17033 4120 17038 4176
rect 17094 4120 20626 4176
rect 20682 4120 20687 4176
rect 17033 4118 20687 4120
rect 17033 4115 17099 4118
rect 20621 4115 20687 4118
rect 38193 4178 38259 4181
rect 39200 4178 39800 4208
rect 38193 4176 39800 4178
rect 38193 4120 38198 4176
rect 38254 4120 39800 4176
rect 38193 4118 39800 4120
rect 38193 4115 38259 4118
rect 6545 4042 6611 4045
rect 6862 4042 6868 4044
rect 6545 4040 6868 4042
rect 6545 3984 6550 4040
rect 6606 3984 6868 4040
rect 6545 3982 6868 3984
rect 6545 3979 6611 3982
rect 6862 3980 6868 3982
rect 6932 3980 6938 4044
rect 7281 4042 7347 4045
rect 8477 4044 8543 4045
rect 7414 4042 7420 4044
rect 7281 4040 7420 4042
rect 7281 3984 7286 4040
rect 7342 3984 7420 4040
rect 7281 3982 7420 3984
rect 7281 3979 7347 3982
rect 7414 3980 7420 3982
rect 7484 3980 7490 4044
rect 8477 4042 8524 4044
rect 8432 4040 8524 4042
rect 8432 3984 8482 4040
rect 8432 3982 8524 3984
rect 8477 3980 8524 3982
rect 8588 3980 8594 4044
rect 9029 4042 9095 4045
rect 12160 4042 12220 4115
rect 39200 4088 39800 4118
rect 9029 4040 12220 4042
rect 9029 3984 9034 4040
rect 9090 3984 12220 4040
rect 9029 3982 12220 3984
rect 12525 4042 12591 4045
rect 14089 4042 14155 4045
rect 14273 4044 14339 4045
rect 12525 4040 14155 4042
rect 12525 3984 12530 4040
rect 12586 3984 14094 4040
rect 14150 3984 14155 4040
rect 12525 3982 14155 3984
rect 8477 3979 8543 3980
rect 9029 3979 9095 3982
rect 12525 3979 12591 3982
rect 14089 3979 14155 3982
rect 14222 3980 14228 4044
rect 14292 4042 14339 4044
rect 14457 4042 14523 4045
rect 15837 4042 15903 4045
rect 14292 4040 14384 4042
rect 14334 3984 14384 4040
rect 14292 3982 14384 3984
rect 14457 4040 15903 4042
rect 14457 3984 14462 4040
rect 14518 3984 15842 4040
rect 15898 3984 15903 4040
rect 14457 3982 15903 3984
rect 14292 3980 14339 3982
rect 14273 3979 14339 3980
rect 14457 3979 14523 3982
rect 15837 3979 15903 3982
rect 17534 3980 17540 4044
rect 17604 4042 17610 4044
rect 19517 4042 19583 4045
rect 17604 4040 19583 4042
rect 17604 3984 19522 4040
rect 19578 3984 19583 4040
rect 17604 3982 19583 3984
rect 17604 3980 17610 3982
rect 19517 3979 19583 3982
rect 19885 4042 19951 4045
rect 21725 4042 21791 4045
rect 22001 4044 22067 4045
rect 21950 4042 21956 4044
rect 19885 4040 21791 4042
rect 19885 3984 19890 4040
rect 19946 3984 21730 4040
rect 21786 3984 21791 4040
rect 19885 3982 21791 3984
rect 21910 3982 21956 4042
rect 22020 4040 22067 4044
rect 22062 3984 22067 4040
rect 19885 3979 19951 3982
rect 21725 3979 21791 3982
rect 21950 3980 21956 3982
rect 22020 3980 22067 3984
rect 22001 3979 22067 3980
rect 7741 3906 7807 3909
rect 15561 3906 15627 3909
rect 7741 3904 15627 3906
rect 7741 3848 7746 3904
rect 7802 3848 15566 3904
rect 15622 3848 15627 3904
rect 7741 3846 15627 3848
rect 7741 3843 7807 3846
rect 15561 3843 15627 3846
rect 16062 3844 16068 3908
rect 16132 3906 16138 3908
rect 23933 3906 23999 3909
rect 16132 3904 23999 3906
rect 16132 3848 23938 3904
rect 23994 3848 23999 3904
rect 16132 3846 23999 3848
rect 16132 3844 16138 3846
rect 23933 3843 23999 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 7925 3770 7991 3773
rect 12525 3770 12591 3773
rect 7925 3768 12591 3770
rect 7925 3712 7930 3768
rect 7986 3712 12530 3768
rect 12586 3712 12591 3768
rect 7925 3710 12591 3712
rect 7925 3707 7991 3710
rect 12525 3707 12591 3710
rect 14089 3770 14155 3773
rect 18638 3770 18644 3772
rect 14089 3768 18644 3770
rect 14089 3712 14094 3768
rect 14150 3712 18644 3768
rect 14089 3710 18644 3712
rect 14089 3707 14155 3710
rect 18638 3708 18644 3710
rect 18708 3708 18714 3772
rect 18822 3708 18828 3772
rect 18892 3770 18898 3772
rect 21357 3770 21423 3773
rect 18892 3768 21423 3770
rect 18892 3712 21362 3768
rect 21418 3712 21423 3768
rect 18892 3710 21423 3712
rect 18892 3708 18898 3710
rect 21357 3707 21423 3710
rect 2957 3634 3023 3637
rect 2957 3632 8816 3634
rect 2957 3576 2962 3632
rect 3018 3576 8816 3632
rect 2957 3574 8816 3576
rect 2957 3571 3023 3574
rect 200 3498 800 3528
rect 3785 3498 3851 3501
rect 200 3496 3851 3498
rect 200 3440 3790 3496
rect 3846 3440 3851 3496
rect 200 3438 3851 3440
rect 8756 3498 8816 3574
rect 8886 3572 8892 3636
rect 8956 3634 8962 3636
rect 9029 3634 9095 3637
rect 8956 3632 9095 3634
rect 8956 3576 9034 3632
rect 9090 3576 9095 3632
rect 8956 3574 9095 3576
rect 8956 3572 8962 3574
rect 9029 3571 9095 3574
rect 9213 3634 9279 3637
rect 16205 3634 16271 3637
rect 9213 3632 16271 3634
rect 9213 3576 9218 3632
rect 9274 3576 16210 3632
rect 16266 3576 16271 3632
rect 9213 3574 16271 3576
rect 9213 3571 9279 3574
rect 16205 3571 16271 3574
rect 16389 3634 16455 3637
rect 20621 3634 20687 3637
rect 16389 3632 20687 3634
rect 16389 3576 16394 3632
rect 16450 3576 20626 3632
rect 20682 3576 20687 3632
rect 16389 3574 20687 3576
rect 16389 3571 16455 3574
rect 20621 3571 20687 3574
rect 9673 3498 9739 3501
rect 8756 3496 9739 3498
rect 8756 3440 9678 3496
rect 9734 3440 9739 3496
rect 8756 3438 9739 3440
rect 200 3408 800 3438
rect 3785 3435 3851 3438
rect 9673 3435 9739 3438
rect 9806 3436 9812 3500
rect 9876 3498 9882 3500
rect 10317 3498 10383 3501
rect 9876 3496 10383 3498
rect 9876 3440 10322 3496
rect 10378 3440 10383 3496
rect 9876 3438 10383 3440
rect 9876 3436 9882 3438
rect 10317 3435 10383 3438
rect 10685 3498 10751 3501
rect 20253 3498 20319 3501
rect 24025 3498 24091 3501
rect 10685 3496 20178 3498
rect 10685 3440 10690 3496
rect 10746 3440 20178 3496
rect 10685 3438 20178 3440
rect 10685 3435 10751 3438
rect 2957 3362 3023 3365
rect 18781 3362 18847 3365
rect 2957 3360 18847 3362
rect 2957 3304 2962 3360
rect 3018 3304 18786 3360
rect 18842 3304 18847 3360
rect 2957 3302 18847 3304
rect 20118 3362 20178 3438
rect 20253 3496 24091 3498
rect 20253 3440 20258 3496
rect 20314 3440 24030 3496
rect 24086 3440 24091 3496
rect 20253 3438 24091 3440
rect 20253 3435 20319 3438
rect 24025 3435 24091 3438
rect 26049 3362 26115 3365
rect 20118 3360 26115 3362
rect 20118 3304 26054 3360
rect 26110 3304 26115 3360
rect 20118 3302 26115 3304
rect 2957 3299 3023 3302
rect 18781 3299 18847 3302
rect 26049 3299 26115 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4245 3226 4311 3229
rect 8201 3226 8267 3229
rect 12985 3226 13051 3229
rect 16297 3228 16363 3229
rect 4245 3224 5642 3226
rect 4245 3168 4250 3224
rect 4306 3168 5642 3224
rect 4245 3166 5642 3168
rect 4245 3163 4311 3166
rect 3509 3090 3575 3093
rect 5349 3090 5415 3093
rect 3509 3088 5415 3090
rect 3509 3032 3514 3088
rect 3570 3032 5354 3088
rect 5410 3032 5415 3088
rect 3509 3030 5415 3032
rect 5582 3090 5642 3166
rect 8201 3224 13051 3226
rect 8201 3168 8206 3224
rect 8262 3168 12990 3224
rect 13046 3168 13051 3224
rect 8201 3166 13051 3168
rect 8201 3163 8267 3166
rect 12985 3163 13051 3166
rect 16246 3164 16252 3228
rect 16316 3226 16363 3228
rect 16573 3226 16639 3229
rect 19149 3226 19215 3229
rect 16316 3224 16408 3226
rect 16358 3168 16408 3224
rect 16316 3166 16408 3168
rect 16573 3224 19215 3226
rect 16573 3168 16578 3224
rect 16634 3168 19154 3224
rect 19210 3168 19215 3224
rect 16573 3166 19215 3168
rect 16316 3164 16363 3166
rect 16297 3163 16363 3164
rect 16573 3163 16639 3166
rect 19149 3163 19215 3166
rect 25405 3090 25471 3093
rect 5582 3088 25471 3090
rect 5582 3032 25410 3088
rect 25466 3032 25471 3088
rect 5582 3030 25471 3032
rect 3509 3027 3575 3030
rect 5349 3027 5415 3030
rect 25405 3027 25471 3030
rect 5533 2956 5599 2957
rect 5533 2954 5580 2956
rect 5488 2952 5580 2954
rect 5488 2896 5538 2952
rect 5488 2894 5580 2896
rect 5533 2892 5580 2894
rect 5644 2892 5650 2956
rect 6545 2954 6611 2957
rect 25037 2954 25103 2957
rect 6545 2952 25103 2954
rect 6545 2896 6550 2952
rect 6606 2896 25042 2952
rect 25098 2896 25103 2952
rect 6545 2894 25103 2896
rect 5533 2891 5599 2892
rect 6545 2891 6611 2894
rect 25037 2891 25103 2894
rect 200 2818 800 2848
rect 3969 2818 4035 2821
rect 200 2816 4035 2818
rect 200 2760 3974 2816
rect 4030 2760 4035 2816
rect 200 2758 4035 2760
rect 200 2728 800 2758
rect 3969 2755 4035 2758
rect 6361 2818 6427 2821
rect 16665 2818 16731 2821
rect 6361 2816 16731 2818
rect 6361 2760 6366 2816
rect 6422 2760 16670 2816
rect 16726 2760 16731 2816
rect 6361 2758 16731 2760
rect 6361 2755 6427 2758
rect 16665 2755 16731 2758
rect 18965 2818 19031 2821
rect 21817 2818 21883 2821
rect 18965 2816 21883 2818
rect 18965 2760 18970 2816
rect 19026 2760 21822 2816
rect 21878 2760 21883 2816
rect 18965 2758 21883 2760
rect 18965 2755 19031 2758
rect 21817 2755 21883 2758
rect 36905 2818 36971 2821
rect 39200 2818 39800 2848
rect 36905 2816 39800 2818
rect 36905 2760 36910 2816
rect 36966 2760 39800 2816
rect 36905 2758 39800 2760
rect 36905 2755 36971 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 39800 2758
rect 34930 2687 35246 2688
rect 5257 2682 5323 2685
rect 8334 2682 8340 2684
rect 5257 2680 8340 2682
rect 5257 2624 5262 2680
rect 5318 2624 8340 2680
rect 5257 2622 8340 2624
rect 5257 2619 5323 2622
rect 8334 2620 8340 2622
rect 8404 2620 8410 2684
rect 10869 2682 10935 2685
rect 23289 2682 23355 2685
rect 10869 2680 23355 2682
rect 10869 2624 10874 2680
rect 10930 2624 23294 2680
rect 23350 2624 23355 2680
rect 10869 2622 23355 2624
rect 10869 2619 10935 2622
rect 23289 2619 23355 2622
rect 4613 2546 4679 2549
rect 5206 2546 5212 2548
rect 4613 2544 5212 2546
rect 4613 2488 4618 2544
rect 4674 2488 5212 2544
rect 4613 2486 5212 2488
rect 4613 2483 4679 2486
rect 5206 2484 5212 2486
rect 5276 2484 5282 2548
rect 6821 2546 6887 2549
rect 19057 2546 19123 2549
rect 6821 2544 19123 2546
rect 6821 2488 6826 2544
rect 6882 2488 19062 2544
rect 19118 2488 19123 2544
rect 6821 2486 19123 2488
rect 6821 2483 6887 2486
rect 19057 2483 19123 2486
rect 19241 2546 19307 2549
rect 20294 2546 20300 2548
rect 19241 2544 20300 2546
rect 19241 2488 19246 2544
rect 19302 2488 20300 2544
rect 19241 2486 20300 2488
rect 19241 2483 19307 2486
rect 20294 2484 20300 2486
rect 20364 2484 20370 2548
rect 21766 2484 21772 2548
rect 21836 2546 21842 2548
rect 23289 2546 23355 2549
rect 21836 2544 23355 2546
rect 21836 2488 23294 2544
rect 23350 2488 23355 2544
rect 21836 2486 23355 2488
rect 21836 2484 21842 2486
rect 23289 2483 23355 2486
rect 10961 2410 11027 2413
rect 20529 2410 20595 2413
rect 10961 2408 20595 2410
rect 10961 2352 10966 2408
rect 11022 2352 20534 2408
rect 20590 2352 20595 2408
rect 10961 2350 20595 2352
rect 10961 2347 11027 2350
rect 20529 2347 20595 2350
rect 21582 2348 21588 2412
rect 21652 2410 21658 2412
rect 30373 2410 30439 2413
rect 21652 2408 30439 2410
rect 21652 2352 30378 2408
rect 30434 2352 30439 2408
rect 21652 2350 30439 2352
rect 21652 2348 21658 2350
rect 30373 2347 30439 2350
rect 6085 2274 6151 2277
rect 15469 2274 15535 2277
rect 6085 2272 15535 2274
rect 6085 2216 6090 2272
rect 6146 2216 15474 2272
rect 15530 2216 15535 2272
rect 6085 2214 15535 2216
rect 6085 2211 6151 2214
rect 15469 2211 15535 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 10225 2138 10291 2141
rect 15009 2138 15075 2141
rect 19241 2138 19307 2141
rect 10225 2136 19307 2138
rect 10225 2080 10230 2136
rect 10286 2080 15014 2136
rect 15070 2080 19246 2136
rect 19302 2080 19307 2136
rect 10225 2078 19307 2080
rect 10225 2075 10291 2078
rect 15009 2075 15075 2078
rect 19241 2075 19307 2078
rect 37181 2138 37247 2141
rect 39200 2138 39800 2168
rect 37181 2136 39800 2138
rect 37181 2080 37186 2136
rect 37242 2080 39800 2136
rect 37181 2078 39800 2080
rect 37181 2075 37247 2078
rect 39200 2048 39800 2078
rect 8385 2002 8451 2005
rect 22277 2002 22343 2005
rect 8385 2000 22343 2002
rect 8385 1944 8390 2000
rect 8446 1944 22282 2000
rect 22338 1944 22343 2000
rect 8385 1942 22343 1944
rect 8385 1939 8451 1942
rect 22277 1939 22343 1942
rect 5165 1866 5231 1869
rect 20253 1866 20319 1869
rect 5165 1864 20319 1866
rect 5165 1808 5170 1864
rect 5226 1808 20258 1864
rect 20314 1808 20319 1864
rect 5165 1806 20319 1808
rect 5165 1803 5231 1806
rect 20253 1803 20319 1806
rect 8293 1730 8359 1733
rect 17493 1730 17559 1733
rect 8293 1728 17559 1730
rect 8293 1672 8298 1728
rect 8354 1672 17498 1728
rect 17554 1672 17559 1728
rect 8293 1670 17559 1672
rect 8293 1667 8359 1670
rect 17493 1667 17559 1670
rect 200 1458 800 1488
rect 6453 1458 6519 1461
rect 200 1456 6519 1458
rect 200 1400 6458 1456
rect 6514 1400 6519 1456
rect 200 1398 6519 1400
rect 200 1368 800 1398
rect 6453 1395 6519 1398
rect 5022 1260 5028 1324
rect 5092 1322 5098 1324
rect 23381 1322 23447 1325
rect 5092 1320 23447 1322
rect 5092 1264 23386 1320
rect 23442 1264 23447 1320
rect 5092 1262 23447 1264
rect 5092 1260 5098 1262
rect 23381 1259 23447 1262
rect 200 778 800 808
rect 3509 778 3575 781
rect 200 776 3575 778
rect 200 720 3514 776
rect 3570 720 3575 776
rect 200 718 3575 720
rect 200 688 800 718
rect 3509 715 3575 718
rect 38285 778 38351 781
rect 39200 778 39800 808
rect 38285 776 39800 778
rect 38285 720 38290 776
rect 38346 720 39800 776
rect 38285 718 39800 720
rect 38285 715 38351 718
rect 39200 688 39800 718
rect 37273 98 37339 101
rect 39200 98 39800 128
rect 37273 96 39800 98
rect 37273 40 37278 96
rect 37334 40 39800 96
rect 37273 38 39800 40
rect 37273 35 37339 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 8524 36484 8588 36548
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 27292 33084 27356 33148
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 1164 30364 1228 30428
rect 2084 30424 2148 30428
rect 2084 30368 2098 30424
rect 2098 30368 2148 30424
rect 2084 30364 2148 30368
rect 4844 30364 4908 30428
rect 5396 30364 5460 30428
rect 12756 30364 12820 30428
rect 22692 30364 22756 30428
rect 21588 30228 21652 30292
rect 16252 30152 16316 30156
rect 16252 30096 16302 30152
rect 16302 30096 16316 30152
rect 16252 30092 16316 30096
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 3556 29276 3620 29340
rect 7420 29140 7484 29204
rect 1900 29004 1964 29068
rect 6500 29004 6564 29068
rect 11652 29004 11716 29068
rect 21956 28868 22020 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 5212 28596 5276 28660
rect 4660 28460 4724 28524
rect 6684 28460 6748 28524
rect 16988 28324 17052 28388
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 16252 28052 16316 28116
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 2820 27644 2884 27708
rect 7052 27704 7116 27708
rect 7052 27648 7066 27704
rect 7066 27648 7116 27704
rect 7052 27644 7116 27648
rect 9812 27644 9876 27708
rect 10732 27704 10796 27708
rect 10732 27648 10746 27704
rect 10746 27648 10796 27704
rect 10732 27644 10796 27648
rect 14964 27644 15028 27708
rect 14780 27508 14844 27572
rect 8340 27432 8404 27436
rect 8340 27376 8390 27432
rect 8390 27376 8404 27432
rect 8340 27372 8404 27376
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 3740 27100 3804 27164
rect 5028 27024 5092 27028
rect 5028 26968 5042 27024
rect 5042 26968 5092 27024
rect 5028 26964 5092 26968
rect 5580 26828 5644 26892
rect 6868 26692 6932 26756
rect 16068 26828 16132 26892
rect 8708 26692 8772 26756
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 9260 26692 9324 26756
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 13676 26556 13740 26620
rect 10916 26480 10980 26484
rect 10916 26424 10966 26480
rect 10966 26424 10980 26480
rect 10916 26420 10980 26424
rect 3372 26284 3436 26348
rect 6132 26284 6196 26348
rect 7604 26284 7668 26348
rect 12572 26284 12636 26348
rect 17724 26344 17788 26348
rect 17724 26288 17738 26344
rect 17738 26288 17788 26344
rect 17724 26284 17788 26288
rect 20116 26284 20180 26348
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 23060 25876 23124 25940
rect 7236 25800 7300 25804
rect 7236 25744 7286 25800
rect 7286 25744 7300 25800
rect 7236 25740 7300 25744
rect 15516 25664 15580 25668
rect 15516 25608 15530 25664
rect 15530 25608 15580 25664
rect 15516 25604 15580 25608
rect 22876 25604 22940 25668
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 5212 24924 5276 24988
rect 5948 24984 6012 24988
rect 5948 24928 5962 24984
rect 5962 24928 6012 24984
rect 5948 24924 6012 24928
rect 13860 24924 13924 24988
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 5580 24652 5644 24716
rect 9996 24652 10060 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 20116 24380 20180 24444
rect 11284 24244 11348 24308
rect 12756 24108 12820 24172
rect 16804 23972 16868 24036
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 5580 23428 5644 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 8892 23488 8956 23492
rect 8892 23432 8906 23488
rect 8906 23432 8956 23488
rect 8892 23428 8956 23432
rect 10548 23428 10612 23492
rect 21772 23428 21836 23492
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 12940 23292 13004 23356
rect 5028 23216 5092 23220
rect 5028 23160 5078 23216
rect 5078 23160 5092 23216
rect 5028 23156 5092 23160
rect 5212 23156 5276 23220
rect 5028 23020 5092 23084
rect 9812 23080 9876 23084
rect 9812 23024 9826 23080
rect 9826 23024 9876 23080
rect 9812 23020 9876 23024
rect 8340 22884 8404 22948
rect 7420 22748 7484 22812
rect 16988 22748 17052 22812
rect 24716 22884 24780 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 12940 22340 13004 22404
rect 13124 22340 13188 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 5764 22204 5828 22268
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 9444 22068 9508 22132
rect 12388 22068 12452 22132
rect 5764 21932 5828 21996
rect 12756 22068 12820 22132
rect 13492 21932 13556 21996
rect 22692 22068 22756 22132
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 1900 21584 1964 21588
rect 1900 21528 1950 21584
rect 1950 21528 1964 21584
rect 1900 21524 1964 21528
rect 9628 21524 9692 21588
rect 26924 21992 26988 21996
rect 26924 21936 26938 21992
rect 26938 21936 26988 21992
rect 26924 21932 26988 21936
rect 14596 21388 14660 21452
rect 18828 21388 18892 21452
rect 3740 21252 3804 21316
rect 5396 21252 5460 21316
rect 12756 21252 12820 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 5028 21116 5092 21180
rect 19196 21116 19260 21180
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 10180 20980 10244 21044
rect 19196 20980 19260 21044
rect 9260 20844 9324 20908
rect 9812 20844 9876 20908
rect 6684 20708 6748 20772
rect 15516 20768 15580 20772
rect 15516 20712 15566 20768
rect 15566 20712 15580 20768
rect 15516 20708 15580 20712
rect 20116 20768 20180 20772
rect 20116 20712 20166 20768
rect 20166 20712 20180 20768
rect 20116 20708 20180 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 12204 20572 12268 20636
rect 12388 20572 12452 20636
rect 20484 20436 20548 20500
rect 6868 20300 6932 20364
rect 11836 20300 11900 20364
rect 17356 20300 17420 20364
rect 6500 20224 6564 20228
rect 6500 20168 6514 20224
rect 6514 20168 6564 20224
rect 6500 20164 6564 20168
rect 6868 20164 6932 20228
rect 27108 20164 27172 20228
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 20668 20028 20732 20092
rect 4844 19816 4908 19820
rect 4844 19760 4894 19816
rect 4894 19760 4908 19816
rect 4844 19756 4908 19760
rect 7788 19756 7852 19820
rect 10180 19816 10244 19820
rect 10180 19760 10230 19816
rect 10230 19760 10244 19816
rect 10180 19756 10244 19760
rect 12388 19756 12452 19820
rect 18828 19892 18892 19956
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 20116 19816 20180 19820
rect 20116 19760 20166 19816
rect 20166 19760 20180 19816
rect 20116 19756 20180 19760
rect 20668 19756 20732 19820
rect 20116 19620 20180 19684
rect 2820 19408 2884 19412
rect 2820 19352 2870 19408
rect 2870 19352 2884 19408
rect 2820 19348 2884 19352
rect 4660 19348 4724 19412
rect 9996 19212 10060 19276
rect 11652 19076 11716 19140
rect 20116 19348 20180 19412
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 9260 18940 9324 19004
rect 10364 18940 10428 19004
rect 10916 18940 10980 19004
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 10916 18804 10980 18868
rect 17724 18668 17788 18732
rect 12020 18532 12084 18596
rect 14780 18396 14844 18460
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 7420 18260 7484 18324
rect 21036 18260 21100 18324
rect 22140 18260 22204 18324
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 13860 17988 13924 18052
rect 16804 17988 16868 18052
rect 17172 17988 17236 18052
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 10548 17852 10612 17916
rect 16068 17852 16132 17916
rect 8892 17580 8956 17644
rect 16988 17716 17052 17780
rect 20116 17716 20180 17780
rect 21220 17852 21284 17916
rect 26372 17716 26436 17780
rect 7604 17444 7668 17508
rect 17540 17444 17604 17508
rect 21220 17444 21284 17508
rect 22140 17444 22204 17508
rect 22324 17444 22388 17508
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 13860 17308 13924 17372
rect 11284 17172 11348 17236
rect 18276 17232 18340 17236
rect 18276 17176 18326 17232
rect 18326 17176 18340 17232
rect 18276 17172 18340 17176
rect 18828 17172 18892 17236
rect 17356 17036 17420 17100
rect 19012 17036 19076 17100
rect 21220 17036 21284 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 14964 16764 15028 16828
rect 7236 16628 7300 16692
rect 8708 16628 8772 16692
rect 9260 16628 9324 16692
rect 20484 16628 20548 16692
rect 20852 16628 20916 16692
rect 6868 16356 6932 16420
rect 12388 16356 12452 16420
rect 9076 16220 9140 16284
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 20852 16084 20916 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 3556 15676 3620 15740
rect 13860 15812 13924 15876
rect 14596 15812 14660 15876
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 17908 15676 17972 15740
rect 18092 15736 18156 15740
rect 18092 15680 18142 15736
rect 18142 15680 18156 15736
rect 18092 15676 18156 15680
rect 24900 15736 24964 15740
rect 24900 15680 24914 15736
rect 24914 15680 24964 15736
rect 24900 15676 24964 15680
rect 14780 15404 14844 15468
rect 17356 15404 17420 15468
rect 17908 15404 17972 15468
rect 7788 15192 7852 15196
rect 7788 15136 7838 15192
rect 7838 15136 7852 15192
rect 7788 15132 7852 15136
rect 9444 15132 9508 15196
rect 12020 15268 12084 15332
rect 18460 15268 18524 15332
rect 20852 15328 20916 15332
rect 20852 15272 20902 15328
rect 20902 15272 20916 15328
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 12204 15132 12268 15196
rect 18828 15132 18892 15196
rect 20116 15132 20180 15196
rect 20852 15268 20916 15272
rect 3924 14996 3988 15060
rect 10732 14860 10796 14924
rect 26188 14996 26252 15060
rect 27292 15056 27356 15060
rect 27292 15000 27342 15056
rect 27342 15000 27356 15056
rect 27292 14996 27356 15000
rect 19196 14724 19260 14788
rect 21036 14724 21100 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 18460 14588 18524 14652
rect 22508 14724 22572 14788
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 14780 14452 14844 14516
rect 15884 14452 15948 14516
rect 21036 14512 21100 14516
rect 21036 14456 21086 14512
rect 21086 14456 21100 14512
rect 21036 14452 21100 14456
rect 6132 14044 6196 14108
rect 14964 14044 15028 14108
rect 18828 14180 18892 14244
rect 19196 14180 19260 14244
rect 19380 14240 19444 14244
rect 19380 14184 19394 14240
rect 19394 14184 19444 14240
rect 19380 14180 19444 14184
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 18460 14044 18524 14108
rect 18828 14044 18892 14108
rect 26372 14240 26436 14244
rect 26372 14184 26422 14240
rect 26422 14184 26436 14240
rect 26372 14180 26436 14184
rect 5948 13908 6012 13972
rect 16620 13908 16684 13972
rect 26004 13908 26068 13972
rect 27108 13772 27172 13836
rect 27660 13832 27724 13836
rect 27660 13776 27674 13832
rect 27674 13776 27724 13832
rect 27660 13772 27724 13776
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 10364 13500 10428 13564
rect 14780 13500 14844 13564
rect 21036 13696 21100 13700
rect 21036 13640 21086 13696
rect 21086 13640 21100 13696
rect 21036 13636 21100 13640
rect 21404 13636 21468 13700
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 14228 13364 14292 13428
rect 13124 13092 13188 13156
rect 19012 13152 19076 13156
rect 19012 13096 19062 13152
rect 19062 13096 19076 13152
rect 19012 13092 19076 13096
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 15700 12956 15764 13020
rect 3924 12820 3988 12884
rect 5396 12880 5460 12884
rect 5396 12824 5446 12880
rect 5446 12824 5460 12880
rect 5028 12684 5092 12748
rect 5396 12820 5460 12824
rect 19012 12820 19076 12884
rect 20116 12956 20180 13020
rect 21036 12820 21100 12884
rect 16804 12684 16868 12748
rect 18092 12684 18156 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 9628 12412 9692 12476
rect 11468 12412 11532 12476
rect 16620 12412 16684 12476
rect 8524 12336 8588 12340
rect 8524 12280 8574 12336
rect 8574 12280 8588 12336
rect 8524 12276 8588 12280
rect 11100 12276 11164 12340
rect 20116 12276 20180 12340
rect 20668 12064 20732 12068
rect 20668 12008 20682 12064
rect 20682 12008 20732 12064
rect 20668 12004 20732 12008
rect 22324 12004 22388 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 8340 11656 8404 11660
rect 8340 11600 8390 11656
rect 8390 11600 8404 11656
rect 8340 11596 8404 11600
rect 11468 11596 11532 11660
rect 12388 11596 12452 11660
rect 17724 11596 17788 11660
rect 18276 11656 18340 11660
rect 18276 11600 18290 11656
rect 18290 11600 18340 11656
rect 18276 11596 18340 11600
rect 19380 11868 19444 11932
rect 20116 11868 20180 11932
rect 22876 11868 22940 11932
rect 21588 11732 21652 11796
rect 5396 11520 5460 11524
rect 5396 11464 5446 11520
rect 5446 11464 5460 11520
rect 5396 11460 5460 11464
rect 19978 11460 20042 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 13124 11324 13188 11388
rect 17540 11324 17604 11388
rect 17724 11324 17788 11388
rect 21404 11460 21468 11524
rect 22324 11460 22388 11524
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 20484 11324 20548 11388
rect 9260 10916 9324 10980
rect 10732 10780 10796 10844
rect 14412 10976 14476 10980
rect 18644 11052 18708 11116
rect 14412 10920 14462 10976
rect 14462 10920 14476 10976
rect 14412 10916 14476 10920
rect 17908 10916 17972 10980
rect 18644 10916 18708 10980
rect 19196 10976 19260 10980
rect 19196 10920 19246 10976
rect 19246 10920 19260 10976
rect 19196 10916 19260 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 12940 10780 13004 10844
rect 13492 10780 13556 10844
rect 19380 10780 19444 10844
rect 20116 10780 20180 10844
rect 14228 10644 14292 10708
rect 17724 10508 17788 10572
rect 17908 10508 17972 10572
rect 14964 10372 15028 10436
rect 16436 10372 16500 10436
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 11100 10236 11164 10300
rect 3372 10100 3436 10164
rect 13860 10100 13924 10164
rect 17540 10100 17604 10164
rect 20116 10100 20180 10164
rect 20852 10100 20916 10164
rect 12940 9964 13004 10028
rect 16620 9964 16684 10028
rect 10916 9828 10980 9892
rect 11468 9828 11532 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 14412 9692 14476 9756
rect 15516 9692 15580 9756
rect 1164 9556 1228 9620
rect 18644 9692 18708 9756
rect 19380 9692 19444 9756
rect 22140 9692 22204 9756
rect 9076 9420 9140 9484
rect 20484 9420 20548 9484
rect 16068 9284 16132 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 12020 9012 12084 9076
rect 12204 9012 12268 9076
rect 17540 9012 17604 9076
rect 18092 9012 18156 9076
rect 24900 9012 24964 9076
rect 16436 8740 16500 8804
rect 11468 8604 11532 8668
rect 19196 8740 19260 8804
rect 20484 8740 20548 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 17356 8604 17420 8668
rect 9444 8332 9508 8396
rect 14044 8332 14108 8396
rect 14596 8332 14660 8396
rect 15884 8332 15948 8396
rect 13676 8256 13740 8260
rect 13676 8200 13690 8256
rect 13690 8200 13740 8256
rect 13676 8196 13740 8200
rect 19012 8196 19076 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 7052 8060 7116 8124
rect 12204 7924 12268 7988
rect 16804 7924 16868 7988
rect 17356 8120 17420 8124
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 17356 8064 17370 8120
rect 17370 8064 17420 8120
rect 17356 8060 17420 8064
rect 20668 8060 20732 8124
rect 9812 7788 9876 7852
rect 11284 7788 11348 7852
rect 19380 7788 19444 7852
rect 21404 7788 21468 7852
rect 16804 7652 16868 7716
rect 17172 7652 17236 7716
rect 17724 7652 17788 7716
rect 8892 7516 8956 7580
rect 16620 7516 16684 7580
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 19196 7516 19260 7580
rect 20300 7516 20364 7580
rect 22140 7244 22204 7308
rect 22508 7108 22572 7172
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 9812 6972 9876 7036
rect 10364 7032 10428 7036
rect 10364 6976 10414 7032
rect 10414 6976 10428 7032
rect 10364 6972 10428 6976
rect 10916 7032 10980 7036
rect 10916 6976 10930 7032
rect 10930 6976 10980 7032
rect 10916 6972 10980 6976
rect 11652 6972 11716 7036
rect 18460 6972 18524 7036
rect 18644 7032 18708 7036
rect 18644 6976 18658 7032
rect 18658 6976 18708 7032
rect 18644 6972 18708 6976
rect 19196 6972 19260 7036
rect 20300 6972 20364 7036
rect 5580 6428 5644 6492
rect 15700 6836 15764 6900
rect 23060 6836 23124 6900
rect 24716 6896 24780 6900
rect 24716 6840 24730 6896
rect 24730 6840 24780 6896
rect 24716 6836 24780 6840
rect 12204 6700 12268 6764
rect 18276 6700 18340 6764
rect 18644 6700 18708 6764
rect 20852 6700 20916 6764
rect 22324 6700 22388 6764
rect 12388 6564 12452 6628
rect 17724 6564 17788 6628
rect 20116 6564 20180 6628
rect 21220 6564 21284 6628
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 19012 6428 19076 6492
rect 9996 6292 10060 6356
rect 10364 6292 10428 6356
rect 17908 6292 17972 6356
rect 21036 6428 21100 6492
rect 10364 6156 10428 6220
rect 10548 6156 10612 6220
rect 15516 6020 15580 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12204 5884 12268 5948
rect 12388 5884 12452 5948
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 16988 5944 17052 5948
rect 16988 5888 17038 5944
rect 17038 5888 17052 5944
rect 16988 5884 17052 5888
rect 10180 5476 10244 5540
rect 10548 5476 10612 5540
rect 12204 5612 12268 5676
rect 12756 5612 12820 5676
rect 17724 5612 17788 5676
rect 18092 5612 18156 5676
rect 8524 5400 8588 5404
rect 8524 5344 8538 5400
rect 8538 5344 8588 5400
rect 8524 5340 8588 5344
rect 10364 5340 10428 5404
rect 13860 5476 13924 5540
rect 14044 5536 14108 5540
rect 14044 5480 14058 5536
rect 14058 5480 14108 5536
rect 14044 5476 14108 5480
rect 27660 5612 27724 5676
rect 26924 5476 26988 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 18828 5340 18892 5404
rect 7052 4932 7116 4996
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 10180 4932 10244 4996
rect 18276 5068 18340 5132
rect 12020 4932 12084 4996
rect 9260 4796 9324 4860
rect 9996 4796 10060 4860
rect 13124 4796 13188 4860
rect 2084 4660 2148 4724
rect 12388 4720 12452 4724
rect 12388 4664 12402 4720
rect 12402 4664 12452 4720
rect 12388 4660 12452 4664
rect 12572 4660 12636 4724
rect 14780 4796 14844 4860
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 13492 4660 13556 4724
rect 15700 4660 15764 4724
rect 17356 4660 17420 4724
rect 15700 4388 15764 4452
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 18092 4252 18156 4316
rect 12020 4116 12084 4180
rect 6868 3980 6932 4044
rect 7420 3980 7484 4044
rect 8524 4040 8588 4044
rect 8524 3984 8538 4040
rect 8538 3984 8588 4040
rect 8524 3980 8588 3984
rect 14228 4040 14292 4044
rect 14228 3984 14278 4040
rect 14278 3984 14292 4040
rect 14228 3980 14292 3984
rect 17540 3980 17604 4044
rect 21956 4040 22020 4044
rect 21956 3984 22006 4040
rect 22006 3984 22020 4040
rect 21956 3980 22020 3984
rect 16068 3844 16132 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 18644 3708 18708 3772
rect 18828 3708 18892 3772
rect 8892 3572 8956 3636
rect 9812 3436 9876 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 16252 3224 16316 3228
rect 16252 3168 16302 3224
rect 16302 3168 16316 3224
rect 16252 3164 16316 3168
rect 5580 2952 5644 2956
rect 5580 2896 5594 2952
rect 5594 2896 5644 2952
rect 5580 2892 5644 2896
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 8340 2620 8404 2684
rect 5212 2484 5276 2548
rect 20300 2484 20364 2548
rect 21772 2484 21836 2548
rect 21588 2348 21652 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 5028 1260 5092 1324
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 8523 36548 8589 36549
rect 8523 36484 8524 36548
rect 8588 36484 8589 36548
rect 8523 36483 8589 36484
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 1163 30428 1229 30429
rect 1163 30364 1164 30428
rect 1228 30364 1229 30428
rect 1163 30363 1229 30364
rect 2083 30428 2149 30429
rect 2083 30364 2084 30428
rect 2148 30364 2149 30428
rect 2083 30363 2149 30364
rect 1166 9621 1226 30363
rect 1899 29068 1965 29069
rect 1899 29004 1900 29068
rect 1964 29004 1965 29068
rect 1899 29003 1965 29004
rect 1902 21589 1962 29003
rect 1899 21588 1965 21589
rect 1899 21524 1900 21588
rect 1964 21524 1965 21588
rect 1899 21523 1965 21524
rect 1163 9620 1229 9621
rect 1163 9556 1164 9620
rect 1228 9556 1229 9620
rect 1163 9555 1229 9556
rect 2086 4725 2146 30363
rect 4208 29952 4528 30976
rect 4843 30428 4909 30429
rect 4843 30364 4844 30428
rect 4908 30364 4909 30428
rect 4843 30363 4909 30364
rect 5395 30428 5461 30429
rect 5395 30364 5396 30428
rect 5460 30364 5461 30428
rect 5395 30363 5461 30364
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 3555 29340 3621 29341
rect 3555 29276 3556 29340
rect 3620 29276 3621 29340
rect 3555 29275 3621 29276
rect 2819 27708 2885 27709
rect 2819 27644 2820 27708
rect 2884 27644 2885 27708
rect 2819 27643 2885 27644
rect 2822 19413 2882 27643
rect 3371 26348 3437 26349
rect 3371 26284 3372 26348
rect 3436 26284 3437 26348
rect 3371 26283 3437 26284
rect 2819 19412 2885 19413
rect 2819 19348 2820 19412
rect 2884 19348 2885 19412
rect 2819 19347 2885 19348
rect 3374 10165 3434 26283
rect 3558 15741 3618 29275
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4659 28524 4725 28525
rect 4659 28460 4660 28524
rect 4724 28460 4725 28524
rect 4659 28459 4725 28460
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 3739 27164 3805 27165
rect 3739 27100 3740 27164
rect 3804 27100 3805 27164
rect 3739 27099 3805 27100
rect 3742 21317 3802 27099
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 3739 21316 3805 21317
rect 3739 21252 3740 21316
rect 3804 21252 3805 21316
rect 3739 21251 3805 21252
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4662 19413 4722 28459
rect 4846 19821 4906 30363
rect 5211 28660 5277 28661
rect 5211 28596 5212 28660
rect 5276 28596 5277 28660
rect 5211 28595 5277 28596
rect 5027 27028 5093 27029
rect 5027 26964 5028 27028
rect 5092 26964 5093 27028
rect 5027 26963 5093 26964
rect 5030 23221 5090 26963
rect 5214 24989 5274 28595
rect 5211 24988 5277 24989
rect 5211 24924 5212 24988
rect 5276 24924 5277 24988
rect 5211 24923 5277 24924
rect 5027 23220 5093 23221
rect 5027 23156 5028 23220
rect 5092 23156 5093 23220
rect 5027 23155 5093 23156
rect 5211 23220 5277 23221
rect 5211 23156 5212 23220
rect 5276 23156 5277 23220
rect 5211 23155 5277 23156
rect 5027 23084 5093 23085
rect 5027 23020 5028 23084
rect 5092 23020 5093 23084
rect 5027 23019 5093 23020
rect 5030 21181 5090 23019
rect 5027 21180 5093 21181
rect 5027 21116 5028 21180
rect 5092 21116 5093 21180
rect 5027 21115 5093 21116
rect 4843 19820 4909 19821
rect 4843 19756 4844 19820
rect 4908 19756 4909 19820
rect 4843 19755 4909 19756
rect 4659 19412 4725 19413
rect 4659 19348 4660 19412
rect 4724 19348 4725 19412
rect 4659 19347 4725 19348
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 3555 15740 3621 15741
rect 3555 15676 3556 15740
rect 3620 15676 3621 15740
rect 3555 15675 3621 15676
rect 3923 15060 3989 15061
rect 3923 14996 3924 15060
rect 3988 14996 3989 15060
rect 3923 14995 3989 14996
rect 3926 12885 3986 14995
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 4208 12544 4528 13568
rect 5027 12748 5093 12749
rect 5027 12684 5028 12748
rect 5092 12684 5093 12748
rect 5027 12683 5093 12684
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 3371 10164 3437 10165
rect 3371 10100 3372 10164
rect 3436 10100 3437 10164
rect 3371 10099 3437 10100
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 2083 4724 2149 4725
rect 2083 4660 2084 4724
rect 2148 4660 2149 4724
rect 2083 4659 2149 4660
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 5030 1325 5090 12683
rect 5214 2549 5274 23155
rect 5398 21317 5458 30363
rect 7419 29204 7485 29205
rect 7419 29140 7420 29204
rect 7484 29140 7485 29204
rect 7419 29139 7485 29140
rect 6499 29068 6565 29069
rect 6499 29004 6500 29068
rect 6564 29004 6565 29068
rect 6499 29003 6565 29004
rect 5579 26892 5645 26893
rect 5579 26828 5580 26892
rect 5644 26828 5645 26892
rect 5579 26827 5645 26828
rect 5582 24717 5642 26827
rect 6131 26348 6197 26349
rect 6131 26284 6132 26348
rect 6196 26284 6197 26348
rect 6131 26283 6197 26284
rect 5947 24988 6013 24989
rect 5947 24924 5948 24988
rect 6012 24924 6013 24988
rect 5947 24923 6013 24924
rect 5579 24716 5645 24717
rect 5579 24652 5580 24716
rect 5644 24652 5645 24716
rect 5579 24651 5645 24652
rect 5582 23493 5642 24651
rect 5579 23492 5645 23493
rect 5579 23428 5580 23492
rect 5644 23428 5645 23492
rect 5579 23427 5645 23428
rect 5763 22268 5829 22269
rect 5763 22204 5764 22268
rect 5828 22204 5829 22268
rect 5763 22203 5829 22204
rect 5766 21997 5826 22203
rect 5763 21996 5829 21997
rect 5763 21932 5764 21996
rect 5828 21932 5829 21996
rect 5763 21931 5829 21932
rect 5395 21316 5461 21317
rect 5395 21252 5396 21316
rect 5460 21252 5461 21316
rect 5395 21251 5461 21252
rect 5950 13973 6010 24923
rect 6134 14109 6194 26283
rect 6502 20229 6562 29003
rect 6683 28524 6749 28525
rect 6683 28460 6684 28524
rect 6748 28460 6749 28524
rect 6683 28459 6749 28460
rect 6686 20773 6746 28459
rect 7051 27708 7117 27709
rect 7051 27644 7052 27708
rect 7116 27644 7117 27708
rect 7051 27643 7117 27644
rect 6867 26756 6933 26757
rect 6867 26692 6868 26756
rect 6932 26692 6933 26756
rect 6867 26691 6933 26692
rect 6683 20772 6749 20773
rect 6683 20708 6684 20772
rect 6748 20708 6749 20772
rect 6683 20707 6749 20708
rect 6870 20365 6930 26691
rect 6867 20364 6933 20365
rect 6867 20300 6868 20364
rect 6932 20300 6933 20364
rect 6867 20299 6933 20300
rect 6499 20228 6565 20229
rect 6499 20164 6500 20228
rect 6564 20164 6565 20228
rect 6499 20163 6565 20164
rect 6867 20228 6933 20229
rect 6867 20164 6868 20228
rect 6932 20164 6933 20228
rect 6867 20163 6933 20164
rect 6870 16421 6930 20163
rect 6867 16420 6933 16421
rect 6867 16356 6868 16420
rect 6932 16356 6933 16420
rect 6867 16355 6933 16356
rect 6131 14108 6197 14109
rect 6131 14044 6132 14108
rect 6196 14044 6197 14108
rect 6131 14043 6197 14044
rect 5947 13972 6013 13973
rect 5947 13908 5948 13972
rect 6012 13908 6013 13972
rect 5947 13907 6013 13908
rect 5395 12884 5461 12885
rect 5395 12820 5396 12884
rect 5460 12820 5461 12884
rect 5395 12819 5461 12820
rect 5398 11525 5458 12819
rect 7054 12450 7114 27643
rect 7235 25804 7301 25805
rect 7235 25740 7236 25804
rect 7300 25740 7301 25804
rect 7235 25739 7301 25740
rect 7238 16693 7298 25739
rect 7422 22813 7482 29139
rect 8339 27436 8405 27437
rect 8339 27372 8340 27436
rect 8404 27372 8405 27436
rect 8339 27371 8405 27372
rect 7603 26348 7669 26349
rect 7603 26284 7604 26348
rect 7668 26284 7669 26348
rect 7603 26283 7669 26284
rect 7419 22812 7485 22813
rect 7419 22748 7420 22812
rect 7484 22748 7485 22812
rect 7419 22747 7485 22748
rect 7419 18324 7485 18325
rect 7419 18260 7420 18324
rect 7484 18260 7485 18324
rect 7419 18259 7485 18260
rect 7235 16692 7301 16693
rect 7235 16628 7236 16692
rect 7300 16628 7301 16692
rect 7235 16627 7301 16628
rect 6870 12390 7114 12450
rect 5395 11524 5461 11525
rect 5395 11460 5396 11524
rect 5460 11460 5461 11524
rect 5395 11459 5461 11460
rect 5579 6492 5645 6493
rect 5579 6428 5580 6492
rect 5644 6428 5645 6492
rect 5579 6427 5645 6428
rect 5582 2957 5642 6427
rect 6870 4045 6930 12390
rect 7051 8124 7117 8125
rect 7051 8060 7052 8124
rect 7116 8060 7117 8124
rect 7051 8059 7117 8060
rect 7054 4997 7114 8059
rect 7051 4996 7117 4997
rect 7051 4932 7052 4996
rect 7116 4932 7117 4996
rect 7051 4931 7117 4932
rect 7422 4045 7482 18259
rect 7606 17509 7666 26283
rect 8342 22949 8402 27371
rect 8339 22948 8405 22949
rect 8339 22884 8340 22948
rect 8404 22884 8405 22948
rect 8339 22883 8405 22884
rect 7787 19820 7853 19821
rect 7787 19756 7788 19820
rect 7852 19756 7853 19820
rect 7787 19755 7853 19756
rect 7603 17508 7669 17509
rect 7603 17444 7604 17508
rect 7668 17444 7669 17508
rect 7603 17443 7669 17444
rect 7790 15197 7850 19755
rect 7787 15196 7853 15197
rect 7787 15132 7788 15196
rect 7852 15132 7853 15196
rect 7787 15131 7853 15132
rect 8526 12341 8586 36483
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 27291 33148 27357 33149
rect 27291 33084 27292 33148
rect 27356 33084 27357 33148
rect 27291 33083 27357 33084
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 12755 30428 12821 30429
rect 12755 30364 12756 30428
rect 12820 30364 12821 30428
rect 12755 30363 12821 30364
rect 11651 29068 11717 29069
rect 11651 29004 11652 29068
rect 11716 29004 11717 29068
rect 11651 29003 11717 29004
rect 9811 27708 9877 27709
rect 9811 27644 9812 27708
rect 9876 27644 9877 27708
rect 9811 27643 9877 27644
rect 10731 27708 10797 27709
rect 10731 27644 10732 27708
rect 10796 27644 10797 27708
rect 10731 27643 10797 27644
rect 8707 26756 8773 26757
rect 8707 26692 8708 26756
rect 8772 26692 8773 26756
rect 8707 26691 8773 26692
rect 9259 26756 9325 26757
rect 9259 26692 9260 26756
rect 9324 26692 9325 26756
rect 9259 26691 9325 26692
rect 8710 16693 8770 26691
rect 8891 23492 8957 23493
rect 8891 23428 8892 23492
rect 8956 23428 8957 23492
rect 8891 23427 8957 23428
rect 8894 17645 8954 23427
rect 9262 20909 9322 26691
rect 9814 23085 9874 27643
rect 9995 24716 10061 24717
rect 9995 24652 9996 24716
rect 10060 24652 10061 24716
rect 9995 24651 10061 24652
rect 9811 23084 9877 23085
rect 9811 23020 9812 23084
rect 9876 23020 9877 23084
rect 9811 23019 9877 23020
rect 9443 22132 9509 22133
rect 9443 22068 9444 22132
rect 9508 22068 9509 22132
rect 9443 22067 9509 22068
rect 9259 20908 9325 20909
rect 9259 20844 9260 20908
rect 9324 20844 9325 20908
rect 9259 20843 9325 20844
rect 9259 19004 9325 19005
rect 9259 18940 9260 19004
rect 9324 18940 9325 19004
rect 9259 18939 9325 18940
rect 8891 17644 8957 17645
rect 8891 17580 8892 17644
rect 8956 17580 8957 17644
rect 8891 17579 8957 17580
rect 9262 16693 9322 18939
rect 8707 16692 8773 16693
rect 8707 16628 8708 16692
rect 8772 16628 8773 16692
rect 8707 16627 8773 16628
rect 9259 16692 9325 16693
rect 9259 16628 9260 16692
rect 9324 16628 9325 16692
rect 9259 16627 9325 16628
rect 9075 16284 9141 16285
rect 9075 16220 9076 16284
rect 9140 16220 9141 16284
rect 9075 16219 9141 16220
rect 8523 12340 8589 12341
rect 8523 12276 8524 12340
rect 8588 12276 8589 12340
rect 8523 12275 8589 12276
rect 8339 11660 8405 11661
rect 8339 11596 8340 11660
rect 8404 11596 8405 11660
rect 8339 11595 8405 11596
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 7419 4044 7485 4045
rect 7419 3980 7420 4044
rect 7484 3980 7485 4044
rect 7419 3979 7485 3980
rect 5579 2956 5645 2957
rect 5579 2892 5580 2956
rect 5644 2892 5645 2956
rect 5579 2891 5645 2892
rect 8342 2685 8402 11595
rect 9078 9485 9138 16219
rect 9446 15197 9506 22067
rect 9627 21588 9693 21589
rect 9627 21524 9628 21588
rect 9692 21524 9693 21588
rect 9627 21523 9693 21524
rect 9443 15196 9509 15197
rect 9443 15132 9444 15196
rect 9508 15132 9509 15196
rect 9443 15131 9509 15132
rect 9630 12477 9690 21523
rect 9811 20908 9877 20909
rect 9811 20844 9812 20908
rect 9876 20844 9877 20908
rect 9811 20843 9877 20844
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 9259 10980 9325 10981
rect 9259 10916 9260 10980
rect 9324 10916 9325 10980
rect 9259 10915 9325 10916
rect 9075 9484 9141 9485
rect 9075 9420 9076 9484
rect 9140 9420 9141 9484
rect 9075 9419 9141 9420
rect 8891 7580 8957 7581
rect 8891 7516 8892 7580
rect 8956 7516 8957 7580
rect 8891 7515 8957 7516
rect 8523 5404 8589 5405
rect 8523 5340 8524 5404
rect 8588 5340 8589 5404
rect 8523 5339 8589 5340
rect 8526 4045 8586 5339
rect 8523 4044 8589 4045
rect 8523 3980 8524 4044
rect 8588 3980 8589 4044
rect 8523 3979 8589 3980
rect 8894 3637 8954 7515
rect 9262 4861 9322 10915
rect 9443 8396 9509 8397
rect 9443 8332 9444 8396
rect 9508 8394 9509 8396
rect 9508 8334 9690 8394
rect 9508 8332 9509 8334
rect 9443 8331 9509 8332
rect 9630 7170 9690 8334
rect 9814 7853 9874 20843
rect 9998 19277 10058 24651
rect 10547 23492 10613 23493
rect 10547 23428 10548 23492
rect 10612 23428 10613 23492
rect 10547 23427 10613 23428
rect 10179 21044 10245 21045
rect 10179 20980 10180 21044
rect 10244 20980 10245 21044
rect 10179 20979 10245 20980
rect 10182 19821 10242 20979
rect 10179 19820 10245 19821
rect 10179 19756 10180 19820
rect 10244 19756 10245 19820
rect 10179 19755 10245 19756
rect 9995 19276 10061 19277
rect 9995 19212 9996 19276
rect 10060 19212 10061 19276
rect 9995 19211 10061 19212
rect 10363 19004 10429 19005
rect 10363 18940 10364 19004
rect 10428 18940 10429 19004
rect 10363 18939 10429 18940
rect 10366 13565 10426 18939
rect 10550 17917 10610 23427
rect 10547 17916 10613 17917
rect 10547 17852 10548 17916
rect 10612 17852 10613 17916
rect 10547 17851 10613 17852
rect 10734 14925 10794 27643
rect 10915 26484 10981 26485
rect 10915 26420 10916 26484
rect 10980 26420 10981 26484
rect 10915 26419 10981 26420
rect 10918 19005 10978 26419
rect 11283 24308 11349 24309
rect 11283 24244 11284 24308
rect 11348 24244 11349 24308
rect 11283 24243 11349 24244
rect 10915 19004 10981 19005
rect 10915 18940 10916 19004
rect 10980 18940 10981 19004
rect 10915 18939 10981 18940
rect 10915 18868 10981 18869
rect 10915 18804 10916 18868
rect 10980 18804 10981 18868
rect 10915 18803 10981 18804
rect 10731 14924 10797 14925
rect 10731 14860 10732 14924
rect 10796 14860 10797 14924
rect 10731 14859 10797 14860
rect 10363 13564 10429 13565
rect 10363 13500 10364 13564
rect 10428 13500 10429 13564
rect 10363 13499 10429 13500
rect 10731 10844 10797 10845
rect 10731 10780 10732 10844
rect 10796 10780 10797 10844
rect 10731 10779 10797 10780
rect 9811 7852 9877 7853
rect 9811 7788 9812 7852
rect 9876 7788 9877 7852
rect 9811 7787 9877 7788
rect 9630 7110 10610 7170
rect 9811 7036 9877 7037
rect 9811 6972 9812 7036
rect 9876 6972 9877 7036
rect 9811 6971 9877 6972
rect 10363 7036 10429 7037
rect 10363 6972 10364 7036
rect 10428 6972 10429 7036
rect 10363 6971 10429 6972
rect 9259 4860 9325 4861
rect 9259 4796 9260 4860
rect 9324 4796 9325 4860
rect 9259 4795 9325 4796
rect 8891 3636 8957 3637
rect 8891 3572 8892 3636
rect 8956 3572 8957 3636
rect 8891 3571 8957 3572
rect 9814 3501 9874 6971
rect 10366 6357 10426 6971
rect 9995 6356 10061 6357
rect 9995 6292 9996 6356
rect 10060 6292 10061 6356
rect 9995 6291 10061 6292
rect 10363 6356 10429 6357
rect 10363 6292 10364 6356
rect 10428 6292 10429 6356
rect 10363 6291 10429 6292
rect 9998 4861 10058 6291
rect 10550 6221 10610 7110
rect 10363 6220 10429 6221
rect 10363 6156 10364 6220
rect 10428 6156 10429 6220
rect 10363 6155 10429 6156
rect 10547 6220 10613 6221
rect 10547 6156 10548 6220
rect 10612 6156 10613 6220
rect 10547 6155 10613 6156
rect 10179 5540 10245 5541
rect 10179 5476 10180 5540
rect 10244 5476 10245 5540
rect 10179 5475 10245 5476
rect 10182 4997 10242 5475
rect 10366 5405 10426 6155
rect 10547 5540 10613 5541
rect 10547 5476 10548 5540
rect 10612 5476 10613 5540
rect 10547 5475 10613 5476
rect 10363 5404 10429 5405
rect 10363 5340 10364 5404
rect 10428 5340 10429 5404
rect 10363 5339 10429 5340
rect 10179 4996 10245 4997
rect 10179 4932 10180 4996
rect 10244 4932 10245 4996
rect 10179 4931 10245 4932
rect 9995 4860 10061 4861
rect 9995 4796 9996 4860
rect 10060 4796 10061 4860
rect 9995 4795 10061 4796
rect 10550 4722 10610 5475
rect 10734 5130 10794 10779
rect 10918 9893 10978 18803
rect 11286 17237 11346 24243
rect 11654 19141 11714 29003
rect 12571 26348 12637 26349
rect 12571 26284 12572 26348
rect 12636 26284 12637 26348
rect 12571 26283 12637 26284
rect 12387 22132 12453 22133
rect 12387 22068 12388 22132
rect 12452 22130 12453 22132
rect 12574 22130 12634 26283
rect 12758 24173 12818 30363
rect 16251 30156 16317 30157
rect 16251 30092 16252 30156
rect 16316 30092 16317 30156
rect 16251 30091 16317 30092
rect 16254 28117 16314 30091
rect 19568 29408 19888 30432
rect 22691 30428 22757 30429
rect 22691 30364 22692 30428
rect 22756 30364 22757 30428
rect 22691 30363 22757 30364
rect 21587 30292 21653 30293
rect 21587 30228 21588 30292
rect 21652 30228 21653 30292
rect 21587 30227 21653 30228
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 16987 28388 17053 28389
rect 16987 28324 16988 28388
rect 17052 28324 17053 28388
rect 16987 28323 17053 28324
rect 16251 28116 16317 28117
rect 16251 28052 16252 28116
rect 16316 28052 16317 28116
rect 16251 28051 16317 28052
rect 14963 27708 15029 27709
rect 14963 27644 14964 27708
rect 15028 27644 15029 27708
rect 14963 27643 15029 27644
rect 14779 27572 14845 27573
rect 14779 27508 14780 27572
rect 14844 27508 14845 27572
rect 14779 27507 14845 27508
rect 13675 26620 13741 26621
rect 13675 26556 13676 26620
rect 13740 26556 13741 26620
rect 13675 26555 13741 26556
rect 12755 24172 12821 24173
rect 12755 24108 12756 24172
rect 12820 24108 12821 24172
rect 12755 24107 12821 24108
rect 12758 22133 12818 24107
rect 12939 23356 13005 23357
rect 12939 23292 12940 23356
rect 13004 23292 13005 23356
rect 12939 23291 13005 23292
rect 12942 22405 13002 23291
rect 12939 22404 13005 22405
rect 12939 22340 12940 22404
rect 13004 22340 13005 22404
rect 12939 22339 13005 22340
rect 13123 22404 13189 22405
rect 13123 22340 13124 22404
rect 13188 22340 13189 22404
rect 13123 22339 13189 22340
rect 12452 22070 12634 22130
rect 12755 22132 12821 22133
rect 12452 22068 12453 22070
rect 12387 22067 12453 22068
rect 12755 22068 12756 22132
rect 12820 22068 12821 22132
rect 12755 22067 12821 22068
rect 12755 21316 12821 21317
rect 12755 21252 12756 21316
rect 12820 21314 12821 21316
rect 13126 21314 13186 22339
rect 13491 21996 13557 21997
rect 13491 21932 13492 21996
rect 13556 21932 13557 21996
rect 13491 21931 13557 21932
rect 12820 21254 13186 21314
rect 12820 21252 12821 21254
rect 12755 21251 12821 21252
rect 11838 20710 12450 20770
rect 11838 20365 11898 20710
rect 12390 20637 12450 20710
rect 12203 20636 12269 20637
rect 12203 20572 12204 20636
rect 12268 20572 12269 20636
rect 12203 20571 12269 20572
rect 12387 20636 12453 20637
rect 12387 20572 12388 20636
rect 12452 20572 12453 20636
rect 12387 20571 12453 20572
rect 11835 20364 11901 20365
rect 11835 20300 11836 20364
rect 11900 20300 11901 20364
rect 11835 20299 11901 20300
rect 12206 19818 12266 20571
rect 12387 19820 12453 19821
rect 12387 19818 12388 19820
rect 12206 19758 12388 19818
rect 12387 19756 12388 19758
rect 12452 19756 12453 19820
rect 12387 19755 12453 19756
rect 11651 19140 11717 19141
rect 11651 19076 11652 19140
rect 11716 19076 11717 19140
rect 11651 19075 11717 19076
rect 12019 18596 12085 18597
rect 12019 18532 12020 18596
rect 12084 18532 12085 18596
rect 12019 18531 12085 18532
rect 11283 17236 11349 17237
rect 11283 17172 11284 17236
rect 11348 17172 11349 17236
rect 11283 17171 11349 17172
rect 11099 12340 11165 12341
rect 11099 12276 11100 12340
rect 11164 12276 11165 12340
rect 11099 12275 11165 12276
rect 11102 10301 11162 12275
rect 11099 10300 11165 10301
rect 11099 10236 11100 10300
rect 11164 10236 11165 10300
rect 11099 10235 11165 10236
rect 10915 9892 10981 9893
rect 10915 9828 10916 9892
rect 10980 9828 10981 9892
rect 10915 9827 10981 9828
rect 10918 7037 10978 9827
rect 11286 7853 11346 17171
rect 12022 15333 12082 18531
rect 12387 16420 12453 16421
rect 12387 16356 12388 16420
rect 12452 16356 12453 16420
rect 12387 16355 12453 16356
rect 12019 15332 12085 15333
rect 12019 15268 12020 15332
rect 12084 15268 12085 15332
rect 12019 15267 12085 15268
rect 12203 15196 12269 15197
rect 12203 15132 12204 15196
rect 12268 15132 12269 15196
rect 12203 15131 12269 15132
rect 11467 12476 11533 12477
rect 11467 12412 11468 12476
rect 11532 12412 11533 12476
rect 11467 12411 11533 12412
rect 11470 11661 11530 12411
rect 11467 11660 11533 11661
rect 11467 11596 11468 11660
rect 11532 11596 11533 11660
rect 11467 11595 11533 11596
rect 11470 9893 11530 11595
rect 11467 9892 11533 9893
rect 11467 9828 11468 9892
rect 11532 9828 11533 9892
rect 11467 9827 11533 9828
rect 12206 9077 12266 15131
rect 12390 11661 12450 16355
rect 13123 13156 13189 13157
rect 13123 13092 13124 13156
rect 13188 13092 13189 13156
rect 13123 13091 13189 13092
rect 13126 12450 13186 13091
rect 13126 12390 13370 12450
rect 12387 11660 12453 11661
rect 12387 11596 12388 11660
rect 12452 11596 12453 11660
rect 12387 11595 12453 11596
rect 13123 11388 13189 11389
rect 13123 11324 13124 11388
rect 13188 11324 13189 11388
rect 13123 11323 13189 11324
rect 12939 10844 13005 10845
rect 12939 10780 12940 10844
rect 13004 10780 13005 10844
rect 12939 10779 13005 10780
rect 12942 10029 13002 10779
rect 12939 10028 13005 10029
rect 12939 9964 12940 10028
rect 13004 9964 13005 10028
rect 12939 9963 13005 9964
rect 12019 9076 12085 9077
rect 12019 9012 12020 9076
rect 12084 9012 12085 9076
rect 12019 9011 12085 9012
rect 12203 9076 12269 9077
rect 12203 9012 12204 9076
rect 12268 9012 12269 9076
rect 12203 9011 12269 9012
rect 11467 8668 11533 8669
rect 11467 8604 11468 8668
rect 11532 8604 11533 8668
rect 11467 8603 11533 8604
rect 11283 7852 11349 7853
rect 11283 7788 11284 7852
rect 11348 7788 11349 7852
rect 11470 7850 11530 8603
rect 12022 7986 12082 9011
rect 12203 7988 12269 7989
rect 12203 7986 12204 7988
rect 12022 7926 12204 7986
rect 12203 7924 12204 7926
rect 12268 7924 12269 7988
rect 12203 7923 12269 7924
rect 11470 7790 12450 7850
rect 11283 7787 11349 7788
rect 10915 7036 10981 7037
rect 10915 6972 10916 7036
rect 10980 6972 10981 7036
rect 10915 6971 10981 6972
rect 11651 7036 11717 7037
rect 11651 6972 11652 7036
rect 11716 6972 11717 7036
rect 11651 6971 11717 6972
rect 11654 5538 11714 6971
rect 12203 6764 12269 6765
rect 12203 6700 12204 6764
rect 12268 6700 12269 6764
rect 12203 6699 12269 6700
rect 12206 5949 12266 6699
rect 12390 6629 12450 7790
rect 12387 6628 12453 6629
rect 12387 6564 12388 6628
rect 12452 6564 12453 6628
rect 12387 6563 12453 6564
rect 12203 5948 12269 5949
rect 12203 5884 12204 5948
rect 12268 5884 12269 5948
rect 12203 5883 12269 5884
rect 12387 5948 12453 5949
rect 12387 5884 12388 5948
rect 12452 5884 12453 5948
rect 12387 5883 12453 5884
rect 12390 5810 12450 5883
rect 12206 5750 12450 5810
rect 12206 5677 12266 5750
rect 12203 5676 12269 5677
rect 12203 5612 12204 5676
rect 12268 5612 12269 5676
rect 12203 5611 12269 5612
rect 12755 5676 12821 5677
rect 12755 5612 12756 5676
rect 12820 5612 12821 5676
rect 12755 5611 12821 5612
rect 12758 5538 12818 5611
rect 11654 5478 12818 5538
rect 10734 5070 12082 5130
rect 12022 4997 12082 5070
rect 12019 4996 12085 4997
rect 12019 4932 12020 4996
rect 12084 4932 12085 4996
rect 12019 4931 12085 4932
rect 13126 4861 13186 11323
rect 13123 4860 13189 4861
rect 13123 4796 13124 4860
rect 13188 4796 13189 4860
rect 13123 4795 13189 4796
rect 12387 4724 12453 4725
rect 12387 4722 12388 4724
rect 10550 4662 12388 4722
rect 12387 4660 12388 4662
rect 12452 4660 12453 4724
rect 12387 4659 12453 4660
rect 12571 4724 12637 4725
rect 12571 4660 12572 4724
rect 12636 4660 12637 4724
rect 13310 4722 13370 12390
rect 13494 10845 13554 21931
rect 13491 10844 13557 10845
rect 13491 10780 13492 10844
rect 13556 10780 13557 10844
rect 13491 10779 13557 10780
rect 13678 8261 13738 26555
rect 13859 24988 13925 24989
rect 13859 24924 13860 24988
rect 13924 24924 13925 24988
rect 13859 24923 13925 24924
rect 13862 18053 13922 24923
rect 14595 21452 14661 21453
rect 14595 21388 14596 21452
rect 14660 21388 14661 21452
rect 14595 21387 14661 21388
rect 13859 18052 13925 18053
rect 13859 17988 13860 18052
rect 13924 17988 13925 18052
rect 13859 17987 13925 17988
rect 13862 17373 13922 17987
rect 13859 17372 13925 17373
rect 13859 17308 13860 17372
rect 13924 17308 13925 17372
rect 13859 17307 13925 17308
rect 14598 15877 14658 21387
rect 14782 18461 14842 27507
rect 14779 18460 14845 18461
rect 14779 18396 14780 18460
rect 14844 18396 14845 18460
rect 14779 18395 14845 18396
rect 14966 16829 15026 27643
rect 16067 26892 16133 26893
rect 16067 26828 16068 26892
rect 16132 26828 16133 26892
rect 16067 26827 16133 26828
rect 15515 25668 15581 25669
rect 15515 25604 15516 25668
rect 15580 25604 15581 25668
rect 15515 25603 15581 25604
rect 15518 20773 15578 25603
rect 15515 20772 15581 20773
rect 15515 20708 15516 20772
rect 15580 20708 15581 20772
rect 15515 20707 15581 20708
rect 16070 17917 16130 26827
rect 16067 17916 16133 17917
rect 16067 17852 16068 17916
rect 16132 17852 16133 17916
rect 16067 17851 16133 17852
rect 14963 16828 15029 16829
rect 14963 16764 14964 16828
rect 15028 16764 15029 16828
rect 14963 16763 15029 16764
rect 13859 15876 13925 15877
rect 13859 15812 13860 15876
rect 13924 15812 13925 15876
rect 13859 15811 13925 15812
rect 14595 15876 14661 15877
rect 14595 15812 14596 15876
rect 14660 15812 14661 15876
rect 14595 15811 14661 15812
rect 13862 10165 13922 15811
rect 14779 15468 14845 15469
rect 14779 15404 14780 15468
rect 14844 15404 14845 15468
rect 14779 15403 14845 15404
rect 14782 14517 14842 15403
rect 14779 14516 14845 14517
rect 14779 14452 14780 14516
rect 14844 14452 14845 14516
rect 14779 14451 14845 14452
rect 15883 14516 15949 14517
rect 15883 14452 15884 14516
rect 15948 14452 15949 14516
rect 15883 14451 15949 14452
rect 14963 14108 15029 14109
rect 14963 14044 14964 14108
rect 15028 14044 15029 14108
rect 14963 14043 15029 14044
rect 14779 13564 14845 13565
rect 14779 13500 14780 13564
rect 14844 13500 14845 13564
rect 14779 13499 14845 13500
rect 14227 13428 14293 13429
rect 14227 13364 14228 13428
rect 14292 13364 14293 13428
rect 14227 13363 14293 13364
rect 14230 11250 14290 13363
rect 14230 11190 14658 11250
rect 14411 10980 14477 10981
rect 14411 10916 14412 10980
rect 14476 10916 14477 10980
rect 14411 10915 14477 10916
rect 14227 10708 14293 10709
rect 14227 10644 14228 10708
rect 14292 10644 14293 10708
rect 14227 10643 14293 10644
rect 13859 10164 13925 10165
rect 13859 10100 13860 10164
rect 13924 10100 13925 10164
rect 13859 10099 13925 10100
rect 13675 8260 13741 8261
rect 13675 8196 13676 8260
rect 13740 8196 13741 8260
rect 13675 8195 13741 8196
rect 13862 5541 13922 10099
rect 14043 8396 14109 8397
rect 14043 8332 14044 8396
rect 14108 8332 14109 8396
rect 14043 8331 14109 8332
rect 14046 5541 14106 8331
rect 13859 5540 13925 5541
rect 13859 5476 13860 5540
rect 13924 5476 13925 5540
rect 13859 5475 13925 5476
rect 14043 5540 14109 5541
rect 14043 5476 14044 5540
rect 14108 5476 14109 5540
rect 14043 5475 14109 5476
rect 13491 4724 13557 4725
rect 13491 4722 13492 4724
rect 13310 4662 13492 4722
rect 12571 4659 12637 4660
rect 13491 4660 13492 4662
rect 13556 4660 13557 4724
rect 13491 4659 13557 4660
rect 12574 4314 12634 4659
rect 12022 4254 12634 4314
rect 12022 4181 12082 4254
rect 12019 4180 12085 4181
rect 12019 4116 12020 4180
rect 12084 4116 12085 4180
rect 12019 4115 12085 4116
rect 14230 4045 14290 10643
rect 14414 9757 14474 10915
rect 14411 9756 14477 9757
rect 14411 9692 14412 9756
rect 14476 9692 14477 9756
rect 14411 9691 14477 9692
rect 14598 8397 14658 11190
rect 14595 8396 14661 8397
rect 14595 8332 14596 8396
rect 14660 8332 14661 8396
rect 14595 8331 14661 8332
rect 14782 4861 14842 13499
rect 14966 10437 15026 14043
rect 15699 13020 15765 13021
rect 15699 12956 15700 13020
rect 15764 12956 15765 13020
rect 15699 12955 15765 12956
rect 14963 10436 15029 10437
rect 14963 10372 14964 10436
rect 15028 10372 15029 10436
rect 14963 10371 15029 10372
rect 15515 9756 15581 9757
rect 15515 9692 15516 9756
rect 15580 9692 15581 9756
rect 15515 9691 15581 9692
rect 15518 6085 15578 9691
rect 15702 6901 15762 12955
rect 15886 8397 15946 14451
rect 16067 9348 16133 9349
rect 16067 9284 16068 9348
rect 16132 9284 16133 9348
rect 16067 9283 16133 9284
rect 15883 8396 15949 8397
rect 15883 8332 15884 8396
rect 15948 8332 15949 8396
rect 15883 8331 15949 8332
rect 15699 6900 15765 6901
rect 15699 6836 15700 6900
rect 15764 6836 15765 6900
rect 15699 6835 15765 6836
rect 15515 6084 15581 6085
rect 15515 6020 15516 6084
rect 15580 6020 15581 6084
rect 15515 6019 15581 6020
rect 14779 4860 14845 4861
rect 14779 4796 14780 4860
rect 14844 4796 14845 4860
rect 14779 4795 14845 4796
rect 15699 4724 15765 4725
rect 15699 4660 15700 4724
rect 15764 4660 15765 4724
rect 15699 4659 15765 4660
rect 15702 4453 15762 4659
rect 15699 4452 15765 4453
rect 15699 4388 15700 4452
rect 15764 4388 15765 4452
rect 15699 4387 15765 4388
rect 14227 4044 14293 4045
rect 14227 3980 14228 4044
rect 14292 3980 14293 4044
rect 14227 3979 14293 3980
rect 16070 3909 16130 9283
rect 16067 3908 16133 3909
rect 16067 3844 16068 3908
rect 16132 3844 16133 3908
rect 16067 3843 16133 3844
rect 9811 3500 9877 3501
rect 9811 3436 9812 3500
rect 9876 3436 9877 3500
rect 9811 3435 9877 3436
rect 16254 3229 16314 28051
rect 16803 24036 16869 24037
rect 16803 23972 16804 24036
rect 16868 23972 16869 24036
rect 16803 23971 16869 23972
rect 16806 18053 16866 23971
rect 16990 22813 17050 28323
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 17723 26348 17789 26349
rect 17723 26284 17724 26348
rect 17788 26284 17789 26348
rect 17723 26283 17789 26284
rect 16987 22812 17053 22813
rect 16987 22748 16988 22812
rect 17052 22748 17053 22812
rect 16987 22747 17053 22748
rect 17355 20364 17421 20365
rect 17355 20300 17356 20364
rect 17420 20300 17421 20364
rect 17355 20299 17421 20300
rect 16803 18052 16869 18053
rect 16803 17988 16804 18052
rect 16868 17988 16869 18052
rect 16803 17987 16869 17988
rect 17171 18052 17237 18053
rect 17171 17988 17172 18052
rect 17236 17988 17237 18052
rect 17171 17987 17237 17988
rect 16619 13972 16685 13973
rect 16619 13908 16620 13972
rect 16684 13908 16685 13972
rect 16619 13907 16685 13908
rect 16622 12477 16682 13907
rect 16806 12749 16866 17987
rect 16987 17780 17053 17781
rect 16987 17716 16988 17780
rect 17052 17716 17053 17780
rect 16987 17715 17053 17716
rect 16803 12748 16869 12749
rect 16803 12684 16804 12748
rect 16868 12684 16869 12748
rect 16803 12683 16869 12684
rect 16619 12476 16685 12477
rect 16619 12412 16620 12476
rect 16684 12412 16685 12476
rect 16619 12411 16685 12412
rect 16435 10436 16501 10437
rect 16435 10372 16436 10436
rect 16500 10372 16501 10436
rect 16435 10371 16501 10372
rect 16438 8805 16498 10371
rect 16619 10028 16685 10029
rect 16619 9964 16620 10028
rect 16684 9964 16685 10028
rect 16619 9963 16685 9964
rect 16435 8804 16501 8805
rect 16435 8740 16436 8804
rect 16500 8740 16501 8804
rect 16435 8739 16501 8740
rect 16622 7581 16682 9963
rect 16803 7988 16869 7989
rect 16803 7924 16804 7988
rect 16868 7924 16869 7988
rect 16803 7923 16869 7924
rect 16806 7717 16866 7923
rect 16803 7716 16869 7717
rect 16803 7652 16804 7716
rect 16868 7652 16869 7716
rect 16803 7651 16869 7652
rect 16619 7580 16685 7581
rect 16619 7516 16620 7580
rect 16684 7516 16685 7580
rect 16619 7515 16685 7516
rect 16990 5949 17050 17715
rect 17174 7717 17234 17987
rect 17358 17101 17418 20299
rect 17726 18733 17786 26283
rect 19568 26144 19888 27168
rect 20115 26348 20181 26349
rect 20115 26284 20116 26348
rect 20180 26284 20181 26348
rect 20115 26283 20181 26284
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 20118 24445 20178 26283
rect 20115 24444 20181 24445
rect 20115 24380 20116 24444
rect 20180 24380 20181 24444
rect 20115 24379 20181 24380
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 18827 21452 18893 21453
rect 18827 21388 18828 21452
rect 18892 21388 18893 21452
rect 18827 21387 18893 21388
rect 19198 21390 19442 21450
rect 18830 19957 18890 21387
rect 19198 21181 19258 21390
rect 19195 21180 19261 21181
rect 19195 21116 19196 21180
rect 19260 21116 19261 21180
rect 19195 21115 19261 21116
rect 19195 21044 19261 21045
rect 19195 20980 19196 21044
rect 19260 20980 19261 21044
rect 19195 20979 19261 20980
rect 18827 19956 18893 19957
rect 18827 19892 18828 19956
rect 18892 19892 18893 19956
rect 18827 19891 18893 19892
rect 17723 18732 17789 18733
rect 17723 18668 17724 18732
rect 17788 18668 17789 18732
rect 17723 18667 17789 18668
rect 17539 17508 17605 17509
rect 17539 17444 17540 17508
rect 17604 17444 17605 17508
rect 17539 17443 17605 17444
rect 17355 17100 17421 17101
rect 17355 17036 17356 17100
rect 17420 17036 17421 17100
rect 17355 17035 17421 17036
rect 17355 15468 17421 15469
rect 17355 15404 17356 15468
rect 17420 15404 17421 15468
rect 17355 15403 17421 15404
rect 17358 8669 17418 15403
rect 17542 11389 17602 17443
rect 18275 17236 18341 17237
rect 18275 17172 18276 17236
rect 18340 17172 18341 17236
rect 18275 17171 18341 17172
rect 18827 17236 18893 17237
rect 18827 17172 18828 17236
rect 18892 17172 18893 17236
rect 18827 17171 18893 17172
rect 17907 15740 17973 15741
rect 17907 15676 17908 15740
rect 17972 15676 17973 15740
rect 17907 15675 17973 15676
rect 18091 15740 18157 15741
rect 18091 15676 18092 15740
rect 18156 15676 18157 15740
rect 18091 15675 18157 15676
rect 17910 15469 17970 15675
rect 17907 15468 17973 15469
rect 17907 15404 17908 15468
rect 17972 15404 17973 15468
rect 17907 15403 17973 15404
rect 18094 12749 18154 15675
rect 18278 14786 18338 17171
rect 18459 15332 18525 15333
rect 18459 15268 18460 15332
rect 18524 15268 18525 15332
rect 18459 15267 18525 15268
rect 18462 14922 18522 15267
rect 18830 15197 18890 17171
rect 19011 17100 19077 17101
rect 19011 17036 19012 17100
rect 19076 17036 19077 17100
rect 19011 17035 19077 17036
rect 18827 15196 18893 15197
rect 18827 15132 18828 15196
rect 18892 15132 18893 15196
rect 18827 15131 18893 15132
rect 18462 14862 18890 14922
rect 18278 14726 18706 14786
rect 18459 14652 18525 14653
rect 18459 14588 18460 14652
rect 18524 14588 18525 14652
rect 18459 14587 18525 14588
rect 18462 14109 18522 14587
rect 18459 14108 18525 14109
rect 18459 14044 18460 14108
rect 18524 14044 18525 14108
rect 18459 14043 18525 14044
rect 18091 12748 18157 12749
rect 18091 12684 18092 12748
rect 18156 12684 18157 12748
rect 18091 12683 18157 12684
rect 17723 11660 17789 11661
rect 17723 11596 17724 11660
rect 17788 11658 17789 11660
rect 18275 11660 18341 11661
rect 17788 11598 18154 11658
rect 17788 11596 17789 11598
rect 17723 11595 17789 11596
rect 17539 11388 17605 11389
rect 17539 11324 17540 11388
rect 17604 11324 17605 11388
rect 17539 11323 17605 11324
rect 17723 11388 17789 11389
rect 17723 11324 17724 11388
rect 17788 11324 17789 11388
rect 17723 11323 17789 11324
rect 17726 10573 17786 11323
rect 17907 10980 17973 10981
rect 17907 10916 17908 10980
rect 17972 10916 17973 10980
rect 17907 10915 17973 10916
rect 17910 10573 17970 10915
rect 17723 10572 17789 10573
rect 17723 10508 17724 10572
rect 17788 10508 17789 10572
rect 17723 10507 17789 10508
rect 17907 10572 17973 10573
rect 17907 10508 17908 10572
rect 17972 10508 17973 10572
rect 17907 10507 17973 10508
rect 18094 10434 18154 11598
rect 18275 11596 18276 11660
rect 18340 11596 18341 11660
rect 18275 11595 18341 11596
rect 17726 10374 18154 10434
rect 17539 10164 17605 10165
rect 17539 10100 17540 10164
rect 17604 10100 17605 10164
rect 17539 10099 17605 10100
rect 17542 9210 17602 10099
rect 17726 9690 17786 10374
rect 17726 9630 17970 9690
rect 17542 9150 17786 9210
rect 17539 9076 17605 9077
rect 17539 9012 17540 9076
rect 17604 9012 17605 9076
rect 17539 9011 17605 9012
rect 17355 8668 17421 8669
rect 17355 8604 17356 8668
rect 17420 8604 17421 8668
rect 17355 8603 17421 8604
rect 17355 8124 17421 8125
rect 17355 8060 17356 8124
rect 17420 8060 17421 8124
rect 17355 8059 17421 8060
rect 17171 7716 17237 7717
rect 17171 7652 17172 7716
rect 17236 7652 17237 7716
rect 17171 7651 17237 7652
rect 16987 5948 17053 5949
rect 16987 5884 16988 5948
rect 17052 5884 17053 5948
rect 16987 5883 17053 5884
rect 17358 4725 17418 8059
rect 17355 4724 17421 4725
rect 17355 4660 17356 4724
rect 17420 4660 17421 4724
rect 17355 4659 17421 4660
rect 17542 4045 17602 9011
rect 17726 7717 17786 9150
rect 17723 7716 17789 7717
rect 17723 7652 17724 7716
rect 17788 7652 17789 7716
rect 17723 7651 17789 7652
rect 17723 6628 17789 6629
rect 17723 6564 17724 6628
rect 17788 6564 17789 6628
rect 17723 6563 17789 6564
rect 17726 5677 17786 6563
rect 17910 6357 17970 9630
rect 18091 9076 18157 9077
rect 18091 9012 18092 9076
rect 18156 9012 18157 9076
rect 18091 9011 18157 9012
rect 18094 6626 18154 9011
rect 18278 6765 18338 11595
rect 18462 9210 18522 14043
rect 18646 11117 18706 14726
rect 18830 14245 18890 14862
rect 18827 14244 18893 14245
rect 18827 14180 18828 14244
rect 18892 14180 18893 14244
rect 18827 14179 18893 14180
rect 18827 14108 18893 14109
rect 18827 14044 18828 14108
rect 18892 14044 18893 14108
rect 18827 14043 18893 14044
rect 18643 11116 18709 11117
rect 18643 11052 18644 11116
rect 18708 11052 18709 11116
rect 18643 11051 18709 11052
rect 18643 10980 18709 10981
rect 18643 10916 18644 10980
rect 18708 10916 18709 10980
rect 18643 10915 18709 10916
rect 18646 9757 18706 10915
rect 18643 9756 18709 9757
rect 18643 9692 18644 9756
rect 18708 9692 18709 9756
rect 18643 9691 18709 9692
rect 18462 9150 18706 9210
rect 18646 7037 18706 9150
rect 18459 7036 18525 7037
rect 18459 6972 18460 7036
rect 18524 6972 18525 7036
rect 18459 6971 18525 6972
rect 18643 7036 18709 7037
rect 18643 6972 18644 7036
rect 18708 6972 18709 7036
rect 18643 6971 18709 6972
rect 18275 6764 18341 6765
rect 18275 6700 18276 6764
rect 18340 6700 18341 6764
rect 18275 6699 18341 6700
rect 18094 6566 18338 6626
rect 17907 6356 17973 6357
rect 17907 6292 17908 6356
rect 17972 6292 17973 6356
rect 17907 6291 17973 6292
rect 17723 5676 17789 5677
rect 17723 5612 17724 5676
rect 17788 5612 17789 5676
rect 17723 5611 17789 5612
rect 18091 5676 18157 5677
rect 18091 5612 18092 5676
rect 18156 5612 18157 5676
rect 18091 5611 18157 5612
rect 18094 4317 18154 5611
rect 18278 5133 18338 6566
rect 18275 5132 18341 5133
rect 18275 5068 18276 5132
rect 18340 5068 18341 5132
rect 18275 5067 18341 5068
rect 18091 4316 18157 4317
rect 18091 4252 18092 4316
rect 18156 4252 18157 4316
rect 18091 4251 18157 4252
rect 17539 4044 17605 4045
rect 17539 3980 17540 4044
rect 17604 3980 17605 4044
rect 17539 3979 17605 3980
rect 16251 3228 16317 3229
rect 16251 3164 16252 3228
rect 16316 3164 16317 3228
rect 16251 3163 16317 3164
rect 18462 3090 18522 6971
rect 18643 6764 18709 6765
rect 18643 6700 18644 6764
rect 18708 6700 18709 6764
rect 18643 6699 18709 6700
rect 18646 3773 18706 6699
rect 18830 5405 18890 14043
rect 19014 13157 19074 17035
rect 19198 14789 19258 20979
rect 19195 14788 19261 14789
rect 19195 14724 19196 14788
rect 19260 14724 19261 14788
rect 19195 14723 19261 14724
rect 19382 14245 19442 21390
rect 19568 20704 19888 21728
rect 20115 20772 20181 20773
rect 20115 20708 20116 20772
rect 20180 20708 20181 20772
rect 20115 20707 20181 20708
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 20118 19821 20178 20707
rect 20483 20500 20549 20501
rect 20483 20436 20484 20500
rect 20548 20436 20549 20500
rect 20483 20435 20549 20436
rect 20115 19820 20181 19821
rect 20115 19756 20116 19820
rect 20180 19756 20181 19820
rect 20115 19755 20181 19756
rect 20115 19684 20181 19685
rect 20115 19620 20116 19684
rect 20180 19620 20181 19684
rect 20115 19619 20181 19620
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 20118 19413 20178 19619
rect 20115 19412 20181 19413
rect 20115 19348 20116 19412
rect 20180 19348 20181 19412
rect 20115 19347 20181 19348
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 20115 17780 20181 17781
rect 20115 17716 20116 17780
rect 20180 17778 20181 17780
rect 20180 17718 20362 17778
rect 20180 17716 20181 17718
rect 20115 17715 20181 17716
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19195 14244 19261 14245
rect 19195 14180 19196 14244
rect 19260 14180 19261 14244
rect 19195 14179 19261 14180
rect 19379 14244 19445 14245
rect 19379 14180 19380 14244
rect 19444 14180 19445 14244
rect 19379 14179 19445 14180
rect 19011 13156 19077 13157
rect 19011 13092 19012 13156
rect 19076 13092 19077 13156
rect 19011 13091 19077 13092
rect 19011 12884 19077 12885
rect 19011 12820 19012 12884
rect 19076 12820 19077 12884
rect 19011 12819 19077 12820
rect 19014 8261 19074 12819
rect 19198 10981 19258 14179
rect 19568 14176 19888 15200
rect 20115 15196 20181 15197
rect 20115 15132 20116 15196
rect 20180 15132 20181 15196
rect 20115 15131 20181 15132
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 20118 13021 20178 15131
rect 20115 13020 20181 13021
rect 20115 12956 20116 13020
rect 20180 12956 20181 13020
rect 20115 12955 20181 12956
rect 20115 12340 20181 12341
rect 20115 12276 20116 12340
rect 20180 12276 20181 12340
rect 20115 12275 20181 12276
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19379 11932 19445 11933
rect 19379 11868 19380 11932
rect 19444 11868 19445 11932
rect 19379 11867 19445 11868
rect 19195 10980 19261 10981
rect 19195 10916 19196 10980
rect 19260 10916 19261 10980
rect 19195 10915 19261 10916
rect 19382 10845 19442 11867
rect 19568 10912 19888 11936
rect 20118 11933 20178 12275
rect 20115 11932 20181 11933
rect 20115 11868 20116 11932
rect 20180 11868 20181 11932
rect 20115 11867 20181 11868
rect 19977 11524 20043 11525
rect 19977 11460 19978 11524
rect 20042 11522 20043 11524
rect 20042 11462 20178 11522
rect 20042 11460 20043 11462
rect 19977 11459 20043 11460
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19379 10844 19445 10845
rect 19379 10780 19380 10844
rect 19444 10780 19445 10844
rect 19379 10779 19445 10780
rect 19568 9824 19888 10848
rect 20118 10845 20178 11462
rect 20115 10844 20181 10845
rect 20115 10780 20116 10844
rect 20180 10780 20181 10844
rect 20115 10779 20181 10780
rect 20115 10164 20181 10165
rect 20115 10100 20116 10164
rect 20180 10100 20181 10164
rect 20115 10099 20181 10100
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19379 9756 19445 9757
rect 19379 9692 19380 9756
rect 19444 9692 19445 9756
rect 19379 9691 19445 9692
rect 19195 8804 19261 8805
rect 19195 8740 19196 8804
rect 19260 8740 19261 8804
rect 19195 8739 19261 8740
rect 19011 8260 19077 8261
rect 19011 8196 19012 8260
rect 19076 8196 19077 8260
rect 19011 8195 19077 8196
rect 19198 7714 19258 8739
rect 19382 7853 19442 9691
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19379 7852 19445 7853
rect 19379 7788 19380 7852
rect 19444 7788 19445 7852
rect 19379 7787 19445 7788
rect 19014 7654 19258 7714
rect 19014 6493 19074 7654
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19195 7580 19261 7581
rect 19195 7516 19196 7580
rect 19260 7516 19261 7580
rect 19195 7515 19261 7516
rect 19198 7037 19258 7515
rect 19195 7036 19261 7037
rect 19195 6972 19196 7036
rect 19260 6972 19261 7036
rect 19195 6971 19261 6972
rect 19568 6560 19888 7584
rect 20118 6629 20178 10099
rect 20302 7581 20362 17718
rect 20486 16693 20546 20435
rect 20667 20092 20733 20093
rect 20667 20028 20668 20092
rect 20732 20028 20733 20092
rect 20667 20027 20733 20028
rect 20670 19821 20730 20027
rect 20667 19820 20733 19821
rect 20667 19756 20668 19820
rect 20732 19756 20733 19820
rect 20667 19755 20733 19756
rect 21035 18324 21101 18325
rect 21035 18260 21036 18324
rect 21100 18260 21101 18324
rect 21035 18259 21101 18260
rect 20483 16692 20549 16693
rect 20483 16628 20484 16692
rect 20548 16628 20549 16692
rect 20483 16627 20549 16628
rect 20851 16692 20917 16693
rect 20851 16628 20852 16692
rect 20916 16628 20917 16692
rect 20851 16627 20917 16628
rect 20854 16149 20914 16627
rect 20851 16148 20917 16149
rect 20851 16084 20852 16148
rect 20916 16084 20917 16148
rect 20851 16083 20917 16084
rect 20851 15332 20917 15333
rect 20851 15268 20852 15332
rect 20916 15268 20917 15332
rect 20851 15267 20917 15268
rect 20854 13834 20914 15267
rect 21038 14789 21098 18259
rect 21219 17916 21285 17917
rect 21219 17852 21220 17916
rect 21284 17852 21285 17916
rect 21219 17851 21285 17852
rect 21222 17509 21282 17851
rect 21219 17508 21285 17509
rect 21219 17444 21220 17508
rect 21284 17444 21285 17508
rect 21219 17443 21285 17444
rect 21219 17100 21285 17101
rect 21219 17036 21220 17100
rect 21284 17036 21285 17100
rect 21219 17035 21285 17036
rect 21035 14788 21101 14789
rect 21035 14724 21036 14788
rect 21100 14724 21101 14788
rect 21035 14723 21101 14724
rect 21035 14516 21101 14517
rect 21035 14452 21036 14516
rect 21100 14452 21101 14516
rect 21035 14451 21101 14452
rect 20670 13774 20914 13834
rect 20670 12069 20730 13774
rect 21038 13701 21098 14451
rect 21035 13700 21101 13701
rect 21035 13636 21036 13700
rect 21100 13636 21101 13700
rect 21035 13635 21101 13636
rect 21035 12884 21101 12885
rect 21035 12820 21036 12884
rect 21100 12820 21101 12884
rect 21035 12819 21101 12820
rect 20667 12068 20733 12069
rect 20667 12004 20668 12068
rect 20732 12004 20733 12068
rect 20667 12003 20733 12004
rect 20483 11388 20549 11389
rect 20483 11324 20484 11388
rect 20548 11386 20549 11388
rect 20548 11326 20730 11386
rect 20548 11324 20549 11326
rect 20483 11323 20549 11324
rect 20483 9484 20549 9485
rect 20483 9420 20484 9484
rect 20548 9420 20549 9484
rect 20483 9419 20549 9420
rect 20486 8805 20546 9419
rect 20483 8804 20549 8805
rect 20483 8740 20484 8804
rect 20548 8740 20549 8804
rect 20483 8739 20549 8740
rect 20670 8125 20730 11326
rect 20851 10164 20917 10165
rect 20851 10100 20852 10164
rect 20916 10100 20917 10164
rect 20851 10099 20917 10100
rect 20667 8124 20733 8125
rect 20667 8060 20668 8124
rect 20732 8060 20733 8124
rect 20667 8059 20733 8060
rect 20299 7580 20365 7581
rect 20299 7516 20300 7580
rect 20364 7516 20365 7580
rect 20299 7515 20365 7516
rect 20299 7036 20365 7037
rect 20299 6972 20300 7036
rect 20364 6972 20365 7036
rect 20299 6971 20365 6972
rect 20115 6628 20181 6629
rect 20115 6564 20116 6628
rect 20180 6564 20181 6628
rect 20115 6563 20181 6564
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19011 6492 19077 6493
rect 19011 6428 19012 6492
rect 19076 6428 19077 6492
rect 19011 6427 19077 6428
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 18827 5404 18893 5405
rect 18827 5340 18828 5404
rect 18892 5340 18893 5404
rect 18827 5339 18893 5340
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 18643 3772 18709 3773
rect 18643 3708 18644 3772
rect 18708 3708 18709 3772
rect 18643 3707 18709 3708
rect 18827 3772 18893 3773
rect 18827 3708 18828 3772
rect 18892 3708 18893 3772
rect 18827 3707 18893 3708
rect 18830 3090 18890 3707
rect 18462 3030 18890 3090
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 8339 2684 8405 2685
rect 8339 2620 8340 2684
rect 8404 2620 8405 2684
rect 8339 2619 8405 2620
rect 5211 2548 5277 2549
rect 5211 2484 5212 2548
rect 5276 2484 5277 2548
rect 5211 2483 5277 2484
rect 19568 2208 19888 3232
rect 20302 2549 20362 6971
rect 20854 6765 20914 10099
rect 20851 6764 20917 6765
rect 20851 6700 20852 6764
rect 20916 6700 20917 6764
rect 20851 6699 20917 6700
rect 21038 6493 21098 12819
rect 21222 6629 21282 17035
rect 21403 13700 21469 13701
rect 21403 13636 21404 13700
rect 21468 13636 21469 13700
rect 21403 13635 21469 13636
rect 21406 11525 21466 13635
rect 21590 11797 21650 30227
rect 21955 28932 22021 28933
rect 21955 28868 21956 28932
rect 22020 28868 22021 28932
rect 21955 28867 22021 28868
rect 21771 23492 21837 23493
rect 21771 23428 21772 23492
rect 21836 23428 21837 23492
rect 21771 23427 21837 23428
rect 21587 11796 21653 11797
rect 21587 11732 21588 11796
rect 21652 11732 21653 11796
rect 21587 11731 21653 11732
rect 21403 11524 21469 11525
rect 21403 11460 21404 11524
rect 21468 11460 21469 11524
rect 21403 11459 21469 11460
rect 21406 7853 21466 11459
rect 21403 7852 21469 7853
rect 21403 7788 21404 7852
rect 21468 7788 21469 7852
rect 21403 7787 21469 7788
rect 21219 6628 21285 6629
rect 21219 6564 21220 6628
rect 21284 6564 21285 6628
rect 21219 6563 21285 6564
rect 21035 6492 21101 6493
rect 21035 6428 21036 6492
rect 21100 6428 21101 6492
rect 21035 6427 21101 6428
rect 20299 2548 20365 2549
rect 20299 2484 20300 2548
rect 20364 2484 20365 2548
rect 20299 2483 20365 2484
rect 21590 2413 21650 11731
rect 21774 2549 21834 23427
rect 21958 4045 22018 28867
rect 22694 22133 22754 30363
rect 23059 25940 23125 25941
rect 23059 25876 23060 25940
rect 23124 25876 23125 25940
rect 23059 25875 23125 25876
rect 22875 25668 22941 25669
rect 22875 25604 22876 25668
rect 22940 25604 22941 25668
rect 22875 25603 22941 25604
rect 22691 22132 22757 22133
rect 22691 22068 22692 22132
rect 22756 22068 22757 22132
rect 22691 22067 22757 22068
rect 22139 18324 22205 18325
rect 22139 18260 22140 18324
rect 22204 18260 22205 18324
rect 22139 18259 22205 18260
rect 22142 17509 22202 18259
rect 22139 17508 22205 17509
rect 22139 17444 22140 17508
rect 22204 17444 22205 17508
rect 22139 17443 22205 17444
rect 22323 17508 22389 17509
rect 22323 17444 22324 17508
rect 22388 17444 22389 17508
rect 22323 17443 22389 17444
rect 22326 12069 22386 17443
rect 22507 14788 22573 14789
rect 22507 14724 22508 14788
rect 22572 14724 22573 14788
rect 22507 14723 22573 14724
rect 22323 12068 22389 12069
rect 22323 12004 22324 12068
rect 22388 12004 22389 12068
rect 22323 12003 22389 12004
rect 22323 11524 22389 11525
rect 22323 11460 22324 11524
rect 22388 11460 22389 11524
rect 22323 11459 22389 11460
rect 22139 9756 22205 9757
rect 22139 9692 22140 9756
rect 22204 9692 22205 9756
rect 22139 9691 22205 9692
rect 22142 7309 22202 9691
rect 22139 7308 22205 7309
rect 22139 7244 22140 7308
rect 22204 7244 22205 7308
rect 22139 7243 22205 7244
rect 22326 6765 22386 11459
rect 22510 7173 22570 14723
rect 22878 11933 22938 25603
rect 22875 11932 22941 11933
rect 22875 11868 22876 11932
rect 22940 11868 22941 11932
rect 22875 11867 22941 11868
rect 22507 7172 22573 7173
rect 22507 7108 22508 7172
rect 22572 7108 22573 7172
rect 22507 7107 22573 7108
rect 23062 6901 23122 25875
rect 24715 22948 24781 22949
rect 24715 22884 24716 22948
rect 24780 22884 24781 22948
rect 24715 22883 24781 22884
rect 24718 6901 24778 22883
rect 26923 21996 26989 21997
rect 26923 21932 26924 21996
rect 26988 21932 26989 21996
rect 26923 21931 26989 21932
rect 26371 17780 26437 17781
rect 26371 17716 26372 17780
rect 26436 17716 26437 17780
rect 26371 17715 26437 17716
rect 24899 15740 24965 15741
rect 24899 15676 24900 15740
rect 24964 15676 24965 15740
rect 24899 15675 24965 15676
rect 24902 9077 24962 15675
rect 26187 15060 26253 15061
rect 26187 14996 26188 15060
rect 26252 14996 26253 15060
rect 26187 14995 26253 14996
rect 26003 13972 26069 13973
rect 26003 13908 26004 13972
rect 26068 13970 26069 13972
rect 26190 13970 26250 14995
rect 26374 14245 26434 17715
rect 26371 14244 26437 14245
rect 26371 14180 26372 14244
rect 26436 14180 26437 14244
rect 26371 14179 26437 14180
rect 26068 13910 26250 13970
rect 26068 13908 26069 13910
rect 26003 13907 26069 13908
rect 24899 9076 24965 9077
rect 24899 9012 24900 9076
rect 24964 9012 24965 9076
rect 24899 9011 24965 9012
rect 23059 6900 23125 6901
rect 23059 6836 23060 6900
rect 23124 6836 23125 6900
rect 23059 6835 23125 6836
rect 24715 6900 24781 6901
rect 24715 6836 24716 6900
rect 24780 6836 24781 6900
rect 24715 6835 24781 6836
rect 22323 6764 22389 6765
rect 22323 6700 22324 6764
rect 22388 6700 22389 6764
rect 22323 6699 22389 6700
rect 26926 5541 26986 21931
rect 27107 20228 27173 20229
rect 27107 20164 27108 20228
rect 27172 20164 27173 20228
rect 27107 20163 27173 20164
rect 27110 13837 27170 20163
rect 27294 15061 27354 33083
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 27291 15060 27357 15061
rect 27291 14996 27292 15060
rect 27356 14996 27357 15060
rect 27291 14995 27357 14996
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 27107 13836 27173 13837
rect 27107 13772 27108 13836
rect 27172 13772 27173 13836
rect 27107 13771 27173 13772
rect 27659 13836 27725 13837
rect 27659 13772 27660 13836
rect 27724 13772 27725 13836
rect 27659 13771 27725 13772
rect 27662 5677 27722 13771
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 27659 5676 27725 5677
rect 27659 5612 27660 5676
rect 27724 5612 27725 5676
rect 27659 5611 27725 5612
rect 26923 5540 26989 5541
rect 26923 5476 26924 5540
rect 26988 5476 26989 5540
rect 26923 5475 26989 5476
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 21955 4044 22021 4045
rect 21955 3980 21956 4044
rect 22020 3980 22021 4044
rect 21955 3979 22021 3980
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 21771 2548 21837 2549
rect 21771 2484 21772 2548
rect 21836 2484 21837 2548
rect 21771 2483 21837 2484
rect 21587 2412 21653 2413
rect 21587 2348 21588 2412
rect 21652 2348 21653 2412
rect 21587 2347 21653 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 5027 1324 5093 1325
rect 5027 1260 5028 1324
rect 5092 1260 5093 1324
rect 5027 1259 5093 1260
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 24840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1667941163
transform 1 0 22264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1667941163
transform 1 0 23552 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1667941163
transform 1 0 25484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1667941163
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1667941163
transform 1 0 22264 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1667941163
transform 1 0 30728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1667941163
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1667941163
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1667941163
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1667941163
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1667941163
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1667941163
transform 1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1667941163
transform 1 0 22264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1667941163
transform 1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1667941163
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1667941163
transform 1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1667941163
transform 1 0 2116 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1667941163
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1667941163
transform 1 0 10948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1667941163
transform 1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39
timestamp 1667941163
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1667941163
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1667941163
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_126
timestamp 1667941163
transform 1 0 12696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1667941163
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1667941163
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1667941163
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1667941163
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_231
timestamp 1667941163
transform 1 0 22356 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 1667941163
transform 1 0 23092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1667941163
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1667941163
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1667941163
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_287
timestamp 1667941163
transform 1 0 27508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_295
timestamp 1667941163
transform 1 0 28244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1667941163
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1667941163
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_320
timestamp 1667941163
transform 1 0 30544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_324
timestamp 1667941163
transform 1 0 30912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1667941163
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_343
timestamp 1667941163
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1667941163
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_379
timestamp 1667941163
transform 1 0 35972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_385
timestamp 1667941163
transform 1 0 36524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1667941163
transform 1 0 3404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1667941163
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_71
timestamp 1667941163
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_79
timestamp 1667941163
transform 1 0 8372 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1667941163
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1667941163
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_119
timestamp 1667941163
transform 1 0 12052 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_130
timestamp 1667941163
transform 1 0 13064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1667941163
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1667941163
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1667941163
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1667941163
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1667941163
transform 1 0 17204 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_183
timestamp 1667941163
transform 1 0 17940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1667941163
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1667941163
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_203
timestamp 1667941163
transform 1 0 19780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1667941163
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1667941163
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1667941163
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_252
timestamp 1667941163
transform 1 0 24288 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_262
timestamp 1667941163
transform 1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_266
timestamp 1667941163
transform 1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1667941163
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1667941163
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_289
timestamp 1667941163
transform 1 0 27692 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_345
timestamp 1667941163
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1667941163
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1667941163
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_63
timestamp 1667941163
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_71
timestamp 1667941163
transform 1 0 7636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1667941163
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1667941163
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1667941163
transform 1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1667941163
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1667941163
transform 1 0 11868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1667941163
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_131
timestamp 1667941163
transform 1 0 13156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1667941163
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1667941163
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1667941163
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1667941163
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1667941163
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1667941163
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1667941163
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_190
timestamp 1667941163
transform 1 0 18584 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1667941163
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1667941163
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_216
timestamp 1667941163
transform 1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_223
timestamp 1667941163
transform 1 0 21620 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_228
timestamp 1667941163
transform 1 0 22080 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_232
timestamp 1667941163
transform 1 0 22448 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_237
timestamp 1667941163
transform 1 0 22908 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1667941163
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_258
timestamp 1667941163
transform 1 0 24840 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_270
timestamp 1667941163
transform 1 0 25944 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_282
timestamp 1667941163
transform 1 0 27048 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_294
timestamp 1667941163
transform 1 0 28152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1667941163
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_385
timestamp 1667941163
transform 1 0 36524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_390
timestamp 1667941163
transform 1 0 36984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1667941163
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1667941163
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1667941163
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1667941163
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_63
timestamp 1667941163
transform 1 0 6900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_71
timestamp 1667941163
transform 1 0 7636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1667941163
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_82
timestamp 1667941163
transform 1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1667941163
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1667941163
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1667941163
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1667941163
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1667941163
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1667941163
transform 1 0 13156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1667941163
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1667941163
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1667941163
transform 1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1667941163
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1667941163
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_174
timestamp 1667941163
transform 1 0 17112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1667941163
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1667941163
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1667941163
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_209
timestamp 1667941163
transform 1 0 20332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1667941163
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1667941163
transform 1 0 22264 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1667941163
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1667941163
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_263
timestamp 1667941163
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1667941163
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1667941163
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_33
timestamp 1667941163
transform 1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1667941163
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_43
timestamp 1667941163
transform 1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp 1667941163
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1667941163
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_75
timestamp 1667941163
transform 1 0 8004 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1667941163
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_90
timestamp 1667941163
transform 1 0 9384 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_98
timestamp 1667941163
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1667941163
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1667941163
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1667941163
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1667941163
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_131
timestamp 1667941163
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1667941163
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1667941163
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1667941163
transform 1 0 14812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_156
timestamp 1667941163
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1667941163
transform 1 0 16100 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp 1667941163
transform 1 0 16744 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_184
timestamp 1667941163
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1667941163
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_202
timestamp 1667941163
transform 1 0 19688 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_216
timestamp 1667941163
transform 1 0 20976 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1667941163
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_230
timestamp 1667941163
transform 1 0 22264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1667941163
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1667941163
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_325
timestamp 1667941163
transform 1 0 31004 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_329
timestamp 1667941163
transform 1 0 31372 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_341
timestamp 1667941163
transform 1 0 32476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_353
timestamp 1667941163
transform 1 0 33580 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1667941163
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1667941163
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1667941163
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1667941163
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1667941163
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1667941163
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_99
timestamp 1667941163
transform 1 0 10212 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1667941163
transform 1 0 10580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1667941163
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_124
timestamp 1667941163
transform 1 0 12512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1667941163
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1667941163
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1667941163
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_152
timestamp 1667941163
transform 1 0 15088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_159
timestamp 1667941163
transform 1 0 15732 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1667941163
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_180
timestamp 1667941163
transform 1 0 17664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1667941163
transform 1 0 18308 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1667941163
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_201
timestamp 1667941163
transform 1 0 19596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp 1667941163
transform 1 0 20332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_216
timestamp 1667941163
transform 1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_228
timestamp 1667941163
transform 1 0 22080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_232
timestamp 1667941163
transform 1 0 22448 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_244
timestamp 1667941163
transform 1 0 23552 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_256
timestamp 1667941163
transform 1 0 24656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_268
timestamp 1667941163
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1667941163
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1667941163
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1667941163
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1667941163
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_90
timestamp 1667941163
transform 1 0 9384 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_99
timestamp 1667941163
transform 1 0 10212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_110
timestamp 1667941163
transform 1 0 11224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1667941163
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_124
timestamp 1667941163
transform 1 0 12512 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_134
timestamp 1667941163
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1667941163
transform 1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1667941163
transform 1 0 16100 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_174
timestamp 1667941163
transform 1 0 17112 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_182
timestamp 1667941163
transform 1 0 17848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1667941163
transform 1 0 18308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1667941163
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1667941163
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_212
timestamp 1667941163
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_216
timestamp 1667941163
transform 1 0 20976 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1667941163
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1667941163
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_237
timestamp 1667941163
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1667941163
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_395
timestamp 1667941163
transform 1 0 37444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_399
timestamp 1667941163
transform 1 0 37812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1667941163
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_33
timestamp 1667941163
transform 1 0 4140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_41
timestamp 1667941163
transform 1 0 4876 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_49
timestamp 1667941163
transform 1 0 5612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1667941163
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_70
timestamp 1667941163
transform 1 0 7544 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_96
timestamp 1667941163
transform 1 0 9936 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1667941163
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1667941163
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_135
timestamp 1667941163
transform 1 0 13524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_139
timestamp 1667941163
transform 1 0 13892 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_180
timestamp 1667941163
transform 1 0 17664 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_191
timestamp 1667941163
transform 1 0 18676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_197
timestamp 1667941163
transform 1 0 19228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_201
timestamp 1667941163
transform 1 0 19596 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1667941163
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1667941163
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1667941163
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_228
timestamp 1667941163
transform 1 0 22080 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_232
timestamp 1667941163
transform 1 0 22448 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1667941163
transform 1 0 23368 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_246
timestamp 1667941163
transform 1 0 23736 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_251
timestamp 1667941163
transform 1 0 24196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_263
timestamp 1667941163
transform 1 0 25300 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_275
timestamp 1667941163
transform 1 0 26404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_342
timestamp 1667941163
transform 1 0 32568 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_354
timestamp 1667941163
transform 1 0 33672 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_366
timestamp 1667941163
transform 1 0 34776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_378
timestamp 1667941163
transform 1 0 35880 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1667941163
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1667941163
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1667941163
transform 1 0 6348 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1667941163
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1667941163
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_95
timestamp 1667941163
transform 1 0 9844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_124
timestamp 1667941163
transform 1 0 12512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1667941163
transform 1 0 14720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_158
timestamp 1667941163
transform 1 0 15640 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1667941163
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_181
timestamp 1667941163
transform 1 0 17756 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1667941163
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_202
timestamp 1667941163
transform 1 0 19688 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_216
timestamp 1667941163
transform 1 0 20976 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1667941163
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1667941163
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_237
timestamp 1667941163
transform 1 0 22908 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1667941163
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_258
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_266
timestamp 1667941163
transform 1 0 25576 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_272
timestamp 1667941163
transform 1 0 26128 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_284
timestamp 1667941163
transform 1 0 27232 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_293
timestamp 1667941163
transform 1 0 28060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1667941163
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_349
timestamp 1667941163
transform 1 0 33212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1667941163
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_9
timestamp 1667941163
transform 1 0 1932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_13
timestamp 1667941163
transform 1 0 2300 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1667941163
transform 1 0 4508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_45
timestamp 1667941163
transform 1 0 5244 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1667941163
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_64
timestamp 1667941163
transform 1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_70
timestamp 1667941163
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_94
timestamp 1667941163
transform 1 0 9752 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1667941163
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1667941163
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_159
timestamp 1667941163
transform 1 0 15732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1667941163
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1667941163
transform 1 0 18032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1667941163
transform 1 0 19044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_202
timestamp 1667941163
transform 1 0 19688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1667941163
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1667941163
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_230
timestamp 1667941163
transform 1 0 22264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1667941163
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_251
timestamp 1667941163
transform 1 0 24196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_256
timestamp 1667941163
transform 1 0 24656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_260
timestamp 1667941163
transform 1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_265
timestamp 1667941163
transform 1 0 25484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_277
timestamp 1667941163
transform 1 0 26588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1667941163
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_42
timestamp 1667941163
transform 1 0 4968 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_71
timestamp 1667941163
transform 1 0 7636 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1667941163
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1667941163
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_110
timestamp 1667941163
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1667941163
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1667941163
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1667941163
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1667941163
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_202
timestamp 1667941163
transform 1 0 19688 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_208
timestamp 1667941163
transform 1 0 20240 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_212
timestamp 1667941163
transform 1 0 20608 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1667941163
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1667941163
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_237
timestamp 1667941163
transform 1 0 22908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1667941163
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_268
timestamp 1667941163
transform 1 0 25760 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_275
timestamp 1667941163
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_287
timestamp 1667941163
transform 1 0 27508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1667941163
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_28
timestamp 1667941163
transform 1 0 3680 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1667941163
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_83
timestamp 1667941163
transform 1 0 8740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1667941163
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_138
timestamp 1667941163
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_142
timestamp 1667941163
transform 1 0 14168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1667941163
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_180
timestamp 1667941163
transform 1 0 17664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1667941163
transform 1 0 18032 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_198
timestamp 1667941163
transform 1 0 19320 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_204
timestamp 1667941163
transform 1 0 19872 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_208
timestamp 1667941163
transform 1 0 20240 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_229
timestamp 1667941163
transform 1 0 22172 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_243
timestamp 1667941163
transform 1 0 23460 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_250
timestamp 1667941163
transform 1 0 24104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_257
timestamp 1667941163
transform 1 0 24748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_263
timestamp 1667941163
transform 1 0 25300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_267
timestamp 1667941163
transform 1 0 25668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_272
timestamp 1667941163
transform 1 0 26128 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_301
timestamp 1667941163
transform 1 0 28796 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1667941163
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_54
timestamp 1667941163
transform 1 0 6072 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1667941163
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_96
timestamp 1667941163
transform 1 0 9936 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_102
timestamp 1667941163
transform 1 0 10488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_106
timestamp 1667941163
transform 1 0 10856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_154
timestamp 1667941163
transform 1 0 15272 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_162
timestamp 1667941163
transform 1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1667941163
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1667941163
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1667941163
transform 1 0 20884 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_222
timestamp 1667941163
transform 1 0 21528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_230
timestamp 1667941163
transform 1 0 22264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_241
timestamp 1667941163
transform 1 0 23276 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1667941163
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_258
timestamp 1667941163
transform 1 0 24840 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_264
timestamp 1667941163
transform 1 0 25392 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_268
timestamp 1667941163
transform 1 0 25760 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_280
timestamp 1667941163
transform 1 0 26864 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_296
timestamp 1667941163
transform 1 0 28336 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1667941163
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1667941163
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1667941163
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_86
timestamp 1667941163
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1667941163
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_140
timestamp 1667941163
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1667941163
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1667941163
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1667941163
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1667941163
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_195
timestamp 1667941163
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_211
timestamp 1667941163
transform 1 0 20516 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1667941163
transform 1 0 20884 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1667941163
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_236
timestamp 1667941163
transform 1 0 22816 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_244
timestamp 1667941163
transform 1 0 23552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1667941163
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_269
timestamp 1667941163
transform 1 0 25852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1667941163
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_33
timestamp 1667941163
transform 1 0 4140 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_39
timestamp 1667941163
transform 1 0 4692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_66
timestamp 1667941163
transform 1 0 7176 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_72
timestamp 1667941163
transform 1 0 7728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1667941163
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1667941163
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_114
timestamp 1667941163
transform 1 0 11592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1667941163
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1667941163
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1667941163
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1667941163
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_203
timestamp 1667941163
transform 1 0 19780 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_211
timestamp 1667941163
transform 1 0 20516 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1667941163
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_223
timestamp 1667941163
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1667941163
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_237
timestamp 1667941163
transform 1 0 22908 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1667941163
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1667941163
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_272
timestamp 1667941163
transform 1 0 26128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_280
timestamp 1667941163
transform 1 0 26864 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_294
timestamp 1667941163
transform 1 0 28152 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1667941163
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_341
timestamp 1667941163
transform 1 0 32476 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_347
timestamp 1667941163
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_359
timestamp 1667941163
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1667941163
transform 1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_29
timestamp 1667941163
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1667941163
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_83
timestamp 1667941163
transform 1 0 8740 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1667941163
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1667941163
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1667941163
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1667941163
transform 1 0 18032 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_192
timestamp 1667941163
transform 1 0 18768 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1667941163
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1667941163
transform 1 0 20424 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1667941163
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1667941163
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_251
timestamp 1667941163
transform 1 0 24196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_257
timestamp 1667941163
transform 1 0 24748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_267
timestamp 1667941163
transform 1 0 25668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1667941163
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_286
timestamp 1667941163
transform 1 0 27416 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_298
timestamp 1667941163
transform 1 0 28520 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_310
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_322
timestamp 1667941163
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 1667941163
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1667941163
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_44
timestamp 1667941163
transform 1 0 5152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_71
timestamp 1667941163
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_75
timestamp 1667941163
transform 1 0 8004 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1667941163
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_98
timestamp 1667941163
transform 1 0 10120 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_129
timestamp 1667941163
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1667941163
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_164
timestamp 1667941163
transform 1 0 16192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1667941163
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1667941163
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_202
timestamp 1667941163
transform 1 0 19688 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1667941163
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1667941163
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1667941163
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1667941163
transform 1 0 24840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_272
timestamp 1667941163
transform 1 0 26128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_279
timestamp 1667941163
transform 1 0 26772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_286
timestamp 1667941163
transform 1 0 27416 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_293
timestamp 1667941163
transform 1 0 28060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1667941163
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_25
timestamp 1667941163
transform 1 0 3404 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1667941163
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1667941163
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1667941163
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1667941163
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1667941163
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1667941163
transform 1 0 18032 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1667941163
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_204
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_211
timestamp 1667941163
transform 1 0 20516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1667941163
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_234
timestamp 1667941163
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_244
timestamp 1667941163
transform 1 0 23552 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_250
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_264
timestamp 1667941163
transform 1 0 25392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1667941163
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1667941163
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_299
timestamp 1667941163
transform 1 0 28612 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_303
timestamp 1667941163
transform 1 0 28980 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_315
timestamp 1667941163
transform 1 0 30084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_327
timestamp 1667941163
transform 1 0 31188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_360
timestamp 1667941163
transform 1 0 34224 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_372
timestamp 1667941163
transform 1 0 35328 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_384
timestamp 1667941163
transform 1 0 36432 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1667941163
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_44
timestamp 1667941163
transform 1 0 5152 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1667941163
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1667941163
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1667941163
transform 1 0 10120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1667941163
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1667941163
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_161
timestamp 1667941163
transform 1 0 15916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_169
timestamp 1667941163
transform 1 0 16652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1667941163
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1667941163
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_214
timestamp 1667941163
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_221
timestamp 1667941163
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_227
timestamp 1667941163
transform 1 0 21988 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1667941163
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1667941163
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1667941163
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_266
timestamp 1667941163
transform 1 0 25576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_281
timestamp 1667941163
transform 1 0 26956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_288
timestamp 1667941163
transform 1 0 27600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_300
timestamp 1667941163
transform 1 0 28704 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_327
timestamp 1667941163
transform 1 0 31188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_339
timestamp 1667941163
transform 1 0 32292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_351
timestamp 1667941163
transform 1 0 33396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_370
timestamp 1667941163
transform 1 0 35144 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_382
timestamp 1667941163
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_394
timestamp 1667941163
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_34
timestamp 1667941163
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_83
timestamp 1667941163
transform 1 0 8740 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1667941163
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1667941163
transform 1 0 13892 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1667941163
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1667941163
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_198
timestamp 1667941163
transform 1 0 19320 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_204
timestamp 1667941163
transform 1 0 19872 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1667941163
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_236
timestamp 1667941163
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1667941163
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_250
timestamp 1667941163
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1667941163
transform 1 0 24748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1667941163
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_268
timestamp 1667941163
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1667941163
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1667941163
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_303
timestamp 1667941163
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_315
timestamp 1667941163
transform 1 0 30084 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1667941163
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_342
timestamp 1667941163
transform 1 0 32568 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_354
timestamp 1667941163
transform 1 0 33672 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_366
timestamp 1667941163
transform 1 0 34776 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_378
timestamp 1667941163
transform 1 0 35880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1667941163
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1667941163
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1667941163
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1667941163
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_111
timestamp 1667941163
transform 1 0 11316 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1667941163
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_156
timestamp 1667941163
transform 1 0 15456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1667941163
transform 1 0 17020 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1667941163
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_184
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1667941163
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_214
timestamp 1667941163
transform 1 0 20792 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1667941163
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_235
timestamp 1667941163
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_242
timestamp 1667941163
transform 1 0 23368 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_258
timestamp 1667941163
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_266
timestamp 1667941163
transform 1 0 25576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1667941163
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_290
timestamp 1667941163
transform 1 0 27784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1667941163
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_314
timestamp 1667941163
transform 1 0 29992 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_326
timestamp 1667941163
transform 1 0 31096 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_338
timestamp 1667941163
transform 1 0 32200 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_350
timestamp 1667941163
transform 1 0 33304 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1667941163
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_38
timestamp 1667941163
transform 1 0 4600 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_44
timestamp 1667941163
transform 1 0 5152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1667941163
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_63
timestamp 1667941163
transform 1 0 6900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_67
timestamp 1667941163
transform 1 0 7268 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_91
timestamp 1667941163
transform 1 0 9476 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1667941163
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1667941163
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_142
timestamp 1667941163
transform 1 0 14168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1667941163
transform 1 0 15456 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1667941163
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1667941163
transform 1 0 18308 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1667941163
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1667941163
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_216
timestamp 1667941163
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1667941163
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_236
timestamp 1667941163
transform 1 0 22816 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 1667941163
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_257
timestamp 1667941163
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_271
timestamp 1667941163
transform 1 0 26036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1667941163
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1667941163
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_293
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_301
timestamp 1667941163
transform 1 0 28796 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_311
timestamp 1667941163
transform 1 0 29716 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_319
timestamp 1667941163
transform 1 0 30452 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_324
timestamp 1667941163
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1667941163
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1667941163
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_401
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1667941163
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_54
timestamp 1667941163
transform 1 0 6072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_58
timestamp 1667941163
transform 1 0 6440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1667941163
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1667941163
transform 1 0 9292 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1667941163
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_103
timestamp 1667941163
transform 1 0 10580 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1667941163
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1667941163
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1667941163
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_170
timestamp 1667941163
transform 1 0 16744 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1667941163
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_202
timestamp 1667941163
transform 1 0 19688 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1667941163
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_230
timestamp 1667941163
transform 1 0 22264 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_236
timestamp 1667941163
transform 1 0 22816 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_241
timestamp 1667941163
transform 1 0 23276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1667941163
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1667941163
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_277
timestamp 1667941163
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_284
timestamp 1667941163
transform 1 0 27232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1667941163
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1667941163
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1667941163
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_321
timestamp 1667941163
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_334
timestamp 1667941163
transform 1 0 31832 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_346
timestamp 1667941163
transform 1 0 32936 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1667941163
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1667941163
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_393
timestamp 1667941163
transform 1 0 37260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_397
timestamp 1667941163
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_405
timestamp 1667941163
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 1667941163
transform 1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1667941163
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1667941163
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_62
timestamp 1667941163
transform 1 0 6808 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_91
timestamp 1667941163
transform 1 0 9476 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1667941163
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_148
timestamp 1667941163
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1667941163
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_176
timestamp 1667941163
transform 1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_189
timestamp 1667941163
transform 1 0 18492 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_197
timestamp 1667941163
transform 1 0 19228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1667941163
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1667941163
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1667941163
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_257
timestamp 1667941163
transform 1 0 24748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1667941163
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_271
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1667941163
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_315
timestamp 1667941163
transform 1 0 30084 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_322
timestamp 1667941163
transform 1 0 30728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1667941163
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1667941163
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1667941163
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1667941163
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1667941163
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_402
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1667941163
transform 1 0 38456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1667941163
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_44
timestamp 1667941163
transform 1 0 5152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_69
timestamp 1667941163
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1667941163
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_163
timestamp 1667941163
transform 1 0 16100 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1667941163
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_180
timestamp 1667941163
transform 1 0 17664 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_202
timestamp 1667941163
transform 1 0 19688 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_210
timestamp 1667941163
transform 1 0 20424 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1667941163
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_232
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 1667941163
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1667941163
transform 1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_278
timestamp 1667941163
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_285
timestamp 1667941163
transform 1 0 27324 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_293
timestamp 1667941163
transform 1 0 28060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1667941163
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_328
timestamp 1667941163
transform 1 0 31280 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_340
timestamp 1667941163
transform 1 0 32384 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_352
timestamp 1667941163
transform 1 0 33488 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1667941163
transform 1 0 4784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1667941163
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1667941163
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_67
timestamp 1667941163
transform 1 0 7268 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1667941163
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_98
timestamp 1667941163
transform 1 0 10120 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1667941163
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_138
timestamp 1667941163
transform 1 0 13800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_148
timestamp 1667941163
transform 1 0 14720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_152
timestamp 1667941163
transform 1 0 15088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1667941163
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_184
timestamp 1667941163
transform 1 0 18032 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_190
timestamp 1667941163
transform 1 0 18584 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1667941163
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_214
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1667941163
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1667941163
transform 1 0 23184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1667941163
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1667941163
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_268
timestamp 1667941163
transform 1 0 25760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1667941163
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1667941163
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_286
timestamp 1667941163
transform 1 0 27416 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_292
timestamp 1667941163
transform 1 0 27968 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_306
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_319
timestamp 1667941163
transform 1 0 30452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_326
timestamp 1667941163
transform 1 0 31096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1667941163
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1667941163
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1667941163
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_373
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_377
timestamp 1667941163
transform 1 0 35788 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_381
timestamp 1667941163
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1667941163
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1667941163
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_33
timestamp 1667941163
transform 1 0 4140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_55
timestamp 1667941163
transform 1 0 6164 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1667941163
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_98
timestamp 1667941163
transform 1 0 10120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_102
timestamp 1667941163
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1667941163
transform 1 0 12696 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1667941163
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1667941163
transform 1 0 14720 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1667941163
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1667941163
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_208
timestamp 1667941163
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1667941163
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1667941163
transform 1 0 21252 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_240
timestamp 1667941163
transform 1 0 23184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1667941163
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_268
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_285
timestamp 1667941163
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_292
timestamp 1667941163
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_299
timestamp 1667941163
transform 1 0 28612 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_314
timestamp 1667941163
transform 1 0 29992 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1667941163
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_328
timestamp 1667941163
transform 1 0 31280 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_340
timestamp 1667941163
transform 1 0 32384 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_352
timestamp 1667941163
transform 1 0 33488 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1667941163
transform 1 0 1932 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_36
timestamp 1667941163
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1667941163
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1667941163
transform 1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1667941163
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1667941163
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1667941163
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_152
timestamp 1667941163
transform 1 0 15088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1667941163
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_184
timestamp 1667941163
transform 1 0 18032 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_203
timestamp 1667941163
transform 1 0 19780 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1667941163
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 1667941163
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1667941163
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_251
timestamp 1667941163
transform 1 0 24196 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_255
timestamp 1667941163
transform 1 0 24564 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_265
timestamp 1667941163
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_272
timestamp 1667941163
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_292
timestamp 1667941163
transform 1 0 27968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_299
timestamp 1667941163
transform 1 0 28612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_305
timestamp 1667941163
transform 1 0 29164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1667941163
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_322
timestamp 1667941163
transform 1 0 30728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1667941163
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1667941163
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1667941163
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1667941163
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1667941163
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1667941163
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1667941163
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1667941163
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1667941163
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1667941163
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1667941163
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_126
timestamp 1667941163
transform 1 0 12696 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1667941163
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_156
timestamp 1667941163
transform 1 0 15456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_175
timestamp 1667941163
transform 1 0 17204 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1667941163
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1667941163
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1667941163
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1667941163
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1667941163
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_236
timestamp 1667941163
transform 1 0 22816 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_243
timestamp 1667941163
transform 1 0 23460 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1667941163
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1667941163
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1667941163
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1667941163
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_282
timestamp 1667941163
transform 1 0 27048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_296
timestamp 1667941163
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1667941163
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1667941163
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_327
timestamp 1667941163
transform 1 0 31188 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_334
timestamp 1667941163
transform 1 0 31832 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_346
timestamp 1667941163
transform 1 0 32936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1667941163
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1667941163
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1667941163
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1667941163
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1667941163
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_23
timestamp 1667941163
transform 1 0 3220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1667941163
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1667941163
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_85
timestamp 1667941163
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1667941163
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_134
timestamp 1667941163
transform 1 0 13432 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1667941163
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_184
timestamp 1667941163
transform 1 0 18032 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_192
timestamp 1667941163
transform 1 0 18768 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1667941163
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_209
timestamp 1667941163
transform 1 0 20332 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1667941163
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_230
timestamp 1667941163
transform 1 0 22264 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_238
timestamp 1667941163
transform 1 0 23000 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1667941163
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1667941163
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1667941163
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1667941163
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1667941163
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_297
timestamp 1667941163
transform 1 0 28428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_311
timestamp 1667941163
transform 1 0 29716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_318
timestamp 1667941163
transform 1 0 30360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_325
timestamp 1667941163
transform 1 0 31004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1667941163
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1667941163
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1667941163
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1667941163
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1667941163
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1667941163
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1667941163
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 1667941163
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1667941163
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_58
timestamp 1667941163
transform 1 0 6440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1667941163
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1667941163
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_115
timestamp 1667941163
transform 1 0 11684 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1667941163
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_156
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_166
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1667941163
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1667941163
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1667941163
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1667941163
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1667941163
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_268
timestamp 1667941163
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_275
timestamp 1667941163
transform 1 0 26404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_282
timestamp 1667941163
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1667941163
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1667941163
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_320
timestamp 1667941163
transform 1 0 30544 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1667941163
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_346
timestamp 1667941163
transform 1 0 32936 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1667941163
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1667941163
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1667941163
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_401
timestamp 1667941163
transform 1 0 37996 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1667941163
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1667941163
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1667941163
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_92
timestamp 1667941163
transform 1 0 9568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1667941163
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1667941163
transform 1 0 13248 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1667941163
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_188
timestamp 1667941163
transform 1 0 18400 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_209
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1667941163
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1667941163
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_257
timestamp 1667941163
transform 1 0 24748 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1667941163
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1667941163
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_313
timestamp 1667941163
transform 1 0 29900 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_326
timestamp 1667941163
transform 1 0 31096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1667941163
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1667941163
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1667941163
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1667941163
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1667941163
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1667941163
transform 1 0 37904 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1667941163
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1667941163
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_44
timestamp 1667941163
transform 1 0 5152 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_72
timestamp 1667941163
transform 1 0 7728 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_78
timestamp 1667941163
transform 1 0 8280 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_100
timestamp 1667941163
transform 1 0 10304 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_129
timestamp 1667941163
transform 1 0 12972 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1667941163
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1667941163
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_160
timestamp 1667941163
transform 1 0 15824 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1667941163
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1667941163
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1667941163
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1667941163
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1667941163
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_226
timestamp 1667941163
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_230
timestamp 1667941163
transform 1 0 22264 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_240
timestamp 1667941163
transform 1 0 23184 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_247
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1667941163
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_258
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1667941163
transform 1 0 25944 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_277
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1667941163
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_291
timestamp 1667941163
transform 1 0 27876 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_298
timestamp 1667941163
transform 1 0 28520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1667941163
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_321
timestamp 1667941163
transform 1 0 30636 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_328
timestamp 1667941163
transform 1 0 31280 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_340
timestamp 1667941163
transform 1 0 32384 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_352
timestamp 1667941163
transform 1 0 33488 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1667941163
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_401
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_405
timestamp 1667941163
transform 1 0 38364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_31
timestamp 1667941163
transform 1 0 3956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_63
timestamp 1667941163
transform 1 0 6900 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_67
timestamp 1667941163
transform 1 0 7268 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1667941163
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_92
timestamp 1667941163
transform 1 0 9568 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_138
timestamp 1667941163
transform 1 0 13800 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1667941163
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1667941163
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1667941163
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_203
timestamp 1667941163
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1667941163
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1667941163
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1667941163
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_245
timestamp 1667941163
transform 1 0 23644 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_251
timestamp 1667941163
transform 1 0 24196 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_255
timestamp 1667941163
transform 1 0 24564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_269
timestamp 1667941163
transform 1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1667941163
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_286
timestamp 1667941163
transform 1 0 27416 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_294
timestamp 1667941163
transform 1 0 28152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_299
timestamp 1667941163
transform 1 0 28612 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1667941163
transform 1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_313
timestamp 1667941163
transform 1 0 29900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1667941163
transform 1 0 31004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1667941163
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1667941163
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_25
timestamp 1667941163
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_35
timestamp 1667941163
transform 1 0 4324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1667941163
transform 1 0 6992 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_68
timestamp 1667941163
transform 1 0 7360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1667941163
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_100
timestamp 1667941163
transform 1 0 10304 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_106
timestamp 1667941163
transform 1 0 10856 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_127
timestamp 1667941163
transform 1 0 12788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_156
timestamp 1667941163
transform 1 0 15456 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_164
timestamp 1667941163
transform 1 0 16192 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1667941163
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_185
timestamp 1667941163
transform 1 0 18124 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_212
timestamp 1667941163
transform 1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_220
timestamp 1667941163
transform 1 0 21344 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_225
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1667941163
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1667941163
transform 1 0 25944 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1667941163
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_289
timestamp 1667941163
transform 1 0 27692 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_293
timestamp 1667941163
transform 1 0 28060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1667941163
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_326
timestamp 1667941163
transform 1 0 31096 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_338
timestamp 1667941163
transform 1 0 32200 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_350
timestamp 1667941163
transform 1 0 33304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1667941163
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1667941163
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1667941163
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_40
timestamp 1667941163
transform 1 0 4784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_44
timestamp 1667941163
transform 1 0 5152 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1667941163
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1667941163
transform 1 0 7176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1667941163
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_128
timestamp 1667941163
transform 1 0 12880 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_134
timestamp 1667941163
transform 1 0 13432 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_144
timestamp 1667941163
transform 1 0 14352 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_153
timestamp 1667941163
transform 1 0 15180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1667941163
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1667941163
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1667941163
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1667941163
transform 1 0 18032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_197
timestamp 1667941163
transform 1 0 19228 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_214
timestamp 1667941163
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1667941163
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_230
timestamp 1667941163
transform 1 0 22264 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_239
timestamp 1667941163
transform 1 0 23092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_246
timestamp 1667941163
transform 1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1667941163
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_260
timestamp 1667941163
transform 1 0 25024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_267
timestamp 1667941163
transform 1 0 25668 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_296
timestamp 1667941163
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_309
timestamp 1667941163
transform 1 0 29532 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_316
timestamp 1667941163
transform 1 0 30176 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1667941163
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1667941163
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1667941163
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1667941163
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_52
timestamp 1667941163
transform 1 0 5888 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_76
timestamp 1667941163
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_100
timestamp 1667941163
transform 1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_105
timestamp 1667941163
transform 1 0 10764 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1667941163
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1667941163
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_162
timestamp 1667941163
transform 1 0 16008 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_175
timestamp 1667941163
transform 1 0 17204 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_183
timestamp 1667941163
transform 1 0 17940 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_187
timestamp 1667941163
transform 1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1667941163
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_208
timestamp 1667941163
transform 1 0 20240 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_225
timestamp 1667941163
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_232
timestamp 1667941163
transform 1 0 22448 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_240
timestamp 1667941163
transform 1 0 23184 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_258
timestamp 1667941163
transform 1 0 24840 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_270
timestamp 1667941163
transform 1 0 25944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_278
timestamp 1667941163
transform 1 0 26680 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_283
timestamp 1667941163
transform 1 0 27140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1667941163
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1667941163
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1667941163
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1667941163
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1667941163
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 1667941163
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1667941163
transform 1 0 3680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1667941163
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_68
timestamp 1667941163
transform 1 0 7360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1667941163
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1667941163
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_154
timestamp 1667941163
transform 1 0 15272 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_162
timestamp 1667941163
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1667941163
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_180
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_201
timestamp 1667941163
transform 1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_209
timestamp 1667941163
transform 1 0 20332 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_213
timestamp 1667941163
transform 1 0 20700 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1667941163
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1667941163
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_259
timestamp 1667941163
transform 1 0 24932 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_267
timestamp 1667941163
transform 1 0 25668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1667941163
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_290
timestamp 1667941163
transform 1 0 27784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_295
timestamp 1667941163
transform 1 0 28244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_303
timestamp 1667941163
transform 1 0 28980 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_318
timestamp 1667941163
transform 1 0 30360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_325
timestamp 1667941163
transform 1 0 31004 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1667941163
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1667941163
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1667941163
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1667941163
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1667941163
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1667941163
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_51
timestamp 1667941163
transform 1 0 5796 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1667941163
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_156
timestamp 1667941163
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_163
timestamp 1667941163
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1667941163
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_184
timestamp 1667941163
transform 1 0 18032 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1667941163
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_216
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_224
timestamp 1667941163
transform 1 0 21712 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1667941163
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1667941163
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1667941163
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_268
timestamp 1667941163
transform 1 0 25760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_276
timestamp 1667941163
transform 1 0 26496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_291
timestamp 1667941163
transform 1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1667941163
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_314
timestamp 1667941163
transform 1 0 29992 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_326
timestamp 1667941163
transform 1 0 31096 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_338
timestamp 1667941163
transform 1 0 32200 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_350
timestamp 1667941163
transform 1 0 33304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1667941163
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1667941163
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1667941163
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1667941163
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_28
timestamp 1667941163
transform 1 0 3680 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1667941163
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1667941163
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_77
timestamp 1667941163
transform 1 0 8188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1667941163
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1667941163
transform 1 0 13892 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_156
timestamp 1667941163
transform 1 0 15456 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_162
timestamp 1667941163
transform 1 0 16008 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1667941163
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_187
timestamp 1667941163
transform 1 0 18308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1667941163
transform 1 0 19872 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_208
timestamp 1667941163
transform 1 0 20240 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1667941163
transform 1 0 23184 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1667941163
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1667941163
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_261
timestamp 1667941163
transform 1 0 25116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_268
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_292
timestamp 1667941163
transform 1 0 27968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_296
timestamp 1667941163
transform 1 0 28336 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_306
timestamp 1667941163
transform 1 0 29256 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_313
timestamp 1667941163
transform 1 0 29900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1667941163
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1667941163
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1667941163
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1667941163
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1667941163
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1667941163
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_58
timestamp 1667941163
transform 1 0 6440 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_111
timestamp 1667941163
transform 1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1667941163
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_149
timestamp 1667941163
transform 1 0 14812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1667941163
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_182
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_190
timestamp 1667941163
transform 1 0 18584 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_203
timestamp 1667941163
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_220
timestamp 1667941163
transform 1 0 21344 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1667941163
transform 1 0 22080 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1667941163
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1667941163
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_264
timestamp 1667941163
transform 1 0 25392 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_272
timestamp 1667941163
transform 1 0 26128 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_278
timestamp 1667941163
transform 1 0 26680 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_290
timestamp 1667941163
transform 1 0 27784 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_296
timestamp 1667941163
transform 1 0 28336 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1667941163
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1667941163
transform 1 0 30268 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_324
timestamp 1667941163
transform 1 0 30912 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_336
timestamp 1667941163
transform 1 0 32016 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_348
timestamp 1667941163
transform 1 0 33120 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1667941163
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1667941163
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_389
timestamp 1667941163
transform 1 0 36892 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1667941163
transform 1 0 2852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_31
timestamp 1667941163
transform 1 0 3956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_45
timestamp 1667941163
transform 1 0 5244 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1667941163
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_68
timestamp 1667941163
transform 1 0 7360 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_75
timestamp 1667941163
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_99
timestamp 1667941163
transform 1 0 10212 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_135
timestamp 1667941163
transform 1 0 13524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_152
timestamp 1667941163
transform 1 0 15088 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_156
timestamp 1667941163
transform 1 0 15456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_184
timestamp 1667941163
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_188
timestamp 1667941163
transform 1 0 18400 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_192
timestamp 1667941163
transform 1 0 18768 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_209
timestamp 1667941163
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1667941163
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_230
timestamp 1667941163
transform 1 0 22264 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1667941163
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_254
timestamp 1667941163
transform 1 0 24472 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_267
timestamp 1667941163
transform 1 0 25668 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_273
timestamp 1667941163
transform 1 0 26220 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_277
timestamp 1667941163
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_302
timestamp 1667941163
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_314
timestamp 1667941163
transform 1 0 29992 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_326
timestamp 1667941163
transform 1 0 31096 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1667941163
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1667941163
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_399
timestamp 1667941163
transform 1 0 37812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1667941163
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1667941163
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_36
timestamp 1667941163
transform 1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1667941163
transform 1 0 9476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_105
timestamp 1667941163
transform 1 0 10764 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_131
timestamp 1667941163
transform 1 0 13156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1667941163
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_152
timestamp 1667941163
transform 1 0 15088 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1667941163
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_176
timestamp 1667941163
transform 1 0 17296 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_187
timestamp 1667941163
transform 1 0 18308 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_212
timestamp 1667941163
transform 1 0 20608 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_219
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_236
timestamp 1667941163
transform 1 0 22816 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_244
timestamp 1667941163
transform 1 0 23552 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1667941163
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_265
timestamp 1667941163
transform 1 0 25484 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_271
timestamp 1667941163
transform 1 0 26036 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_281
timestamp 1667941163
transform 1 0 26956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_293
timestamp 1667941163
transform 1 0 28060 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_297
timestamp 1667941163
transform 1 0 28428 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1667941163
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_316
timestamp 1667941163
transform 1 0 30176 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_328
timestamp 1667941163
transform 1 0 31280 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_340
timestamp 1667941163
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1667941163
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1667941163
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_389
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_399
timestamp 1667941163
transform 1 0 37812 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_24
timestamp 1667941163
transform 1 0 3312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_30
timestamp 1667941163
transform 1 0 3864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1667941163
transform 1 0 4784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_53
timestamp 1667941163
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_63
timestamp 1667941163
transform 1 0 6900 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_70
timestamp 1667941163
transform 1 0 7544 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_87
timestamp 1667941163
transform 1 0 9108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_95
timestamp 1667941163
transform 1 0 9844 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1667941163
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_128
timestamp 1667941163
transform 1 0 12880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_135
timestamp 1667941163
transform 1 0 13524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_142
timestamp 1667941163
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_156
timestamp 1667941163
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1667941163
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_174
timestamp 1667941163
transform 1 0 17112 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_183
timestamp 1667941163
transform 1 0 17940 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_190
timestamp 1667941163
transform 1 0 18584 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1667941163
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 1667941163
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_230
timestamp 1667941163
transform 1 0 22264 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_244
timestamp 1667941163
transform 1 0 23552 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_256
timestamp 1667941163
transform 1 0 24656 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_292
timestamp 1667941163
transform 1 0 27968 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_304
timestamp 1667941163
transform 1 0 29072 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_316
timestamp 1667941163
transform 1 0 30176 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_323
timestamp 1667941163
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1667941163
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1667941163
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1667941163
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1667941163
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1667941163
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_9
timestamp 1667941163
transform 1 0 1932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1667941163
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_40
timestamp 1667941163
transform 1 0 4784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_47
timestamp 1667941163
transform 1 0 5428 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_54
timestamp 1667941163
transform 1 0 6072 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_63
timestamp 1667941163
transform 1 0 6900 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_67
timestamp 1667941163
transform 1 0 7268 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1667941163
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_96
timestamp 1667941163
transform 1 0 9936 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_104
timestamp 1667941163
transform 1 0 10672 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_119
timestamp 1667941163
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_127
timestamp 1667941163
transform 1 0 12788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_152
timestamp 1667941163
transform 1 0 15088 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_156
timestamp 1667941163
transform 1 0 15456 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_170
timestamp 1667941163
transform 1 0 16744 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_183
timestamp 1667941163
transform 1 0 17940 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_187
timestamp 1667941163
transform 1 0 18308 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1667941163
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_213
timestamp 1667941163
transform 1 0 20700 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_226
timestamp 1667941163
transform 1 0 21896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_233
timestamp 1667941163
transform 1 0 22540 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1667941163
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_261
timestamp 1667941163
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_266
timestamp 1667941163
transform 1 0 25576 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_278
timestamp 1667941163
transform 1 0 26680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_285
timestamp 1667941163
transform 1 0 27324 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_292
timestamp 1667941163
transform 1 0 27968 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_303
timestamp 1667941163
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1667941163
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1667941163
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1667941163
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1667941163
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_377
timestamp 1667941163
transform 1 0 35788 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_386
timestamp 1667941163
transform 1 0 36616 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_398
timestamp 1667941163
transform 1 0 37720 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_12
timestamp 1667941163
transform 1 0 2208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_19
timestamp 1667941163
transform 1 0 2852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_26
timestamp 1667941163
transform 1 0 3496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_33
timestamp 1667941163
transform 1 0 4140 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1667941163
transform 1 0 4784 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_47
timestamp 1667941163
transform 1 0 5428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1667941163
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_63
timestamp 1667941163
transform 1 0 6900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_70
timestamp 1667941163
transform 1 0 7544 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_85
timestamp 1667941163
transform 1 0 8924 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_98
timestamp 1667941163
transform 1 0 10120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_106
timestamp 1667941163
transform 1 0 10856 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1667941163
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_128
timestamp 1667941163
transform 1 0 12880 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_134
timestamp 1667941163
transform 1 0 13432 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_138
timestamp 1667941163
transform 1 0 13800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_145
timestamp 1667941163
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_152
timestamp 1667941163
transform 1 0 15088 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_174
timestamp 1667941163
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_181
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_188
timestamp 1667941163
transform 1 0 18400 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_207
timestamp 1667941163
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_214
timestamp 1667941163
transform 1 0 20792 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_218
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1667941163
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_246
timestamp 1667941163
transform 1 0 23736 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_258
timestamp 1667941163
transform 1 0 24840 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_266
timestamp 1667941163
transform 1 0 25576 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1667941163
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_300
timestamp 1667941163
transform 1 0 28704 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_313
timestamp 1667941163
transform 1 0 29900 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_324
timestamp 1667941163
transform 1 0 30912 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1667941163
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1667941163
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_401
timestamp 1667941163
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_19
timestamp 1667941163
transform 1 0 2852 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_26
timestamp 1667941163
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_33
timestamp 1667941163
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_37
timestamp 1667941163
transform 1 0 4508 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_44
timestamp 1667941163
transform 1 0 5152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_61
timestamp 1667941163
transform 1 0 6716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_72
timestamp 1667941163
transform 1 0 7728 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_78
timestamp 1667941163
transform 1 0 8280 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_100
timestamp 1667941163
transform 1 0 10304 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_117
timestamp 1667941163
transform 1 0 11868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1667941163
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_131
timestamp 1667941163
transform 1 0 13156 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1667941163
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_158
timestamp 1667941163
transform 1 0 15640 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_175
timestamp 1667941163
transform 1 0 17204 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_182
timestamp 1667941163
transform 1 0 17848 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_190
timestamp 1667941163
transform 1 0 18584 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1667941163
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_202
timestamp 1667941163
transform 1 0 19688 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1667941163
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1667941163
transform 1 0 22080 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1667941163
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1667941163
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_292
timestamp 1667941163
transform 1 0 27968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1667941163
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1667941163
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1667941163
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1667941163
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1667941163
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1667941163
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_389
timestamp 1667941163
transform 1 0 36892 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_9
timestamp 1667941163
transform 1 0 1932 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_20
timestamp 1667941163
transform 1 0 2944 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_34
timestamp 1667941163
transform 1 0 4232 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_41
timestamp 1667941163
transform 1 0 4876 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1667941163
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_76
timestamp 1667941163
transform 1 0 8096 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_83
timestamp 1667941163
transform 1 0 8740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1667941163
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_99
timestamp 1667941163
transform 1 0 10212 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_106
timestamp 1667941163
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_120
timestamp 1667941163
transform 1 0 12144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1667941163
transform 1 0 12788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_144
timestamp 1667941163
transform 1 0 14352 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_152
timestamp 1667941163
transform 1 0 15088 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_156
timestamp 1667941163
transform 1 0 15456 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_162
timestamp 1667941163
transform 1 0 16008 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_174
timestamp 1667941163
transform 1 0 17112 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_181
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_187
timestamp 1667941163
transform 1 0 18308 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_201
timestamp 1667941163
transform 1 0 19596 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_240
timestamp 1667941163
transform 1 0 23184 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_247
timestamp 1667941163
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1667941163
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_261
timestamp 1667941163
transform 1 0 25116 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1667941163
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_286
timestamp 1667941163
transform 1 0 27416 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_298
timestamp 1667941163
transform 1 0 28520 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_310
timestamp 1667941163
transform 1 0 29624 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_322
timestamp 1667941163
transform 1 0 30728 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_334
timestamp 1667941163
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1667941163
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1667941163
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1667941163
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1667941163
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1667941163
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_12
timestamp 1667941163
transform 1 0 2208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_19
timestamp 1667941163
transform 1 0 2852 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1667941163
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_34
timestamp 1667941163
transform 1 0 4232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_48
timestamp 1667941163
transform 1 0 5520 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_57
timestamp 1667941163
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_71
timestamp 1667941163
transform 1 0 7636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_75
timestamp 1667941163
transform 1 0 8004 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1667941163
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_91
timestamp 1667941163
transform 1 0 9476 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_100
timestamp 1667941163
transform 1 0 10304 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_104
timestamp 1667941163
transform 1 0 10672 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_108
timestamp 1667941163
transform 1 0 11040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_117
timestamp 1667941163
transform 1 0 11868 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 1667941163
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_156
timestamp 1667941163
transform 1 0 15456 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_167
timestamp 1667941163
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_174
timestamp 1667941163
transform 1 0 17112 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_181
timestamp 1667941163
transform 1 0 17756 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1667941163
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_202
timestamp 1667941163
transform 1 0 19688 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_206
timestamp 1667941163
transform 1 0 20056 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1667941163
transform 1 0 20424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_217
timestamp 1667941163
transform 1 0 21068 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_225
timestamp 1667941163
transform 1 0 21804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_229
timestamp 1667941163
transform 1 0 22172 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_237
timestamp 1667941163
transform 1 0 22908 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_244
timestamp 1667941163
transform 1 0 23552 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_258
timestamp 1667941163
transform 1 0 24840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_275
timestamp 1667941163
transform 1 0 26404 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_282
timestamp 1667941163
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_338
timestamp 1667941163
transform 1 0 32200 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_350
timestamp 1667941163
transform 1 0 33304 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1667941163
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_7
timestamp 1667941163
transform 1 0 1748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1667941163
transform 1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_18
timestamp 1667941163
transform 1 0 2760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_22
timestamp 1667941163
transform 1 0 3128 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_26
timestamp 1667941163
transform 1 0 3496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_30
timestamp 1667941163
transform 1 0 3864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_34
timestamp 1667941163
transform 1 0 4232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_41
timestamp 1667941163
transform 1 0 4876 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_49
timestamp 1667941163
transform 1 0 5612 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_53
timestamp 1667941163
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_68
timestamp 1667941163
transform 1 0 7360 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_76
timestamp 1667941163
transform 1 0 8096 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_89
timestamp 1667941163
transform 1 0 9292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1667941163
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_117
timestamp 1667941163
transform 1 0 11868 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_121
timestamp 1667941163
transform 1 0 12236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_138
timestamp 1667941163
transform 1 0 13800 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_155
timestamp 1667941163
transform 1 0 15364 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1667941163
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_174
timestamp 1667941163
transform 1 0 17112 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_182
timestamp 1667941163
transform 1 0 17848 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_188
timestamp 1667941163
transform 1 0 18400 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_205
timestamp 1667941163
transform 1 0 19964 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_237
timestamp 1667941163
transform 1 0 22908 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_256
timestamp 1667941163
transform 1 0 24656 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1667941163
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1667941163
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1667941163
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1667941163
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1667941163
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1667941163
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1667941163
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1667941163
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1667941163
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1667941163
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1667941163
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_19
timestamp 1667941163
transform 1 0 2852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_26
timestamp 1667941163
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_40
timestamp 1667941163
transform 1 0 4784 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_47
timestamp 1667941163
transform 1 0 5428 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_54
timestamp 1667941163
transform 1 0 6072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_61
timestamp 1667941163
transform 1 0 6716 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_68
timestamp 1667941163
transform 1 0 7360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_75
timestamp 1667941163
transform 1 0 8004 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1667941163
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_90
timestamp 1667941163
transform 1 0 9384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_114
timestamp 1667941163
transform 1 0 11592 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1667941163
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1667941163
transform 1 0 14444 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_149
timestamp 1667941163
transform 1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_157
timestamp 1667941163
transform 1 0 15548 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_161
timestamp 1667941163
transform 1 0 15916 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_168
timestamp 1667941163
transform 1 0 16560 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_180
timestamp 1667941163
transform 1 0 17664 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_188
timestamp 1667941163
transform 1 0 18400 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1667941163
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_212
timestamp 1667941163
transform 1 0 20608 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_216
timestamp 1667941163
transform 1 0 20976 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_224
timestamp 1667941163
transform 1 0 21712 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_230
timestamp 1667941163
transform 1 0 22264 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_242
timestamp 1667941163
transform 1 0 23368 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_258
timestamp 1667941163
transform 1 0 24840 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_270
timestamp 1667941163
transform 1 0 25944 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_274
timestamp 1667941163
transform 1 0 26312 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_281
timestamp 1667941163
transform 1 0 26956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_293
timestamp 1667941163
transform 1 0 28060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1667941163
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1667941163
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1667941163
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1667941163
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1667941163
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1667941163
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_401
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_9
timestamp 1667941163
transform 1 0 1932 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_20
timestamp 1667941163
transform 1 0 2944 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_34
timestamp 1667941163
transform 1 0 4232 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_42
timestamp 1667941163
transform 1 0 4968 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_46
timestamp 1667941163
transform 1 0 5336 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1667941163
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_63
timestamp 1667941163
transform 1 0 6900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_67
timestamp 1667941163
transform 1 0 7268 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_74
timestamp 1667941163
transform 1 0 7912 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_82
timestamp 1667941163
transform 1 0 8648 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_96
timestamp 1667941163
transform 1 0 9936 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1667941163
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1667941163
transform 1 0 11960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_131
timestamp 1667941163
transform 1 0 13156 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_145
timestamp 1667941163
transform 1 0 14444 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_152
timestamp 1667941163
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_159
timestamp 1667941163
transform 1 0 15732 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_189
timestamp 1667941163
transform 1 0 18492 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1667941163
transform 1 0 19044 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_212
timestamp 1667941163
transform 1 0 20608 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_218
timestamp 1667941163
transform 1 0 21160 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1667941163
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_229
timestamp 1667941163
transform 1 0 22172 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_234
timestamp 1667941163
transform 1 0 22632 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_246
timestamp 1667941163
transform 1 0 23736 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_258
timestamp 1667941163
transform 1 0 24840 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_270
timestamp 1667941163
transform 1 0 25944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1667941163
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1667941163
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1667941163
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1667941163
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1667941163
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1667941163
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1667941163
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_7
timestamp 1667941163
transform 1 0 1748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_12
timestamp 1667941163
transform 1 0 2208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_19
timestamp 1667941163
transform 1 0 2852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1667941163
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_35
timestamp 1667941163
transform 1 0 4324 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_39
timestamp 1667941163
transform 1 0 4692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_46
timestamp 1667941163
transform 1 0 5336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_50
timestamp 1667941163
transform 1 0 5704 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_54
timestamp 1667941163
transform 1 0 6072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_61
timestamp 1667941163
transform 1 0 6716 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_68
timestamp 1667941163
transform 1 0 7360 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_75
timestamp 1667941163
transform 1 0 8004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1667941163
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_90
timestamp 1667941163
transform 1 0 9384 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_105
timestamp 1667941163
transform 1 0 10764 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_110
timestamp 1667941163
transform 1 0 11224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_127
timestamp 1667941163
transform 1 0 12788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_131
timestamp 1667941163
transform 1 0 13156 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1667941163
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_149
timestamp 1667941163
transform 1 0 14812 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_154
timestamp 1667941163
transform 1 0 15272 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_166
timestamp 1667941163
transform 1 0 16376 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_178
timestamp 1667941163
transform 1 0 17480 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1667941163
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_216
timestamp 1667941163
transform 1 0 20976 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_228
timestamp 1667941163
transform 1 0 22080 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1667941163
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1667941163
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1667941163
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1667941163
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1667941163
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1667941163
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1667941163
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1667941163
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_7
timestamp 1667941163
transform 1 0 1748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_11
timestamp 1667941163
transform 1 0 2116 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_18
timestamp 1667941163
transform 1 0 2760 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_22
timestamp 1667941163
transform 1 0 3128 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_26
timestamp 1667941163
transform 1 0 3496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_30
timestamp 1667941163
transform 1 0 3864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_34
timestamp 1667941163
transform 1 0 4232 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1667941163
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1667941163
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1667941163
transform 1 0 11960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_122
timestamp 1667941163
transform 1 0 12328 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_126
timestamp 1667941163
transform 1 0 12696 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_138
timestamp 1667941163
transform 1 0 13800 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_150
timestamp 1667941163
transform 1 0 14904 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1667941163
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_189
timestamp 1667941163
transform 1 0 18492 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_194
timestamp 1667941163
transform 1 0 18952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_201
timestamp 1667941163
transform 1 0 19596 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_209
timestamp 1667941163
transform 1 0 20332 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_213
timestamp 1667941163
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 1667941163
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1667941163
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1667941163
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1667941163
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_9
timestamp 1667941163
transform 1 0 1932 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_16
timestamp 1667941163
transform 1 0 2576 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1667941163
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_34
timestamp 1667941163
transform 1 0 4232 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_46
timestamp 1667941163
transform 1 0 5336 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_58
timestamp 1667941163
transform 1 0 6440 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_70
timestamp 1667941163
transform 1 0 7544 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1667941163
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_115
timestamp 1667941163
transform 1 0 11684 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_119
timestamp 1667941163
transform 1 0 12052 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_131
timestamp 1667941163
transform 1 0 13156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_186
timestamp 1667941163
transform 1 0 18216 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1667941163
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1667941163
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1667941163
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1667941163
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1667941163
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1667941163
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1667941163
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1667941163
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1667941163
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1667941163
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_373
timestamp 1667941163
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_389
timestamp 1667941163
transform 1 0 36892 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_17
timestamp 1667941163
transform 1 0 2668 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_22
timestamp 1667941163
transform 1 0 3128 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_29
timestamp 1667941163
transform 1 0 3772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_41
timestamp 1667941163
transform 1 0 4876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1667941163
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1667941163
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1667941163
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_297
timestamp 1667941163
transform 1 0 28428 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_301
timestamp 1667941163
transform 1 0 28796 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_313
timestamp 1667941163
transform 1 0 29900 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_325
timestamp 1667941163
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1667941163
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_16
timestamp 1667941163
transform 1 0 2576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1667941163
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_61
timestamp 1667941163
transform 1 0 6716 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_66
timestamp 1667941163
transform 1 0 7176 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1667941163
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1667941163
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1667941163
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1667941163
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1667941163
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1667941163
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1667941163
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_314
timestamp 1667941163
transform 1 0 29992 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_326
timestamp 1667941163
transform 1 0 31096 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_338
timestamp 1667941163
transform 1 0 32200 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_350
timestamp 1667941163
transform 1 0 33304 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1667941163
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1667941163
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_8
timestamp 1667941163
transform 1 0 1840 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_246
timestamp 1667941163
transform 1 0 23736 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_258
timestamp 1667941163
transform 1 0 24840 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_270
timestamp 1667941163
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_317
timestamp 1667941163
transform 1 0 30268 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_321
timestamp 1667941163
transform 1 0 30636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1667941163
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1667941163
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1667941163
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1667941163
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_108
timestamp 1667941163
transform 1 0 11040 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_120
timestamp 1667941163
transform 1 0 12144 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1667941163
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_237
timestamp 1667941163
transform 1 0 22908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1667941163
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_258
timestamp 1667941163
transform 1 0 24840 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_270
timestamp 1667941163
transform 1 0 25944 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_282
timestamp 1667941163
transform 1 0 27048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_286
timestamp 1667941163
transform 1 0 27416 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_290
timestamp 1667941163
transform 1 0 27784 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_302
timestamp 1667941163
transform 1 0 28888 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1667941163
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1667941163
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1667941163
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1667941163
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_20
timestamp 1667941163
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_32
timestamp 1667941163
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_44
timestamp 1667941163
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_62
timestamp 1667941163
transform 1 0 6808 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_74
timestamp 1667941163
transform 1 0 7912 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_86
timestamp 1667941163
transform 1 0 9016 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_98
timestamp 1667941163
transform 1 0 10120 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_104
timestamp 1667941163
transform 1 0 10672 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1667941163
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_287
timestamp 1667941163
transform 1 0 27508 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_291
timestamp 1667941163
transform 1 0 27876 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_303
timestamp 1667941163
transform 1 0 28980 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_315
timestamp 1667941163
transform 1 0 30084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_327
timestamp 1667941163
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_369
timestamp 1667941163
transform 1 0 35052 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_376
timestamp 1667941163
transform 1 0 35696 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1667941163
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_103
timestamp 1667941163
transform 1 0 10580 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_107
timestamp 1667941163
transform 1 0 10948 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_119
timestamp 1667941163
transform 1 0 12052 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_131
timestamp 1667941163
transform 1 0 13156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_118
timestamp 1667941163
transform 1 0 11960 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_130
timestamp 1667941163
transform 1 0 13064 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_142
timestamp 1667941163
transform 1 0 14168 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_154
timestamp 1667941163
transform 1 0 15272 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1667941163
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_9
timestamp 1667941163
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_16
timestamp 1667941163
transform 1 0 2576 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_45
timestamp 1667941163
transform 1 0 5244 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_49
timestamp 1667941163
transform 1 0 5612 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_61
timestamp 1667941163
transform 1 0 6716 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_73
timestamp 1667941163
transform 1 0 7820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 1667941163
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_90
timestamp 1667941163
transform 1 0 9384 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_102
timestamp 1667941163
transform 1 0 10488 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_114
timestamp 1667941163
transform 1 0 11592 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_126
timestamp 1667941163
transform 1 0 12696 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1667941163
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_229
timestamp 1667941163
transform 1 0 22172 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_234
timestamp 1667941163
transform 1 0 22632 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1667941163
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_384
timestamp 1667941163
transform 1 0 36432 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_392
timestamp 1667941163
transform 1 0 37168 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_9
timestamp 1667941163
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_17
timestamp 1667941163
transform 1 0 2668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_25
timestamp 1667941163
transform 1 0 3404 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_35
timestamp 1667941163
transform 1 0 4324 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_43
timestamp 1667941163
transform 1 0 5060 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 1667941163
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_62
timestamp 1667941163
transform 1 0 6808 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_74
timestamp 1667941163
transform 1 0 7912 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_86
timestamp 1667941163
transform 1 0 9016 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_97
timestamp 1667941163
transform 1 0 10028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1667941163
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_119
timestamp 1667941163
transform 1 0 12052 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_131
timestamp 1667941163
transform 1 0 13156 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_143
timestamp 1667941163
transform 1 0 14260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_155
timestamp 1667941163
transform 1 0 15364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_177
timestamp 1667941163
transform 1 0 17388 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_183
timestamp 1667941163
transform 1 0 17940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_190
timestamp 1667941163
transform 1 0 18584 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_198
timestamp 1667941163
transform 1 0 19320 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_203
timestamp 1667941163
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1667941163
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_231
timestamp 1667941163
transform 1 0 22356 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_239
timestamp 1667941163
transform 1 0 23092 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_245
timestamp 1667941163
transform 1 0 23644 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_257
timestamp 1667941163
transform 1 0 24748 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_265
timestamp 1667941163
transform 1 0 25484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_269
timestamp 1667941163
transform 1 0 25852 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1667941163
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_289
timestamp 1667941163
transform 1 0 27692 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_294
timestamp 1667941163
transform 1 0 28152 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_302
timestamp 1667941163
transform 1 0 28888 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_307
timestamp 1667941163
transform 1 0 29348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_319
timestamp 1667941163
transform 1 0 30452 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_325
timestamp 1667941163
transform 1 0 31004 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_333
timestamp 1667941163
transform 1 0 31740 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1667941163
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_373
timestamp 1667941163
transform 1 0 35420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_377
timestamp 1667941163
transform 1 0 35788 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_382
timestamp 1667941163
transform 1 0 36248 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_13
timestamp 1667941163
transform 1 0 2300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1667941163
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1667941163
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_34
timestamp 1667941163
transform 1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_42
timestamp 1667941163
transform 1 0 4968 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_54
timestamp 1667941163
transform 1 0 6072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_63
timestamp 1667941163
transform 1 0 6900 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_70
timestamp 1667941163
transform 1 0 7544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_91
timestamp 1667941163
transform 1 0 9476 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_99
timestamp 1667941163
transform 1 0 10212 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1667941163
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_119
timestamp 1667941163
transform 1 0 12052 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_127
timestamp 1667941163
transform 1 0 12788 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1667941163
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1667941163
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_146
timestamp 1667941163
transform 1 0 14536 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_160
timestamp 1667941163
transform 1 0 15824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_188
timestamp 1667941163
transform 1 0 18400 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_203
timestamp 1667941163
transform 1 0 19780 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_208
timestamp 1667941163
transform 1 0 20240 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_233
timestamp 1667941163
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1667941163
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_259
timestamp 1667941163
transform 1 0 24932 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_267
timestamp 1667941163
transform 1 0 25668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1667941163
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_295
timestamp 1667941163
transform 1 0 28244 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_302
timestamp 1667941163
transform 1 0 28888 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_315
timestamp 1667941163
transform 1 0 30084 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_323
timestamp 1667941163
transform 1 0 30820 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_359
timestamp 1667941163
transform 1 0 34132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_399
timestamp 1667941163
transform 1 0 37812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0493_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 23736 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 19596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 28244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 26404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 27692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 18400 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 27140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 26956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 28336 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 21620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 30728 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 29716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 26772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 28244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 23920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 25944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 20608 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 13892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 21252 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 22632 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 23920 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 20056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 21620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 15180 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 28336 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 23736 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 5152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 6624 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 11684 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 11592 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 6808 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 23276 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 22908 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 7268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 19412 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 14168 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 6900 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 8464 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 23184 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 8372 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 18032 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 10764 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 10948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 16192 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 20240 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 27784 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 26312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 23552 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 8280 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 21160 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 18308 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 13524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 16100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 23552 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 25484 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 22632 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 23276 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 25760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 20608 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 23276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 1840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 21988 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 22632 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 25484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 25300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 22172 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 22632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 27600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 25760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 23552 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 24564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 21528 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1667941163
transform 1 0 30084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 6624 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 17020 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 10580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 9936 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 4140 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 5152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 8372 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 8372 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1667941163
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 5796 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 7452 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 18124 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 10304 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 24932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 28704 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 28980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 27784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 14536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 17664 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 16008 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 29624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 16100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 20056 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 22264 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 21160 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 24840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 17940 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 6532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 2576 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 4508 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 20976 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1667941163
transform 1 0 23736 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1667941163
transform 1 0 15640 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 19412 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1667941163
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 26128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 23276 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 20976 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 26312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 28704 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 28060 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 18676 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 26128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1667941163
transform 1 0 24104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 26404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 23368 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 30360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 30452 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 31372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 1932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 6992 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 2576 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 2576 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 3220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 3220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 9752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 5244 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 3220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 1840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 20792 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 18676 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 4600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 3220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 3864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 22540 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 25576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 3956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 4600 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 9292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 14536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 12512 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 20884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1667941163
transform 1 0 7728 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1667941163
transform 1 0 24196 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 17480 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 25392 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 27140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 25024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1667941163
transform 1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 19320 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 25208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 26128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1667941163
transform 1 0 27784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 24748 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 28336 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 31464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 22172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 21988 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 27784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1667941163
transform 1 0 31096 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 15456 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 21988 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 19320 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 13524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 18676 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 18676 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 17480 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 26312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 23552 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 22632 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 16100 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1667941163
transform 1 0 18492 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 20424 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 22448 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 18032 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 2668 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 19412 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 14168 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 25116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 6532 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 10672 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1667941163
transform 1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0803_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34684 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 23276 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 33948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 28520 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 6440 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 30636 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 30544 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0813_
timestamp 1667941163
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 6900 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 30728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 16836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 32660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 28520 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 28704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1667941163
transform 1 0 26404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 26036 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 32752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 9384 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 22908 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 29992 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 29716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 10948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 24288 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 31004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 23828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 2576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 10764 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 9108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1667941163
transform 1 0 17480 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1667941163
transform 1 0 19412 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1667941163
transform 1 0 30360 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0847_
timestamp 1667941163
transform 1 0 5060 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1667941163
transform 1 0 23828 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1667941163
transform 1 0 1932 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0850_
timestamp 1667941163
transform 1 0 11868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1667941163
transform 1 0 10948 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1667941163
transform 1 0 21988 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1667941163
transform 1 0 29900 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1667941163
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1667941163
transform 1 0 32936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1667941163
transform 1 0 22816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1667941163
transform 1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1667941163
transform 1 0 14996 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1667941163
transform 1 0 21896 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1667941163
transform 1 0 26864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1667941163
transform 1 0 27048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1667941163
transform 1 0 17940 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1667941163
transform 1 0 2300 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1667941163
transform 1 0 32292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1667941163
transform 1 0 23184 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1667941163
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1667941163
transform 1 0 23276 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1667941163
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0872_
timestamp 1667941163
transform 1 0 5244 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1667941163
transform 1 0 21988 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1667941163
transform 1 0 10488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1667941163
transform 1 0 31556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1667941163
transform 1 0 20516 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1667941163
transform 1 0 27784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1667941163
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1667941163
transform 1 0 22632 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1667941163
transform 1 0 5704 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1667941163
transform 1 0 20700 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1667941163
transform 1 0 3312 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1667941163
transform 1 0 3956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1667941163
transform 1 0 26128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1667941163
transform 1 0 32292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1667941163
transform 1 0 13248 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1667941163
transform 1 0 27416 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1667941163
transform 1 0 7728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1667941163
transform 1 0 30636 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1667941163
transform 1 0 27784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1667941163
transform 1 0 31924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1667941163
transform 1 0 5796 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1667941163
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1667941163
transform 1 0 26772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1667941163
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1667941163
transform 1 0 24472 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1667941163
transform 1 0 18676 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1667941163
transform 1 0 31464 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1667941163
transform 1 0 24380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1667941163
transform 1 0 25116 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1667941163
transform 1 0 31004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1667941163
transform 1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1667941163
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0906_
timestamp 1667941163
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1667941163
transform 1 0 3956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1667941163
transform 1 0 22632 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0909_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 15548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0910_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0911_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 13156 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1667941163
transform 1 0 15640 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1667941163
transform 1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1667941163
transform 1 0 18400 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1667941163
transform 1 0 18032 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1667941163
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1667941163
transform 1 0 28612 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1667941163
transform 1 0 19872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1667941163
transform 1 0 28796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1667941163
transform 1 0 16468 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1667941163
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0922_
timestamp 1667941163
transform 1 0 14168 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1667941163
transform 1 0 27324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1667941163
transform 1 0 15364 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0925_
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1667941163
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1667941163
transform 1 0 18032 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1667941163
transform 1 0 17572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1667941163
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0931_
timestamp 1667941163
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1667941163
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0933_
timestamp 1667941163
transform 1 0 14168 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1667941163
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1667941163
transform 1 0 24472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1667941163
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0937_
timestamp 1667941163
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1667941163
transform 1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1667941163
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1667941163
transform 1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1667941163
transform 1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0944_
timestamp 1667941163
transform 1 0 12880 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1667941163
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1667941163
transform 1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1667941163
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1667941163
transform 1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp 1667941163
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp 1667941163
transform 1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1667941163
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1667941163
transform 1 0 14720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0955_
timestamp 1667941163
transform 1 0 13064 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1667941163
transform 1 0 3220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1667941163
transform 1 0 3220 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1667941163
transform 1 0 3956 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1667941163
transform 1 0 7636 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1667941163
transform 1 0 12328 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp 1667941163
transform 1 0 15732 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1667941163
transform 1 0 10580 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1667941163
transform 1 0 2668 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp 1667941163
transform 1 0 3312 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0966_
timestamp 1667941163
transform 1 0 13064 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1667941163
transform 1 0 3956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1667941163
transform 1 0 5152 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1667941163
transform 1 0 5796 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1667941163
transform 1 0 4508 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1667941163
transform 1 0 4600 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1667941163
transform 1 0 15824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp 1667941163
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1667941163
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1667941163
transform 1 0 15180 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0977_
timestamp 1667941163
transform 1 0 8096 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1667941163
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1667941163
transform 1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp 1667941163
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1667941163
transform 1 0 18032 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1667941163
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1667941163
transform 1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1667941163
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1667941163
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1667941163
transform 1 0 12788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0988_
timestamp 1667941163
transform 1 0 15824 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1667941163
transform 1 0 27784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1667941163
transform 1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1667941163
transform 1 0 26956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp 1667941163
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1667941163
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1667941163
transform 1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1667941163
transform 1 0 27600 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1667941163
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0999_
timestamp 1667941163
transform 1 0 14444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1667941163
transform 1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1667941163
transform 1 0 6440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1667941163
transform 1 0 7728 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1667941163
transform 1 0 6072 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1667941163
transform 1 0 10948 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1667941163
transform 1 0 15640 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1667941163
transform 1 0 22632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1667941163
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1010_
timestamp 1667941163
transform 1 0 15088 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp 1667941163
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp 1667941163
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1667941163
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1667941163
transform 1 0 14260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1667941163
transform 1 0 9108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1667941163
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1667941163
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1667941163
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1667941163
transform 1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1021_
timestamp 1667941163
transform 1 0 19412 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1667941163
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1667941163
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1667941163
transform 1 0 28336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1667941163
transform 1 0 28980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1667941163
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1667941163
transform 1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1667941163
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1667941163
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1032_
timestamp 1667941163
transform 1 0 15824 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1667941163
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1667941163
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1667941163
transform 1 0 14168 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1667941163
transform 1 0 26036 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1667941163
transform 1 0 27140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1667941163
transform 1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1043_
timestamp 1667941163
transform 1 0 18492 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1667941163
transform 1 0 18124 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1667941163
transform 1 0 15824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1667941163
transform 1 0 18676 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1667941163
transform 1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1667941163
transform 1 0 14536 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1667941163
transform 1 0 13248 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1667941163
transform 1 0 17112 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1667941163
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1054_
timestamp 1667941163
transform 1 0 15824 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1667941163
transform 1 0 15364 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1667941163
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1667941163
transform 1 0 26496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1667941163
transform 1 0 14444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1667941163
transform 1 0 29808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1667941163
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1667941163
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1667941163
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1667941163
transform 1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1667941163
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1065_
timestamp 1667941163
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1667941163
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1667941163
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1667941163
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1667941163
transform 1 0 11592 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1667941163
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1667941163
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1667941163
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1667941163
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1667941163
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1667941163
transform 1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1667941163
transform 1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1078_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1656 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1079_
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1080_
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1081_
timestamp 1667941163
transform 1 0 1748 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1082_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 11684 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1083_
timestamp 1667941163
transform 1 0 10580 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1084_
timestamp 1667941163
transform 1 0 7544 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1085_
timestamp 1667941163
transform 1 0 6532 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1086_
timestamp 1667941163
transform 1 0 1656 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1087_
timestamp 1667941163
transform 1 0 1656 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1088_
timestamp 1667941163
transform 1 0 4232 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1089_
timestamp 1667941163
transform 1 0 1656 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1090_
timestamp 1667941163
transform 1 0 6532 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1091_
timestamp 1667941163
transform 1 0 6440 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1092_
timestamp 1667941163
transform 1 0 3956 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1093_
timestamp 1667941163
transform 1 0 3956 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1094_
timestamp 1667941163
transform 1 0 6716 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1095_
timestamp 1667941163
transform 1 0 6256 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1096_
timestamp 1667941163
transform 1 0 4232 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1097_
timestamp 1667941163
transform 1 0 4508 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1098_
timestamp 1667941163
transform 1 0 5520 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1099_
timestamp 1667941163
transform 1 0 3956 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1100_
timestamp 1667941163
transform 1 0 1564 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1101_
timestamp 1667941163
transform 1 0 2392 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1667941163
transform 1 0 11868 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1667941163
transform 1 0 9292 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1667941163
transform 1 0 6624 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1106_
timestamp 1667941163
transform 1 0 11776 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1107_
timestamp 1667941163
transform 1 0 11684 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1108_
timestamp 1667941163
transform 1 0 11868 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1109_
timestamp 1667941163
transform 1 0 11684 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1667941163
transform 1 0 11684 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1667941163
transform 1 0 9384 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1667941163
transform 1 0 6900 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1667941163
transform 1 0 13892 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1114_
timestamp 1667941163
transform 1 0 9108 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1115_
timestamp 1667941163
transform 1 0 11224 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1116_
timestamp 1667941163
transform 1 0 6532 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1117_
timestamp 1667941163
transform 1 0 3956 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1667941163
transform 1 0 1564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1122_
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1123_
timestamp 1667941163
transform 1 0 2300 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1124_
timestamp 1667941163
transform 1 0 7728 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1125_
timestamp 1667941163
transform 1 0 11868 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1667941163
transform 1 0 4140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1667941163
transform 1 0 5888 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1667941163
transform 1 0 4048 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1129_
timestamp 1667941163
transform 1 0 3956 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1130_
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1131_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2852 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1132_
timestamp 1667941163
transform 1 0 1564 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1133_
timestamp 1667941163
transform 1 0 1840 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1667941163
transform 1 0 11316 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1667941163
transform 1 0 9292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1667941163
transform 1 0 9476 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1667941163
transform 1 0 11684 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1138_
timestamp 1667941163
transform 1 0 11684 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1139_
timestamp 1667941163
transform 1 0 9200 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1667941163
transform 1 0 5704 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1141_
timestamp 1667941163
transform 1 0 5336 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1667941163
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1143_
timestamp 1667941163
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1145_
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1146_
timestamp 1667941163
transform 1 0 2024 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1147_
timestamp 1667941163
transform 1 0 11592 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1148_
timestamp 1667941163
transform 1 0 11224 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1149_
timestamp 1667941163
transform 1 0 10856 0 1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1150_
timestamp 1667941163
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1667941163
transform 1 0 9844 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1667941163
transform 1 0 10948 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1667941163
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1154_
timestamp 1667941163
transform 1 0 10672 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1155_
timestamp 1667941163
transform 1 0 10580 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1156_
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1157_
timestamp 1667941163
transform 1 0 1564 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1667941163
transform 1 0 4600 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1667941163
transform 1 0 1564 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1667941163
transform 1 0 1840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1667941163
transform 1 0 1656 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1162_
timestamp 1667941163
transform 1 0 3956 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1163_
timestamp 1667941163
transform 1 0 3956 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1164_
timestamp 1667941163
transform 1 0 6532 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1165_
timestamp 1667941163
transform 1 0 6808 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1667941163
transform 1 0 4324 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1667941163
transform 1 0 5520 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1667941163
transform 1 0 6532 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1667941163
transform 1 0 1656 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1170_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1171_
timestamp 1667941163
transform 1 0 7636 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1172_
timestamp 1667941163
transform 1 0 8832 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1173_
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1667941163
transform 1 0 3772 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1667941163
transform 1 0 3956 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1667941163
transform 1 0 3680 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1178_
timestamp 1667941163
transform 1 0 6624 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1179_
timestamp 1667941163
transform 1 0 3956 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1180_
timestamp 1667941163
transform 1 0 5060 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1181_
timestamp 1667941163
transform 1 0 10396 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1667941163
transform 1 0 1564 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1667941163
transform 1 0 1656 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1667941163
transform 1 0 1656 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1667941163
transform 1 0 6532 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1186_
timestamp 1667941163
transform 1 0 11868 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1187_
timestamp 1667941163
transform 1 0 11684 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1188_
timestamp 1667941163
transform 1 0 7360 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1189_
timestamp 1667941163
transform 1 0 1564 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1667941163
transform 1 0 7360 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1667941163
transform 1 0 6256 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1667941163
transform 1 0 4324 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1667941163
transform 1 0 4048 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1194_
timestamp 1667941163
transform 1 0 4048 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1195_
timestamp 1667941163
transform 1 0 6624 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1196_
timestamp 1667941163
transform 1 0 2116 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1197_
timestamp 1667941163
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1667941163
transform 1 0 8372 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1199_
timestamp 1667941163
transform 1 0 4232 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1667941163
transform 1 0 6348 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1667941163
transform 1 0 6808 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1202_
timestamp 1667941163
transform 1 0 11316 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1203_
timestamp 1667941163
transform 1 0 11776 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1204_
timestamp 1667941163
transform 1 0 11684 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1205_
timestamp 1667941163
transform 1 0 11684 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1667941163
transform 1 0 1656 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1208_
timestamp 1667941163
transform 1 0 2024 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1209_
timestamp 1667941163
transform 1 0 9108 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1210_
timestamp 1667941163
transform 1 0 7360 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1211_
timestamp 1667941163
transform 1 0 6532 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1667941163
transform 1 0 11500 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1667941163
transform 1 0 6716 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1667941163
transform 1 0 9384 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1215_
timestamp 1667941163
transform 1 0 11684 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1216_
timestamp 1667941163
transform 1 0 9108 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1217_
timestamp 1667941163
transform 1 0 9108 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1667941163
transform 1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1667941163
transform 1 0 8096 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1667941163
transform 1 0 11684 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1221_
timestamp 1667941163
transform 1 0 9108 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1222_
timestamp 1667941163
transform 1 0 10856 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1223_
timestamp 1667941163
transform 1 0 7636 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1224_
timestamp 1667941163
transform 1 0 14260 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1667941163
transform 1 0 14260 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1226_
timestamp 1667941163
transform 1 0 4232 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1227_
timestamp 1667941163
transform 1 0 5520 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1228_
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1229_
timestamp 1667941163
transform 1 0 2668 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_2  _1250_
timestamp 1667941163
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1251_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9752 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1667941163
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1254_
timestamp 1667941163
transform 1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1667941163
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1667941163
transform 1 0 9108 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1257_
timestamp 1667941163
transform 1 0 28336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1667941163
transform 1 0 31096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1667941163
transform 1 0 25576 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1260_
timestamp 1667941163
transform 1 0 23460 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1261_
timestamp 1667941163
transform 1 0 36340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1667941163
transform 1 0 29624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1263_
timestamp 1667941163
transform 1 0 30912 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1264_
timestamp 1667941163
transform 1 0 5336 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1667941163
transform 1 0 2944 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1266_
timestamp 1667941163
transform 1 0 6992 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1267_
timestamp 1667941163
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1268_
timestamp 1667941163
transform 1 0 1656 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1269_
timestamp 1667941163
transform 1 0 27876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1667941163
transform 1 0 17664 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1667941163
transform 1 0 27508 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1272_
timestamp 1667941163
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1273_
timestamp 1667941163
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1274_
timestamp 1667941163
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1667941163
transform 1 0 35512 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1276_
timestamp 1667941163
transform 1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1277_
timestamp 1667941163
transform 1 0 22908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1278_
timestamp 1667941163
transform 1 0 6716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1667941163
transform 1 0 4968 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1280_
timestamp 1667941163
transform 1 0 37444 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1667941163
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1282_
timestamp 1667941163
transform 1 0 27876 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1667941163
transform 1 0 5060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1667941163
transform 1 0 21804 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1667941163
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1286_
timestamp 1667941163
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1667941163
transform 1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1288_
timestamp 1667941163
transform 1 0 23184 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1289_
timestamp 1667941163
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1290_
timestamp 1667941163
transform 1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1291_
timestamp 1667941163
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1292_
timestamp 1667941163
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1293_
timestamp 1667941163
transform 1 0 22356 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1667941163
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1295_
timestamp 1667941163
transform 1 0 29900 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1667941163
transform 1 0 2944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1297_
timestamp 1667941163
transform 1 0 37352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1667941163
transform 1 0 11684 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1667941163
transform 1 0 35880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1300_
timestamp 1667941163
transform 1 0 37812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1301_
timestamp 1667941163
transform 1 0 26312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1667941163
transform 1 0 27600 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1303_
timestamp 1667941163
transform 1 0 16100 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1304_
timestamp 1667941163
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1667941163
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1306_
timestamp 1667941163
transform 1 0 2300 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1307_
timestamp 1667941163
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1308_
timestamp 1667941163
transform 1 0 1840 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1309_
timestamp 1667941163
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1310_
timestamp 1667941163
transform 1 0 21712 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1311_
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1312_
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1313_
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1314_
timestamp 1667941163
transform 1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1315_
timestamp 1667941163
transform 1 0 30728 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1316_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1318_
timestamp 1667941163
transform 1 0 20424 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1319_
timestamp 1667941163
transform 1 0 23092 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1320_
timestamp 1667941163
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1321_
timestamp 1667941163
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1322_
timestamp 1667941163
transform 1 0 3220 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1667941163
transform 1 0 20148 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1324_
timestamp 1667941163
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1325_
timestamp 1667941163
transform 1 0 23920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1326_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1327_
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1328__172 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1328_
timestamp 1667941163
transform 1 0 1656 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1329_
timestamp 1667941163
transform 1 0 20148 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1330_
timestamp 1667941163
transform 1 0 16928 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1331_
timestamp 1667941163
transform 1 0 15180 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1332_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 16192 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1333_
timestamp 1667941163
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1334_
timestamp 1667941163
transform 1 0 19320 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1335_
timestamp 1667941163
transform 1 0 18400 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1336_
timestamp 1667941163
transform 1 0 21804 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1337_
timestamp 1667941163
transform 1 0 20332 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1338_
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1339_
timestamp 1667941163
transform 1 0 18952 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1340_
timestamp 1667941163
transform 1 0 14352 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1341_
timestamp 1667941163
transform 1 0 13156 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1342_
timestamp 1667941163
transform 1 0 13616 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1343_
timestamp 1667941163
transform 1 0 14260 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1344_
timestamp 1667941163
transform 1 0 14904 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1344__173
timestamp 1667941163
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1345_
timestamp 1667941163
transform 1 0 14536 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1346_
timestamp 1667941163
transform 1 0 14812 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1347_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1348_
timestamp 1667941163
transform 1 0 18124 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1349_
timestamp 1667941163
transform 1 0 16836 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1350_
timestamp 1667941163
transform 1 0 21988 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1351_
timestamp 1667941163
transform 1 0 14260 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1352_
timestamp 1667941163
transform 1 0 19780 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1353_
timestamp 1667941163
transform 1 0 22632 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1354_
timestamp 1667941163
transform 1 0 14076 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1355_
timestamp 1667941163
transform 1 0 20056 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1356_
timestamp 1667941163
transform 1 0 23092 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1357_
timestamp 1667941163
transform 1 0 13248 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1358_
timestamp 1667941163
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1359_
timestamp 1667941163
transform 1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1360_
timestamp 1667941163
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1360__174
timestamp 1667941163
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1361_
timestamp 1667941163
transform 1 0 5520 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1362_
timestamp 1667941163
transform 1 0 16836 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1363_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1364_
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1365_
timestamp 1667941163
transform 1 0 19412 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1366_
timestamp 1667941163
transform 1 0 9568 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1367_
timestamp 1667941163
transform 1 0 17940 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1368_
timestamp 1667941163
transform 1 0 17940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1369_
timestamp 1667941163
transform 1 0 16836 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1370_
timestamp 1667941163
transform 1 0 15364 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1371_
timestamp 1667941163
transform 1 0 7912 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1372_
timestamp 1667941163
transform 1 0 15548 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1373_
timestamp 1667941163
transform 1 0 23276 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1374_
timestamp 1667941163
transform 1 0 31096 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1375_
timestamp 1667941163
transform 1 0 28704 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1376_
timestamp 1667941163
transform 1 0 27508 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1376__175
timestamp 1667941163
transform 1 0 27692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1377_
timestamp 1667941163
transform 1 0 22356 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1378_
timestamp 1667941163
transform 1 0 29256 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1379_
timestamp 1667941163
transform 1 0 28704 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1380_
timestamp 1667941163
transform 1 0 28244 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1381_
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1382_
timestamp 1667941163
transform 1 0 28428 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1383_
timestamp 1667941163
transform 1 0 26128 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1384_
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1385_
timestamp 1667941163
transform 1 0 23092 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1386_
timestamp 1667941163
transform 1 0 21344 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1387_
timestamp 1667941163
transform 1 0 25116 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1388_
timestamp 1667941163
transform 1 0 29808 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1389_
timestamp 1667941163
transform 1 0 18124 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1390_
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1391_
timestamp 1667941163
transform 1 0 20056 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1392_
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1392__176
timestamp 1667941163
transform 1 0 30912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1393_
timestamp 1667941163
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1394_
timestamp 1667941163
transform 1 0 19780 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1395_
timestamp 1667941163
transform 1 0 20056 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1396_
timestamp 1667941163
transform 1 0 21252 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1397_
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1398_
timestamp 1667941163
transform 1 0 21528 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1399_
timestamp 1667941163
transform 1 0 24196 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1400_
timestamp 1667941163
transform 1 0 16192 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1401_
timestamp 1667941163
transform 1 0 27140 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1402_
timestamp 1667941163
transform 1 0 22080 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1403_
timestamp 1667941163
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1404_
timestamp 1667941163
transform 1 0 26680 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1405_
timestamp 1667941163
transform 1 0 15180 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1406_
timestamp 1667941163
transform 1 0 11684 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1407_
timestamp 1667941163
transform 1 0 11684 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1408__177
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1408_
timestamp 1667941163
transform 1 0 6900 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1409_
timestamp 1667941163
transform 1 0 20700 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1410_
timestamp 1667941163
transform 1 0 12972 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1411_
timestamp 1667941163
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1412_
timestamp 1667941163
transform 1 0 20332 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1413_
timestamp 1667941163
transform 1 0 16652 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1414_
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1415_
timestamp 1667941163
transform 1 0 3956 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1416_
timestamp 1667941163
transform 1 0 18584 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1417_
timestamp 1667941163
transform 1 0 19412 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1418_
timestamp 1667941163
transform 1 0 9108 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1419_
timestamp 1667941163
transform 1 0 21068 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1420_
timestamp 1667941163
transform 1 0 23460 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1421_
timestamp 1667941163
transform 1 0 17204 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1422_
timestamp 1667941163
transform 1 0 2576 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1423_
timestamp 1667941163
transform 1 0 3956 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1424__178
timestamp 1667941163
transform 1 0 5704 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1424_
timestamp 1667941163
transform 1 0 5244 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1425_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1426_
timestamp 1667941163
transform 1 0 3956 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1427_
timestamp 1667941163
transform 1 0 9292 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1428_
timestamp 1667941163
transform 1 0 4784 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1429_
timestamp 1667941163
transform 1 0 4048 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1430_
timestamp 1667941163
transform 1 0 18768 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1431_
timestamp 1667941163
transform 1 0 2024 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1432_
timestamp 1667941163
transform 1 0 3956 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1433_
timestamp 1667941163
transform 1 0 12236 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1434_
timestamp 1667941163
transform 1 0 6532 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1435_
timestamp 1667941163
transform 1 0 8096 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1436_
timestamp 1667941163
transform 1 0 20332 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1437_
timestamp 1667941163
transform 1 0 18492 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1438_
timestamp 1667941163
transform 1 0 30268 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1439_
timestamp 1667941163
transform 1 0 28244 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1440__179
timestamp 1667941163
transform 1 0 30636 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1440_
timestamp 1667941163
transform 1 0 30452 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1441_
timestamp 1667941163
transform 1 0 27140 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1442_
timestamp 1667941163
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1443_
timestamp 1667941163
transform 1 0 28244 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1444_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1445_
timestamp 1667941163
transform 1 0 28612 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1446_
timestamp 1667941163
transform 1 0 29624 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1447_
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1448_
timestamp 1667941163
transform 1 0 29072 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1449_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1450_
timestamp 1667941163
transform 1 0 28428 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1451_
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1452_
timestamp 1667941163
transform 1 0 25852 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1453_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1454_
timestamp 1667941163
transform 1 0 14260 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1455_
timestamp 1667941163
transform 1 0 14260 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1456_
timestamp 1667941163
transform 1 0 9752 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1456__180
timestamp 1667941163
transform 1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1457_
timestamp 1667941163
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1458_
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1459_
timestamp 1667941163
transform 1 0 17664 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1460_
timestamp 1667941163
transform 1 0 22264 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1461_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1462_
timestamp 1667941163
transform 1 0 16560 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1463_
timestamp 1667941163
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1464_
timestamp 1667941163
transform 1 0 17296 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1465_
timestamp 1667941163
transform 1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1466_
timestamp 1667941163
transform 1 0 14260 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1467_
timestamp 1667941163
transform 1 0 18400 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1468_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1469_
timestamp 1667941163
transform 1 0 13984 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1470_
timestamp 1667941163
transform 1 0 19596 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1471_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1472__181
timestamp 1667941163
transform 1 0 23736 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1472_
timestamp 1667941163
transform 1 0 25024 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1473_
timestamp 1667941163
transform 1 0 16100 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1474_
timestamp 1667941163
transform 1 0 28520 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1475_
timestamp 1667941163
transform 1 0 16836 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1476_
timestamp 1667941163
transform 1 0 25208 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1477_
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1478_
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1479_
timestamp 1667941163
transform 1 0 24564 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1480_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1481_
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1482_
timestamp 1667941163
transform 1 0 18584 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1483_
timestamp 1667941163
transform 1 0 19320 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1484_
timestamp 1667941163
transform 1 0 22448 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1485_
timestamp 1667941163
transform 1 0 15180 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1486_
timestamp 1667941163
transform 1 0 10672 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1487_
timestamp 1667941163
transform 1 0 9936 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1488__182
timestamp 1667941163
transform 1 0 11776 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1488_
timestamp 1667941163
transform 1 0 11592 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1489_
timestamp 1667941163
transform 1 0 7452 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1490_
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1491_
timestamp 1667941163
transform 1 0 9108 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1492_
timestamp 1667941163
transform 1 0 15916 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1493_
timestamp 1667941163
transform 1 0 16008 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1494_
timestamp 1667941163
transform 1 0 10396 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1495_
timestamp 1667941163
transform 1 0 7820 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1496_
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1497_
timestamp 1667941163
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1498_
timestamp 1667941163
transform 1 0 9108 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1499_
timestamp 1667941163
transform 1 0 7360 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1500_
timestamp 1667941163
transform 1 0 18400 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1501_
timestamp 1667941163
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1502_
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1503_
timestamp 1667941163
transform 1 0 16836 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1504_
timestamp 1667941163
transform 1 0 13984 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1504__183
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1505_
timestamp 1667941163
transform 1 0 22356 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1506_
timestamp 1667941163
transform 1 0 23736 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1507_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1508_
timestamp 1667941163
transform 1 0 21988 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1509_
timestamp 1667941163
transform 1 0 22172 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1510_
timestamp 1667941163
transform 1 0 27784 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1511_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1512_
timestamp 1667941163
transform 1 0 23276 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1513_
timestamp 1667941163
transform 1 0 19504 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1514_
timestamp 1667941163
transform 1 0 14260 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1515_
timestamp 1667941163
transform 1 0 25576 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1516_
timestamp 1667941163
transform 1 0 27140 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1517_
timestamp 1667941163
transform 1 0 25392 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1518_
timestamp 1667941163
transform 1 0 15180 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1519_
timestamp 1667941163
transform 1 0 15088 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1520__184
timestamp 1667941163
transform 1 0 4416 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1520_
timestamp 1667941163
transform 1 0 4784 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1521_
timestamp 1667941163
transform 1 0 20424 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1522_
timestamp 1667941163
transform 1 0 24564 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1523_
timestamp 1667941163
transform 1 0 16836 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1524_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1525_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1526_
timestamp 1667941163
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1527_
timestamp 1667941163
transform 1 0 4600 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1528_
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1529_
timestamp 1667941163
transform 1 0 17756 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1530_
timestamp 1667941163
transform 1 0 2116 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1531_
timestamp 1667941163
transform 1 0 19412 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1532_
timestamp 1667941163
transform 1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1533_
timestamp 1667941163
transform 1 0 16836 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1534_
timestamp 1667941163
transform 1 0 13892 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1535_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1536__185
timestamp 1667941163
transform 1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1536_
timestamp 1667941163
transform 1 0 8740 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1537_
timestamp 1667941163
transform 1 0 18676 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1538_
timestamp 1667941163
transform 1 0 22172 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1539_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1540_
timestamp 1667941163
transform 1 0 22540 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1541_
timestamp 1667941163
transform 1 0 24564 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1542_
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1543_
timestamp 1667941163
transform 1 0 21988 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1544_
timestamp 1667941163
transform 1 0 25484 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1545_
timestamp 1667941163
transform 1 0 26956 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1546_
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1547_
timestamp 1667941163
transform 1 0 20332 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1548_
timestamp 1667941163
transform 1 0 17112 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1549_
timestamp 1667941163
transform 1 0 17756 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1550_
timestamp 1667941163
transform 1 0 14260 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1551_
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1552__186
timestamp 1667941163
transform 1 0 18768 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1552_
timestamp 1667941163
transform 1 0 19412 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1553_
timestamp 1667941163
transform 1 0 19136 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1554_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1555_
timestamp 1667941163
transform 1 0 22816 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1556_
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1557_
timestamp 1667941163
transform 1 0 15548 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1558_
timestamp 1667941163
transform 1 0 9108 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1559_
timestamp 1667941163
transform 1 0 16376 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1560_
timestamp 1667941163
transform 1 0 18124 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1561_
timestamp 1667941163
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1562_
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1563_
timestamp 1667941163
transform 1 0 4876 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1564_
timestamp 1667941163
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1565_
timestamp 1667941163
transform 1 0 13892 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1566_
timestamp 1667941163
transform 1 0 16008 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1567_
timestamp 1667941163
transform 1 0 10856 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1568__187
timestamp 1667941163
transform 1 0 12420 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1568_
timestamp 1667941163
transform 1 0 12328 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1569_
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1570_
timestamp 1667941163
transform 1 0 25484 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1571_
timestamp 1667941163
transform 1 0 10028 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1572_
timestamp 1667941163
transform 1 0 22080 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1573_
timestamp 1667941163
transform 1 0 22172 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1574_
timestamp 1667941163
transform 1 0 24656 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1575_
timestamp 1667941163
transform 1 0 24840 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1576_
timestamp 1667941163
transform 1 0 27140 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1577_
timestamp 1667941163
transform 1 0 21252 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1578_
timestamp 1667941163
transform 1 0 16468 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1579_
timestamp 1667941163
transform 1 0 27140 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1580_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1581_
timestamp 1667941163
transform 1 0 26128 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1582_
timestamp 1667941163
transform 1 0 16468 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1583_
timestamp 1667941163
transform 1 0 14260 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1584_
timestamp 1667941163
transform 1 0 20700 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1585__188
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1585_
timestamp 1667941163
transform 1 0 13524 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1586_
timestamp 1667941163
transform 1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1587_
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1588_
timestamp 1667941163
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1589_
timestamp 1667941163
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1590_
timestamp 1667941163
transform 1 0 15180 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1591_
timestamp 1667941163
transform 1 0 6532 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1592_
timestamp 1667941163
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1593_
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1594_
timestamp 1667941163
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1595_
timestamp 1667941163
transform 1 0 24932 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1596_
timestamp 1667941163
transform 1 0 27416 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1597__189
timestamp 1667941163
transform 1 0 29716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1597_
timestamp 1667941163
transform 1 0 28888 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1598_
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1599_
timestamp 1667941163
transform 1 0 24840 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1600_
timestamp 1667941163
transform 1 0 23920 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1601_
timestamp 1667941163
transform 1 0 26956 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1602_
timestamp 1667941163
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1603_
timestamp 1667941163
transform 1 0 25760 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1604_
timestamp 1667941163
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1605_
timestamp 1667941163
transform 1 0 25760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1606_
timestamp 1667941163
transform 1 0 18952 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1607_
timestamp 1667941163
transform 1 0 22724 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1608_
timestamp 1667941163
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1609_
timestamp 1667941163
transform 1 0 25208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1609__190
timestamp 1667941163
transform 1 0 27784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1610_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1611_
timestamp 1667941163
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1612_
timestamp 1667941163
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1613_
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1614_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1615_
timestamp 1667941163
transform 1 0 25760 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1616_
timestamp 1667941163
transform 1 0 23644 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1617_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1618_
timestamp 1667941163
transform 1 0 18400 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1619_
timestamp 1667941163
transform 1 0 16928 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1620_
timestamp 1667941163
transform 1 0 18032 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1621_
timestamp 1667941163
transform 1 0 16468 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1621__191
timestamp 1667941163
transform 1 0 16468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1622_
timestamp 1667941163
transform 1 0 20700 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1623_
timestamp 1667941163
transform 1 0 22448 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1624_
timestamp 1667941163
transform 1 0 5152 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1625_
timestamp 1667941163
transform 1 0 20976 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1626_
timestamp 1667941163
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1627_
timestamp 1667941163
transform 1 0 18676 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1628_
timestamp 1667941163
transform 1 0 19412 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1629_
timestamp 1667941163
transform 1 0 20608 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3956 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 6532 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 4140 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 10120 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 4140 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 9108 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 10028 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 10212 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 7268 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 37352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1667941163
transform 1 0 6532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1667941163
transform 1 0 37996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1667941163
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1667941163
transform 1 0 2300 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1667941163
transform 1 0 37996 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1667941163
transform 1 0 3036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 18308 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1667941163
transform 1 0 22632 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1667941163
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1667941163
transform 1 0 37444 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1667941163
transform 1 0 9108 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1667941163
transform 1 0 5152 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1667941163
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 36156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1667941163
transform 1 0 37444 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1667941163
transform 1 0 38088 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1667941163
transform 1 0 38088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1667941163
transform 1 0 10304 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1667941163
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1667941163
transform 1 0 37444 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1667941163
transform 1 0 36708 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1667941163
transform 1 0 14904 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1667941163
transform 1 0 17480 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1667941163
transform 1 0 37444 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1667941163
transform 1 0 3496 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1667941163
transform 1 0 15548 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1667941163
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1667941163
transform 1 0 37996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1667941163
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1667941163
transform 1 0 37444 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1667941163
transform 1 0 36708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1667941163
transform 1 0 1564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 38088 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1667941163
transform 1 0 37996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1667941163
transform 1 0 23920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1667941163
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1667941163
transform 1 0 20608 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1667941163
transform 1 0 3956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1667941163
transform 1 0 38088 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1667941163
transform 1 0 30912 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1667941163
transform 1 0 37444 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1667941163
transform 1 0 32936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1667941163
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1667941163
transform 1 0 16008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 22632 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1667941163
transform 1 0 37444 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1667941163
transform 1 0 37444 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 2208 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 38088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 2852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 38088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1667941163
transform 1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1667941163
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1667941163
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1667941163
transform 1 0 38088 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1667941163
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1667941163
transform 1 0 29072 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1667941163
transform 1 0 28612 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1667941163
transform 1 0 2300 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1667941163
transform 1 0 6532 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1667941163
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1667941163
transform 1 0 25760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output95 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 3220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 4600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 1564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 2668 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 37996 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 23276 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 1564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 4324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 3956 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 37260 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 21988 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1667941163
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1667941163
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1667941163
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1667941163
transform 1 0 12972 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1667941163
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1667941163
transform 1 0 6532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1667941163
transform 1 0 35880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1667941163
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1667941163
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1667941163
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1667941163
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1667941163
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1667941163
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1667941163
transform 1 0 4508 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1667941163
transform 1 0 19412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1667941163
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1667941163
transform 1 0 33764 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 0 nsew signal input
flabel metal2 s 39302 200 39358 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 1 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 2 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 3 nsew signal input
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 ccff_head
port 4 nsew signal input
flabel metal2 s 25134 39200 25190 39800 0 FreeSans 224 90 0 0 ccff_tail
port 5 nsew signal tristate
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 39200 2728 39800 2848 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal2 s 38014 39200 38070 39800 0 FreeSans 224 90 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal2 s 18694 200 18750 800 0 FreeSans 224 90 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 16 nsew signal input
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 17 nsew signal input
flabel metal2 s 17406 39200 17462 39800 0 FreeSans 224 90 0 0 chanx_left_in[3]
port 18 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chanx_left_in[4]
port 19 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 chanx_left_in[5]
port 20 nsew signal input
flabel metal3 s 39200 31288 39800 31408 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 21 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 22 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chanx_left_in[8]
port 23 nsew signal input
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 24 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 25 nsew signal tristate
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 26 nsew signal tristate
flabel metal3 s 39200 38088 39800 38208 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 27 nsew signal tristate
flabel metal2 s 4526 39200 4582 39800 0 FreeSans 224 90 0 0 chanx_left_out[12]
port 28 nsew signal tristate
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chanx_left_out[13]
port 29 nsew signal tristate
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 30 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_left_out[15]
port 31 nsew signal tristate
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_left_out[16]
port 32 nsew signal tristate
flabel metal3 s 200 27888 800 28008 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 33 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 34 nsew signal tristate
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chanx_left_out[1]
port 35 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 36 nsew signal tristate
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chanx_left_out[3]
port 37 nsew signal tristate
flabel metal2 s 1306 39200 1362 39800 0 FreeSans 224 90 0 0 chanx_left_out[4]
port 38 nsew signal tristate
flabel metal2 s 28354 200 28410 800 0 FreeSans 224 90 0 0 chanx_left_out[5]
port 39 nsew signal tristate
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 chanx_left_out[6]
port 40 nsew signal tristate
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 41 nsew signal tristate
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chanx_left_out[8]
port 42 nsew signal tristate
flabel metal2 s 31574 39200 31630 39800 0 FreeSans 224 90 0 0 chanx_left_out[9]
port 43 nsew signal tristate
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 44 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 45 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 46 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 47 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 48 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 49 nsew signal input
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 50 nsew signal input
flabel metal2 s 36726 39200 36782 39800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 51 nsew signal input
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 52 nsew signal input
flabel metal3 s 39200 19728 39800 19848 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 53 nsew signal input
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chanx_right_in[1]
port 54 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 55 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chanx_right_in[3]
port 56 nsew signal input
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 57 nsew signal input
flabel metal2 s 26422 200 26478 800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 58 nsew signal input
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_right_in[6]
port 59 nsew signal input
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chanx_right_in[7]
port 60 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 61 nsew signal input
flabel metal2 s 17406 200 17462 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 62 nsew signal input
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 63 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 64 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 65 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 66 nsew signal tristate
flabel metal3 s 39200 14288 39800 14408 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 67 nsew signal tristate
flabel metal2 s 23846 200 23902 800 0 FreeSans 224 90 0 0 chanx_right_out[14]
port 68 nsew signal tristate
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 69 nsew signal tristate
flabel metal2 s 27066 39200 27122 39800 0 FreeSans 224 90 0 0 chanx_right_out[16]
port 70 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 71 nsew signal tristate
flabel metal2 s 10966 39200 11022 39800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 72 nsew signal tristate
flabel metal3 s 39200 24488 39800 24608 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 73 nsew signal tristate
flabel metal2 s 1306 200 1362 800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 74 nsew signal tristate
flabel metal2 s 12254 200 12310 800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 75 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 76 nsew signal tristate
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 77 nsew signal tristate
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 78 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chanx_right_out[7]
port 79 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 80 nsew signal tristate
flabel metal3 s 200 2728 800 2848 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 81 nsew signal tristate
flabel metal3 s 39200 16328 39800 16448 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 82 nsew signal input
flabel metal3 s 39200 9528 39800 9648 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 83 nsew signal input
flabel metal3 s 200 29928 800 30048 0 FreeSans 480 0 0 0 chany_bottom_in[11]
port 84 nsew signal input
flabel metal2 s 15474 39200 15530 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 85 nsew signal input
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 86 nsew signal input
flabel metal3 s 39200 33328 39800 33448 0 FreeSans 480 0 0 0 chany_bottom_in[14]
port 87 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 88 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 chany_bottom_in[16]
port 89 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[17]
port 90 nsew signal input
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chany_bottom_in[18]
port 91 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 92 nsew signal input
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 chany_bottom_in[2]
port 93 nsew signal input
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 94 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 95 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 96 nsew signal input
flabel metal3 s 39200 21088 39800 21208 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 97 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chany_bottom_in[7]
port 98 nsew signal input
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 99 nsew signal input
flabel metal2 s 20626 39200 20682 39800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 100 nsew signal input
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 101 nsew signal tristate
flabel metal3 s 200 36728 800 36848 0 FreeSans 480 0 0 0 chany_bottom_out[10]
port 102 nsew signal tristate
flabel metal3 s 39200 36728 39800 36848 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 103 nsew signal tristate
flabel metal3 s 200 1368 800 1488 0 FreeSans 480 0 0 0 chany_bottom_out[12]
port 104 nsew signal tristate
flabel metal2 s 21914 39200 21970 39800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 105 nsew signal tristate
flabel metal3 s 200 18368 800 18488 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 106 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 107 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 108 nsew signal tristate
flabel metal2 s 5814 200 5870 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 109 nsew signal tristate
flabel metal3 s 39200 4768 39800 4888 0 FreeSans 480 0 0 0 chany_bottom_out[18]
port 110 nsew signal tristate
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 111 nsew signal tristate
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 112 nsew signal tristate
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 113 nsew signal tristate
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 114 nsew signal tristate
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 115 nsew signal tristate
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chany_bottom_out[6]
port 116 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_bottom_out[7]
port 117 nsew signal tristate
flabel metal2 s 12898 39200 12954 39800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 118 nsew signal tristate
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_bottom_out[9]
port 119 nsew signal tristate
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chany_top_in[0]
port 120 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 121 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_in[11]
port 122 nsew signal input
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chany_top_in[12]
port 123 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chany_top_in[13]
port 124 nsew signal input
flabel metal3 s 39200 11568 39800 11688 0 FreeSans 480 0 0 0 chany_top_in[14]
port 125 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 126 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_top_in[16]
port 127 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 128 nsew signal input
flabel metal2 s 32862 200 32918 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 129 nsew signal input
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 130 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 131 nsew signal input
flabel metal3 s 200 14968 800 15088 0 FreeSans 480 0 0 0 chany_top_in[3]
port 132 nsew signal input
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_in[4]
port 133 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chany_top_in[5]
port 134 nsew signal input
flabel metal2 s 34794 200 34850 800 0 FreeSans 224 90 0 0 chany_top_in[6]
port 135 nsew signal input
flabel metal3 s 200 19728 800 19848 0 FreeSans 480 0 0 0 chany_top_in[7]
port 136 nsew signal input
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chany_top_in[8]
port 137 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chany_top_in[9]
port 138 nsew signal input
flabel metal3 s 200 12928 800 13048 0 FreeSans 480 0 0 0 chany_top_out[0]
port 139 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_top_out[10]
port 140 nsew signal tristate
flabel metal2 s 38014 200 38070 800 0 FreeSans 224 90 0 0 chany_top_out[11]
port 141 nsew signal tristate
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_out[12]
port 142 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_top_out[13]
port 143 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chany_top_out[14]
port 144 nsew signal tristate
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_out[15]
port 145 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[16]
port 146 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_top_out[17]
port 147 nsew signal tristate
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chany_top_out[18]
port 148 nsew signal tristate
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chany_top_out[1]
port 149 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chany_top_out[2]
port 150 nsew signal tristate
flabel metal3 s 200 25168 800 25288 0 FreeSans 480 0 0 0 chany_top_out[3]
port 151 nsew signal tristate
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 152 nsew signal tristate
flabel metal2 s 2594 200 2650 800 0 FreeSans 224 90 0 0 chany_top_out[5]
port 153 nsew signal tristate
flabel metal3 s 200 6128 800 6248 0 FreeSans 480 0 0 0 chany_top_out[6]
port 154 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 155 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 chany_top_out[8]
port 156 nsew signal tristate
flabel metal2 s 33506 39200 33562 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 157 nsew signal tristate
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 158 nsew signal input
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 159 nsew signal input
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 160 nsew signal input
flabel metal2 s 7746 200 7802 800 0 FreeSans 224 90 0 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 161 nsew signal input
flabel metal2 s 14186 200 14242 800 0 FreeSans 224 90 0 0 pReset
port 162 nsew signal input
flabel metal3 s 200 8168 800 8288 0 FreeSans 480 0 0 0 prog_clk
port 163 nsew signal input
flabel metal3 s 39200 26528 39800 26648 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 164 nsew signal input
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 165 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 166 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 167 nsew signal input
flabel metal2 s 18 39200 74 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
port 168 nsew signal input
flabel metal2 s 6458 39200 6514 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
port 169 nsew signal input
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 170 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 171 nsew signal input
flabel metal3 s 200 34688 800 34808 0 FreeSans 480 0 0 0 vccd1
port 172 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 172 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 172 nsew signal bidirectional
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 vssd1
port 173 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 173 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 10810 12206 10810 12206 0 _0000_
rlabel metal1 18400 6970 18400 6970 0 _0001_
rlabel metal1 3365 10642 3365 10642 0 _0002_
rlabel metal1 4646 19448 4646 19448 0 _0003_
rlabel metal1 13439 23018 13439 23018 0 _0004_
rlabel metal1 12151 17578 12151 17578 0 _0005_
rlabel metal2 11086 20468 11086 20468 0 _0006_
rlabel metal1 8103 14314 8103 14314 0 _0007_
rlabel metal1 8234 5032 8234 5032 0 _0008_
rlabel metal2 9982 1870 9982 1870 0 _0009_
rlabel metal3 17204 14960 17204 14960 0 _0010_
rlabel metal1 3457 17578 3457 17578 0 _0011_
rlabel metal2 12558 21165 12558 21165 0 _0012_
rlabel metal3 15985 27676 15985 27676 0 _0013_
rlabel metal1 18216 25126 18216 25126 0 _0014_
rlabel via3 17733 26316 17733 26316 0 _0015_
rlabel metal1 6716 6426 6716 6426 0 _0016_
rlabel metal2 12374 4335 12374 4335 0 _0017_
rlabel via2 7130 5355 7130 5355 0 _0018_
rlabel metal1 14398 1734 14398 1734 0 _0019_
rlabel metal2 13754 4471 13754 4471 0 _0020_
rlabel metal1 5382 8983 5382 8983 0 _0021_
rlabel metal2 7774 4012 7774 4012 0 _0022_
rlabel metal2 4554 7310 4554 7310 0 _0023_
rlabel metal2 12650 17204 12650 17204 0 _0024_
rlabel metal2 6670 13877 6670 13877 0 _0025_
rlabel metal1 6164 7446 6164 7446 0 _0026_
rlabel metal2 9752 14756 9752 14756 0 _0027_
rlabel metal2 14858 5049 14858 5049 0 _0028_
rlabel metal2 13018 6426 13018 6426 0 _0029_
rlabel metal1 11270 3978 11270 3978 0 _0030_
rlabel metal1 12558 8976 12558 8976 0 _0031_
rlabel metal2 13570 5304 13570 5304 0 _0032_
rlabel metal1 8418 3910 8418 3910 0 _0033_
rlabel metal1 8517 8534 8517 8534 0 _0034_
rlabel metal1 13846 7480 13846 7480 0 _0035_
rlabel metal1 11178 3706 11178 3706 0 _0036_
rlabel metal1 10028 3910 10028 3910 0 _0037_
rlabel metal1 7215 13226 7215 13226 0 _0038_
rlabel metal1 5941 11730 5941 11730 0 _0039_
rlabel metal1 3457 20842 3457 20842 0 _0040_
rlabel metal1 1971 22678 1971 22678 0 _0041_
rlabel metal1 3135 24106 3135 24106 0 _0042_
rlabel metal2 2898 19023 2898 19023 0 _0043_
rlabel via3 6509 20196 6509 20196 0 _0044_
rlabel metal2 598 23256 598 23256 0 _0045_
rlabel metal1 15916 29138 15916 29138 0 _0046_
rlabel metal1 11684 9146 11684 9146 0 _0047_
rlabel metal2 5566 25262 5566 25262 0 _0048_
rlabel metal1 7643 19754 7643 19754 0 _0049_
rlabel metal1 4830 22066 4830 22066 0 _0050_
rlabel metal1 5336 29478 5336 29478 0 _0051_
rlabel metal1 6355 20910 6355 20910 0 _0052_
rlabel metal1 4791 21590 4791 21590 0 _0053_
rlabel metal1 3365 23018 3365 23018 0 _0054_
rlabel metal1 3641 20502 3641 20502 0 _0055_
rlabel metal1 14405 25194 14405 25194 0 _0056_
rlabel via2 12466 22763 12466 22763 0 _0057_
rlabel metal1 11323 24106 11323 24106 0 _0058_
rlabel metal1 14536 25806 14536 25806 0 _0059_
rlabel metal2 12466 14773 12466 14773 0 _0060_
rlabel metal1 10817 13226 10817 13226 0 _0061_
rlabel metal1 14858 3910 14858 3910 0 _0062_
rlabel metal2 5980 7140 5980 7140 0 _0063_
rlabel metal1 18032 5882 18032 5882 0 _0064_
rlabel metal2 4094 6987 4094 6987 0 _0065_
rlabel metal1 4646 5576 4646 5576 0 _0066_
rlabel via2 21390 6171 21390 6171 0 _0067_
rlabel metal2 6854 2638 6854 2638 0 _0068_
rlabel metal2 12926 5474 12926 5474 0 _0069_
rlabel metal1 14129 12206 14129 12206 0 _0070_
rlabel metal1 14122 16490 14122 16490 0 _0071_
rlabel metal2 27278 16490 27278 16490 0 _0072_
rlabel metal1 11599 18666 11599 18666 0 _0073_
rlabel metal1 10120 20026 10120 20026 0 _0074_
rlabel metal3 13432 15300 13432 15300 0 _0075_
rlabel via2 14674 4811 14674 4811 0 _0076_
rlabel metal2 13294 16864 13294 16864 0 _0077_
rlabel metal1 13386 20774 13386 20774 0 _0078_
rlabel metal2 18170 5151 18170 5151 0 _0079_
rlabel metal1 6171 24174 6171 24174 0 _0080_
rlabel metal1 2668 26758 2668 26758 0 _0081_
rlabel metal1 5796 29546 5796 29546 0 _0082_
rlabel metal3 7682 21692 7682 21692 0 _0083_
rlabel metal2 5382 17850 5382 17850 0 _0084_
rlabel metal4 13156 12772 13156 12772 0 _0085_
rlabel metal1 8011 23086 8011 23086 0 _0086_
rlabel metal2 15778 29257 15778 29257 0 _0087_
rlabel metal1 14398 1802 14398 1802 0 _0088_
rlabel metal1 9752 3638 9752 3638 0 _0089_
rlabel metal2 8510 3859 8510 3859 0 _0090_
rlabel metal2 7314 8109 7314 8109 0 _0091_
rlabel metal1 13110 13865 13110 13865 0 _0092_
rlabel metal1 9062 16007 9062 16007 0 _0093_
rlabel metal1 9515 17238 9515 17238 0 _0094_
rlabel metal1 13294 17748 13294 17748 0 _0095_
rlabel metal2 13018 3281 13018 3281 0 _0096_
rlabel metal1 3871 2346 3871 2346 0 _0097_
rlabel via1 6946 5117 6946 5117 0 _0098_
rlabel metal2 8234 4233 8234 4233 0 _0099_
rlabel metal1 14030 1496 14030 1496 0 _0100_
rlabel metal1 21436 6358 21436 6358 0 _0101_
rlabel metal1 12282 3706 12282 3706 0 _0102_
rlabel metal1 9706 3094 9706 3094 0 _0103_
rlabel metal1 12466 17544 12466 17544 0 _0104_
rlabel metal2 3910 15419 3910 15419 0 _0105_
rlabel metal4 6900 18292 6900 18292 0 _0106_
rlabel metal1 11178 5678 11178 5678 0 _0107_
rlabel metal2 11086 5899 11086 5899 0 _0108_
rlabel metal2 12466 15997 12466 15997 0 _0109_
rlabel metal1 9430 12206 9430 12206 0 _0110_
rlabel via2 4002 9605 4002 9605 0 _0111_
rlabel via2 27278 18139 27278 18139 0 _0112_
rlabel metal4 19320 21420 19320 21420 0 _0113_
rlabel metal2 17066 15912 17066 15912 0 _0114_
rlabel metal2 9062 4947 9062 4947 0 _0115_
rlabel metal2 14306 4063 14306 4063 0 _0116_
rlabel metal1 8195 12886 8195 12886 0 _0117_
rlabel metal1 16330 12920 16330 12920 0 _0118_
rlabel metal1 19550 6290 19550 6290 0 _0119_
rlabel metal1 10587 24854 10587 24854 0 _0120_
rlabel metal2 18814 25024 18814 25024 0 _0121_
rlabel metal1 8655 25262 8655 25262 0 _0122_
rlabel metal1 9207 24106 9207 24106 0 _0123_
rlabel metal1 17434 20536 17434 20536 0 _0124_
rlabel metal1 14444 22066 14444 22066 0 _0125_
rlabel metal1 13301 20502 13301 20502 0 _0126_
rlabel metal1 13439 24174 13439 24174 0 _0127_
rlabel metal2 14398 1836 14398 1836 0 _0128_
rlabel metal2 2990 3179 2990 3179 0 _0129_
rlabel metal3 10810 2244 10810 2244 0 _0130_
rlabel metal1 14030 2822 14030 2822 0 _0131_
rlabel metal1 14122 14314 14122 14314 0 _0132_
rlabel metal1 8149 16490 8149 16490 0 _0133_
rlabel metal1 28934 15130 28934 15130 0 _0134_
rlabel metal2 15594 5831 15594 5831 0 _0135_
rlabel metal1 10534 4794 10534 4794 0 _0136_
rlabel metal1 11546 4114 11546 4114 0 _0137_
rlabel metal2 13662 5729 13662 5729 0 _0138_
rlabel metal2 11408 9044 11408 9044 0 _0139_
rlabel metal2 13662 1904 13662 1904 0 _0140_
rlabel metal2 9522 4998 9522 4998 0 _0141_
rlabel metal2 17066 4199 17066 4199 0 _0142_
rlabel metal1 11638 4794 11638 4794 0 _0143_
rlabel metal1 13202 4114 13202 4114 0 _0144_
rlabel metal2 9890 5304 9890 5304 0 _0145_
rlabel metal2 14858 11288 14858 11288 0 _0146_
rlabel metal1 20631 5270 20631 5270 0 _0147_
rlabel metal2 17986 5644 17986 5644 0 _0148_
rlabel metal1 2622 4250 2622 4250 0 _0149_
rlabel metal2 17526 5049 17526 5049 0 _0150_
rlabel metal1 7774 15912 7774 15912 0 _0151_
rlabel metal2 15870 13362 15870 13362 0 _0152_
rlabel metal1 8142 11186 8142 11186 0 _0153_
rlabel metal3 12903 22372 12903 22372 0 _0154_
rlabel metal2 17158 21471 17158 21471 0 _0155_
rlabel metal1 6762 7310 6762 7310 0 _0156_
rlabel metal1 13570 3026 13570 3026 0 _0157_
rlabel metal1 7682 30192 7682 30192 0 _0158_
rlabel metal1 13892 17714 13892 17714 0 _0159_
rlabel metal1 20194 4590 20194 4590 0 _0160_
rlabel metal2 8418 20468 8418 20468 0 _0161_
rlabel metal1 15226 29614 15226 29614 0 _0162_
rlabel metal2 20102 5610 20102 5610 0 _0163_
rlabel metal2 27738 13787 27738 13787 0 _0164_
rlabel metal1 14168 4114 14168 4114 0 _0165_
rlabel metal1 16606 2550 16606 2550 0 _0166_
rlabel metal1 29854 14926 29854 14926 0 _0167_
rlabel metal1 2346 4046 2346 4046 0 _0168_
rlabel metal1 14306 12886 14306 12886 0 _0169_
rlabel metal2 8280 22066 8280 22066 0 _0170_
rlabel metal2 1702 27557 1702 27557 0 _0171_
rlabel metal1 20010 24106 20010 24106 0 _0172_
rlabel metal2 13662 20502 13662 20502 0 _0173_
rlabel metal2 15410 15997 15410 15997 0 _0174_
rlabel metal2 22310 13158 22310 13158 0 _0175_
rlabel metal1 20332 16150 20332 16150 0 _0176_
rlabel metal1 19550 15096 19550 15096 0 _0177_
rlabel metal1 18400 22202 18400 22202 0 _0178_
rlabel metal2 22586 23528 22586 23528 0 _0179_
rlabel metal1 20608 22406 20608 22406 0 _0180_
rlabel metal3 11109 20876 11109 20876 0 _0181_
rlabel metal1 19274 27030 19274 27030 0 _0182_
rlabel metal1 14306 9622 14306 9622 0 _0183_
rlabel metal1 13616 28118 13616 28118 0 _0184_
rlabel via2 25990 20859 25990 20859 0 _0185_
rlabel metal1 13984 23766 13984 23766 0 _0186_
rlabel metal1 17986 4726 17986 4726 0 _0187_
rlabel metal1 15180 29206 15180 29206 0 _0188_
rlabel metal1 15134 27370 15134 27370 0 _0189_
rlabel metal1 19642 29512 19642 29512 0 _0190_
rlabel metal2 18354 23800 18354 23800 0 _0191_
rlabel metal1 16652 22678 16652 22678 0 _0192_
rlabel metal1 22540 24922 22540 24922 0 _0193_
rlabel metal1 14720 28458 14720 28458 0 _0194_
rlabel metal2 20010 30872 20010 30872 0 _0195_
rlabel metal1 22494 29818 22494 29818 0 _0196_
rlabel metal2 12742 27302 12742 27302 0 _0197_
rlabel metal1 20286 27336 20286 27336 0 _0198_
rlabel metal2 23690 23970 23690 23970 0 _0199_
rlabel metal1 14536 30294 14536 30294 0 _0200_
rlabel metal1 11822 5542 11822 5542 0 _0201_
rlabel metal1 21344 6834 21344 6834 0 _0202_
rlabel metal1 16376 3706 16376 3706 0 _0203_
rlabel metal1 4784 31858 4784 31858 0 _0204_
rlabel metal2 20102 6545 20102 6545 0 _0205_
rlabel metal1 11914 25976 11914 25976 0 _0206_
rlabel metal1 8786 25670 8786 25670 0 _0207_
rlabel metal2 19366 23290 19366 23290 0 _0208_
rlabel metal1 4416 24378 4416 24378 0 _0209_
rlabel metal2 22034 10880 22034 10880 0 _0210_
rlabel metal2 21022 7769 21022 7769 0 _0211_
rlabel metal1 19734 7922 19734 7922 0 _0212_
rlabel metal1 16468 3910 16468 3910 0 _0213_
rlabel metal1 8234 25942 8234 25942 0 _0214_
rlabel metal1 15410 26282 15410 26282 0 _0215_
rlabel metal2 24058 7939 24058 7939 0 _0216_
rlabel metal1 24748 18054 24748 18054 0 _0217_
rlabel metal1 28934 19448 28934 19448 0 _0218_
rlabel metal1 21252 22406 21252 22406 0 _0219_
rlabel metal2 22586 20043 22586 20043 0 _0220_
rlabel metal2 31602 16728 31602 16728 0 _0221_
rlabel metal1 28704 20570 28704 20570 0 _0222_
rlabel metal2 28474 15640 28474 15640 0 _0223_
rlabel metal2 31234 14552 31234 14552 0 _0224_
rlabel metal1 28658 20808 28658 20808 0 _0225_
rlabel metal1 28727 16490 28727 16490 0 _0226_
rlabel metal1 26496 13974 26496 13974 0 _0227_
rlabel metal1 23690 18326 23690 18326 0 _0228_
rlabel metal1 19642 11322 19642 11322 0 _0229_
rlabel metal2 25346 21080 25346 21080 0 _0230_
rlabel metal2 30038 20026 30038 20026 0 _0231_
rlabel metal1 20194 8058 20194 8058 0 _0232_
rlabel metal2 24150 8228 24150 8228 0 _0233_
rlabel metal2 20190 8466 20190 8466 0 _0234_
rlabel metal2 30866 10574 30866 10574 0 _0235_
rlabel metal1 19228 18394 19228 18394 0 _0236_
rlabel metal1 20976 17850 20976 17850 0 _0237_
rlabel metal1 20700 8602 20700 8602 0 _0238_
rlabel metal1 22356 13498 22356 13498 0 _0239_
rlabel metal1 24380 15062 24380 15062 0 _0240_
rlabel metal2 22586 13090 22586 13090 0 _0241_
rlabel metal2 25346 11016 25346 11016 0 _0242_
rlabel metal2 21390 8704 21390 8704 0 _0243_
rlabel metal2 27370 9112 27370 9112 0 _0244_
rlabel metal1 23874 10234 23874 10234 0 _0245_
rlabel metal1 18584 7310 18584 7310 0 _0246_
rlabel metal1 22172 21318 22172 21318 0 _0247_
rlabel metal1 17894 18224 17894 18224 0 _0248_
rlabel metal1 11408 27030 11408 27030 0 _0249_
rlabel metal1 9522 27976 9522 27976 0 _0250_
rlabel metal1 7038 28118 7038 28118 0 _0251_
rlabel metal1 20976 24854 20976 24854 0 _0252_
rlabel metal1 12880 26282 12880 26282 0 _0253_
rlabel metal1 14582 29478 14582 29478 0 _0254_
rlabel metal2 21666 24174 21666 24174 0 _0255_
rlabel metal1 17250 24106 17250 24106 0 _0256_
rlabel metal1 12466 29206 12466 29206 0 _0257_
rlabel metal1 2438 31382 2438 31382 0 _0258_
rlabel metal1 18814 17272 18814 17272 0 _0259_
rlabel metal1 20064 19754 20064 19754 0 _0260_
rlabel metal4 6900 23528 6900 23528 0 _0261_
rlabel metal2 23414 26112 23414 26112 0 _0262_
rlabel metal1 24058 28186 24058 28186 0 _0263_
rlabel metal1 17848 16490 17848 16490 0 _0264_
rlabel metal2 2806 27676 2806 27676 0 _0265_
rlabel metal2 4186 26350 4186 26350 0 _0266_
rlabel metal1 4692 28118 4692 28118 0 _0267_
rlabel metal2 9338 26418 9338 26418 0 _0268_
rlabel metal1 4186 25976 4186 25976 0 _0269_
rlabel metal2 9522 28798 9522 28798 0 _0270_
rlabel metal2 5014 26010 5014 26010 0 _0271_
rlabel metal1 4462 24854 4462 24854 0 _0272_
rlabel metal1 18906 28730 18906 28730 0 _0273_
rlabel metal1 2346 23290 2346 23290 0 _0274_
rlabel metal2 2714 24038 2714 24038 0 _0275_
rlabel metal1 10810 18224 10810 18224 0 _0276_
rlabel metal1 6394 24854 6394 24854 0 _0277_
rlabel metal1 7774 27030 7774 27030 0 _0278_
rlabel metal1 20428 28118 20428 28118 0 _0279_
rlabel metal1 18768 19414 18768 19414 0 _0280_
rlabel metal1 30544 19414 30544 19414 0 _0281_
rlabel metal2 18814 21760 18814 21760 0 _0282_
rlabel metal1 30728 23766 30728 23766 0 _0283_
rlabel metal2 27370 23902 27370 23902 0 _0284_
rlabel metal2 24242 21794 24242 21794 0 _0285_
rlabel metal1 28474 22984 28474 22984 0 _0286_
rlabel metal1 29946 17544 29946 17544 0 _0287_
rlabel metal1 29716 15062 29716 15062 0 _0288_
rlabel metal1 30176 16150 30176 16150 0 _0289_
rlabel metal1 28244 24378 28244 24378 0 _0290_
rlabel metal2 28842 26792 28842 26792 0 _0291_
rlabel metal2 24978 23970 24978 23970 0 _0292_
rlabel metal2 28658 24582 28658 24582 0 _0293_
rlabel metal1 26174 22678 26174 22678 0 _0294_
rlabel metal1 26680 12886 26680 12886 0 _0295_
rlabel metal1 26910 24922 26910 24922 0 _0296_
rlabel metal1 13202 13770 13202 13770 0 _0297_
rlabel metal2 12742 24293 12742 24293 0 _0298_
rlabel metal1 1978 30770 1978 30770 0 _0299_
rlabel metal1 26496 15674 26496 15674 0 _0300_
rlabel metal4 12604 24208 12604 24208 0 _0301_
rlabel metal1 23644 13498 23644 13498 0 _0302_
rlabel metal1 22954 8058 22954 8058 0 _0303_
rlabel metal1 17059 16184 17059 16184 0 _0304_
rlabel metal1 17940 6698 17940 6698 0 _0305_
rlabel metal1 16698 11662 16698 11662 0 _0306_
rlabel metal1 18768 5882 18768 5882 0 _0307_
rlabel metal2 23782 11798 23782 11798 0 _0308_
rlabel metal1 14904 18666 14904 18666 0 _0309_
rlabel metal1 18975 21590 18975 21590 0 _0310_
rlabel metal2 19412 17170 19412 17170 0 _0311_
rlabel metal2 9982 14620 9982 14620 0 _0312_
rlabel metal2 20194 19635 20194 19635 0 _0313_
rlabel metal1 14766 20570 14766 20570 0 _0314_
rlabel metal1 19274 25704 19274 25704 0 _0315_
rlabel metal2 16330 26520 16330 26520 0 _0316_
rlabel metal1 29256 18326 29256 18326 0 _0317_
rlabel metal1 16606 24378 16606 24378 0 _0318_
rlabel metal1 25208 28186 25208 28186 0 _0319_
rlabel metal1 29624 21114 29624 21114 0 _0320_
rlabel metal1 22402 12308 22402 12308 0 _0321_
rlabel metal1 25208 16490 25208 16490 0 _0322_
rlabel metal2 27370 19822 27370 19822 0 _0323_
rlabel metal2 21298 21794 21298 21794 0 _0324_
rlabel metal2 18814 20944 18814 20944 0 _0325_
rlabel metal1 18676 25942 18676 25942 0 _0326_
rlabel metal2 22402 26962 22402 26962 0 _0327_
rlabel metal2 15410 16966 15410 16966 0 _0328_
rlabel metal1 10902 27336 10902 27336 0 _0329_
rlabel metal2 10166 26180 10166 26180 0 _0330_
rlabel metal1 4508 25262 4508 25262 0 _0331_
rlabel metal1 7314 22066 7314 22066 0 _0332_
rlabel metal1 18860 7446 18860 7446 0 _0333_
rlabel metal1 9522 27370 9522 27370 0 _0334_
rlabel metal1 17434 19856 17434 19856 0 _0335_
rlabel metal1 15916 25466 15916 25466 0 _0336_
rlabel via1 10630 29546 10630 29546 0 _0337_
rlabel metal2 8096 18700 8096 18700 0 _0338_
rlabel metal1 5658 14008 5658 14008 0 _0339_
rlabel metal3 9407 14892 9407 14892 0 _0340_
rlabel metal1 8740 20774 8740 20774 0 _0341_
rlabel metal1 7774 26282 7774 26282 0 _0342_
rlabel metal2 18630 28526 18630 28526 0 _0343_
rlabel metal1 17434 15130 17434 15130 0 _0344_
rlabel metal1 20056 6630 20056 6630 0 _0345_
rlabel metal2 27738 14756 27738 14756 0 _0346_
rlabel metal1 17802 5712 17802 5712 0 _0347_
rlabel metal1 22586 19448 22586 19448 0 _0348_
rlabel metal1 24334 22202 24334 22202 0 _0349_
rlabel metal1 22954 28118 22954 28118 0 _0350_
rlabel metal2 22218 15198 22218 15198 0 _0351_
rlabel metal1 22770 18666 22770 18666 0 _0352_
rlabel metal2 28014 12614 28014 12614 0 _0353_
rlabel metal1 22264 23766 22264 23766 0 _0354_
rlabel metal1 23552 21658 23552 21658 0 _0355_
rlabel metal1 19872 26282 19872 26282 0 _0356_
rlabel metal2 14490 13311 14490 13311 0 _0357_
rlabel metal2 25898 27234 25898 27234 0 _0358_
rlabel metal1 27784 17578 27784 17578 0 _0359_
rlabel metal2 25622 26078 25622 26078 0 _0360_
rlabel metal1 22586 10234 22586 10234 0 _0361_
rlabel metal2 17342 16031 17342 16031 0 _0362_
rlabel metal1 1886 17510 1886 17510 0 _0363_
rlabel metal2 21206 14144 21206 14144 0 _0364_
rlabel metal1 25208 7786 25208 7786 0 _0365_
rlabel metal1 17480 7446 17480 7446 0 _0366_
rlabel metal1 25070 15946 25070 15946 0 _0367_
rlabel metal1 22310 11322 22310 11322 0 _0368_
rlabel metal1 21482 9622 21482 9622 0 _0369_
rlabel metal3 14237 1292 14237 1292 0 _0370_
rlabel viali 20746 9549 20746 9549 0 _0371_
rlabel metal1 18492 8874 18492 8874 0 _0372_
rlabel via2 2346 25925 2346 25925 0 _0373_
rlabel metal2 21022 12614 21022 12614 0 _0374_
rlabel metal2 14582 11985 14582 11985 0 _0375_
rlabel metal2 17066 17000 17066 17000 0 _0376_
rlabel metal2 14122 26078 14122 26078 0 _0377_
rlabel metal1 8694 9622 8694 9622 0 _0378_
rlabel metal1 8694 29274 8694 29274 0 _0379_
rlabel metal1 19090 23766 19090 23766 0 _0380_
rlabel metal1 23046 22678 23046 22678 0 _0381_
rlabel metal2 18262 10438 18262 10438 0 _0382_
rlabel metal2 22770 26520 22770 26520 0 _0383_
rlabel metal1 24886 23018 24886 23018 0 _0384_
rlabel metal2 23690 21114 23690 21114 0 _0385_
rlabel metal1 22724 16150 22724 16150 0 _0386_
rlabel metal1 26082 19414 26082 19414 0 _0387_
rlabel metal1 27554 9962 27554 9962 0 _0388_
rlabel metal1 15732 7514 15732 7514 0 _0389_
rlabel metal1 21114 16150 21114 16150 0 _0390_
rlabel metal1 16790 23766 16790 23766 0 _0391_
rlabel metal1 20286 11866 20286 11866 0 _0392_
rlabel metal1 14720 19754 14720 19754 0 _0393_
rlabel metal1 10718 21352 10718 21352 0 _0394_
rlabel metal1 17112 26894 17112 26894 0 _0395_
rlabel metal1 19320 24854 19320 24854 0 _0396_
rlabel metal1 9384 21930 9384 21930 0 _0397_
rlabel metal1 23184 12954 23184 12954 0 _0398_
rlabel metal1 16422 21862 16422 21862 0 _0399_
rlabel metal2 15778 26622 15778 26622 0 _0400_
rlabel metal3 9223 9452 9223 9452 0 _0401_
rlabel metal1 16514 21114 16514 21114 0 _0402_
rlabel metal1 19136 9146 19136 9146 0 _0403_
rlabel metal1 26726 14790 26726 14790 0 _0404_
rlabel metal1 12144 18938 12144 18938 0 _0405_
rlabel metal1 5290 20502 5290 20502 0 _0406_
rlabel metal1 10672 28390 10672 28390 0 _0407_
rlabel metal3 7521 26316 7521 26316 0 _0408_
rlabel metal2 8326 18496 8326 18496 0 _0409_
rlabel metal1 10902 26282 10902 26282 0 _0410_
rlabel metal1 5750 26826 5750 26826 0 _0411_
rlabel metal1 12466 28424 12466 28424 0 _0412_
rlabel metal1 26496 28118 26496 28118 0 _0413_
rlabel metal2 10258 30158 10258 30158 0 _0414_
rlabel metal1 23092 16762 23092 16762 0 _0415_
rlabel metal2 22402 20638 22402 20638 0 _0416_
rlabel metal1 24150 17238 24150 17238 0 _0417_
rlabel metal2 25070 24990 25070 24990 0 _0418_
rlabel metal1 27370 27336 27370 27336 0 _0419_
rlabel metal1 21436 27098 21436 27098 0 _0420_
rlabel metal2 16698 25500 16698 25500 0 _0421_
rlabel metal1 26956 21590 26956 21590 0 _0422_
rlabel metal1 27968 17238 27968 17238 0 _0423_
rlabel metal1 27002 22746 27002 22746 0 _0424_
rlabel metal1 17296 4794 17296 4794 0 _0425_
rlabel metal3 21252 22984 21252 22984 0 _0426_
rlabel metal2 24058 17748 24058 17748 0 _0427_
rlabel metal1 13018 21590 13018 21590 0 _0428_
rlabel metal2 17802 17306 17802 17306 0 _0429_
rlabel metal1 21482 11322 21482 11322 0 _0430_
rlabel metal1 21896 10574 21896 10574 0 _0431_
rlabel metal1 21666 9146 21666 9146 0 _0432_
rlabel metal1 20240 5882 20240 5882 0 _0433_
rlabel metal1 6716 22678 6716 22678 0 _0434_
rlabel metal1 19964 7242 19964 7242 0 _0435_
rlabel via1 15398 21930 15398 21930 0 _0436_
rlabel metal3 23138 18836 23138 18836 0 _0437_
rlabel metal2 24978 18666 24978 18666 0 _0438_
rlabel metal1 27738 18666 27738 18666 0 _0439_
rlabel metal1 29808 13974 29808 13974 0 _0440_
rlabel metal2 20746 16915 20746 16915 0 _0441_
rlabel metal1 25576 9690 25576 9690 0 _0442_
rlabel metal2 26910 19074 26910 19074 0 _0443_
rlabel metal1 27186 13192 27186 13192 0 _0444_
rlabel metal1 25392 17850 25392 17850 0 _0445_
rlabel metal1 25990 13192 25990 13192 0 _0446_
rlabel metal1 23782 10778 23782 10778 0 _0447_
rlabel metal1 25990 14280 25990 14280 0 _0448_
rlabel metal1 18998 5270 18998 5270 0 _0449_
rlabel metal2 22402 5253 22402 5253 0 _0450_
rlabel metal1 28014 17306 28014 17306 0 _0451_
rlabel metal1 26772 14586 26772 14586 0 _0452_
rlabel metal1 30406 18394 30406 18394 0 _0453_
rlabel metal1 21482 19686 21482 19686 0 _0454_
rlabel metal2 27830 16286 27830 16286 0 _0455_
rlabel metal1 23414 14008 23414 14008 0 _0456_
rlabel metal1 22494 12886 22494 12886 0 _0457_
rlabel metal1 27186 11322 27186 11322 0 _0458_
rlabel metal1 24656 9622 24656 9622 0 _0459_
rlabel metal1 24794 14280 24794 14280 0 _0460_
rlabel metal1 21344 10098 21344 10098 0 _0461_
rlabel metal1 20663 14892 20663 14892 0 _0462_
rlabel metal2 23782 8517 23782 8517 0 _0463_
rlabel metal1 16698 15368 16698 15368 0 _0464_
rlabel metal1 21252 7446 21252 7446 0 _0465_
rlabel metal2 22678 9112 22678 9112 0 _0466_
rlabel metal1 5106 25942 5106 25942 0 _0467_
rlabel metal1 21206 18632 21206 18632 0 _0468_
rlabel metal1 16008 5338 16008 5338 0 _0469_
rlabel metal1 23552 14586 23552 14586 0 _0470_
rlabel metal1 19642 13192 19642 13192 0 _0471_
rlabel metal1 20976 13498 20976 13498 0 _0472_
rlabel metal1 7314 37230 7314 37230 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 38456 3502 38456 3502 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 8418 1367 8418 1367 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 29026 1078 29026 1078 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel via2 37490 17085 37490 17085 0 ccff_head
rlabel metal1 25346 37094 25346 37094 0 ccff_tail
rlabel metal1 2024 37230 2024 37230 0 chanx_left_in[0]
rlabel metal2 4094 20519 4094 20519 0 chanx_left_in[10]
rlabel metal2 36938 2907 36938 2907 0 chanx_left_in[11]
rlabel metal1 38088 36822 38088 36822 0 chanx_left_in[12]
rlabel metal1 3174 4182 3174 4182 0 chanx_left_in[13]
rlabel metal3 1142 22508 1142 22508 0 chanx_left_in[14]
rlabel metal2 18722 1588 18722 1588 0 chanx_left_in[15]
rlabel metal3 1878 39508 1878 39508 0 chanx_left_in[16]
rlabel metal2 38134 7123 38134 7123 0 chanx_left_in[17]
rlabel metal1 18216 37230 18216 37230 0 chanx_left_in[18]
rlabel via2 38134 30651 38134 30651 0 chanx_left_in[1]
rlabel metal3 1924 37468 1924 37468 0 chanx_left_in[2]
rlabel metal1 18538 36788 18538 36788 0 chanx_left_in[3]
rlabel metal1 22632 37298 22632 37298 0 chanx_left_in[4]
rlabel metal2 35466 1554 35466 1554 0 chanx_left_in[5]
rlabel metal1 37352 31790 37352 31790 0 chanx_left_in[6]
rlabel metal3 1786 38828 1786 38828 0 chanx_left_in[7]
rlabel metal1 9108 36754 9108 36754 0 chanx_left_in[8]
rlabel metal3 1188 15708 1188 15708 0 chanx_left_in[9]
rlabel via2 3450 24565 3450 24565 0 chanx_left_out[0]
rlabel metal2 38226 4301 38226 4301 0 chanx_left_out[10]
rlabel metal3 38786 38148 38786 38148 0 chanx_left_out[11]
rlabel metal1 4738 37094 4738 37094 0 chanx_left_out[12]
rlabel metal2 32246 1520 32246 1520 0 chanx_left_out[13]
rlabel via2 1794 7531 1794 7531 0 chanx_left_out[14]
rlabel metal2 33534 1520 33534 1520 0 chanx_left_out[15]
rlabel metal1 11776 2822 11776 2822 0 chanx_left_out[16]
rlabel metal3 1234 27948 1234 27948 0 chanx_left_out[17]
rlabel via2 38226 5525 38226 5525 0 chanx_left_out[18]
rlabel metal2 30958 1520 30958 1520 0 chanx_left_out[1]
rlabel metal3 1234 13668 1234 13668 0 chanx_left_out[2]
rlabel metal1 2852 37094 2852 37094 0 chanx_left_out[3]
rlabel metal1 1564 36890 1564 36890 0 chanx_left_out[4]
rlabel metal2 28382 1520 28382 1520 0 chanx_left_out[5]
rlabel metal1 36156 37094 36156 37094 0 chanx_left_out[6]
rlabel metal3 38740 25908 38740 25908 0 chanx_left_out[7]
rlabel metal1 24656 37094 24656 37094 0 chanx_left_out[8]
rlabel metal1 32154 37094 32154 37094 0 chanx_left_out[9]
rlabel metal2 4094 17204 4094 17204 0 chanx_right_in[0]
rlabel metal1 10442 3026 10442 3026 0 chanx_right_in[10]
rlabel metal1 36294 36142 36294 36142 0 chanx_right_in[11]
rlabel metal2 14858 1588 14858 1588 0 chanx_right_in[12]
rlabel metal2 24518 1588 24518 1588 0 chanx_right_in[13]
rlabel metal2 37490 32181 37490 32181 0 chanx_right_in[14]
rlabel metal2 38318 21913 38318 21913 0 chanx_right_in[15]
rlabel metal1 37168 37230 37168 37230 0 chanx_right_in[16]
rlabel via1 16606 37179 16606 37179 0 chanx_right_in[17]
rlabel via2 38318 19805 38318 19805 0 chanx_right_in[18]
rlabel metal2 10350 38260 10350 38260 0 chanx_right_in[1]
rlabel metal3 1188 5508 1188 5508 0 chanx_right_in[2]
rlabel metal1 14030 37230 14030 37230 0 chanx_right_in[3]
rlabel metal2 37490 27353 37490 27353 0 chanx_right_in[4]
rlabel metal2 26450 1554 26450 1554 0 chanx_right_in[5]
rlabel metal1 34546 37298 34546 37298 0 chanx_right_in[6]
rlabel metal1 38134 35734 38134 35734 0 chanx_right_in[7]
rlabel metal1 14904 37298 14904 37298 0 chanx_right_in[8]
rlabel metal2 17434 1588 17434 1588 0 chanx_right_in[9]
rlabel metal3 38740 12308 38740 12308 0 chanx_right_out[0]
rlabel metal3 38234 2108 38234 2108 0 chanx_right_out[10]
rlabel metal2 23506 37060 23506 37060 0 chanx_right_out[11]
rlabel via2 38226 35445 38226 35445 0 chanx_right_out[12]
rlabel metal2 38226 14297 38226 14297 0 chanx_right_out[13]
rlabel metal1 24012 2822 24012 2822 0 chanx_right_out[14]
rlabel metal3 2108 748 2108 748 0 chanx_right_out[15]
rlabel metal1 27876 37094 27876 37094 0 chanx_right_out[16]
rlabel metal2 38226 36057 38226 36057 0 chanx_right_out[17]
rlabel metal1 11500 36890 11500 36890 0 chanx_right_out[18]
rlabel metal2 38226 24837 38226 24837 0 chanx_right_out[1]
rlabel metal2 1334 1792 1334 1792 0 chanx_right_out[2]
rlabel metal2 12282 1520 12282 1520 0 chanx_right_out[3]
rlabel metal2 1794 30379 1794 30379 0 chanx_right_out[4]
rlabel metal1 32752 37434 32752 37434 0 chanx_right_out[5]
rlabel metal1 4232 10234 4232 10234 0 chanx_right_out[6]
rlabel metal2 36754 1520 36754 1520 0 chanx_right_out[7]
rlabel metal3 1234 32028 1234 32028 0 chanx_right_out[8]
rlabel metal2 4002 3247 4002 3247 0 chanx_right_out[9]
rlabel metal2 38134 16439 38134 16439 0 chany_bottom_in[0]
rlabel metal1 37352 10030 37352 10030 0 chany_bottom_in[10]
rlabel metal3 2200 29988 2200 29988 0 chany_bottom_in[11]
rlabel metal1 15594 36822 15594 36822 0 chany_bottom_in[12]
rlabel metal2 30314 1027 30314 1027 0 chany_bottom_in[13]
rlabel metal2 38134 33439 38134 33439 0 chany_bottom_in[14]
rlabel metal2 12926 976 12926 976 0 chany_bottom_in[15]
rlabel metal3 1142 35428 1142 35428 0 chany_bottom_in[16]
rlabel metal1 37352 29070 37352 29070 0 chany_bottom_in[17]
rlabel metal3 38280 68 38280 68 0 chany_bottom_in[18]
rlabel metal2 38134 10455 38134 10455 0 chany_bottom_in[1]
rlabel metal1 966 33490 966 33490 0 chany_bottom_in[2]
rlabel metal2 38318 18581 38318 18581 0 chany_bottom_in[3]
rlabel metal2 37398 1588 37398 1588 0 chany_bottom_in[4]
rlabel metal2 20010 1588 20010 1588 0 chany_bottom_in[5]
rlabel metal2 38134 21335 38134 21335 0 chany_bottom_in[6]
rlabel metal1 14950 16728 14950 16728 0 chany_bottom_in[7]
rlabel metal2 3910 12087 3910 12087 0 chany_bottom_in[8]
rlabel metal2 20654 38260 20654 38260 0 chany_bottom_in[9]
rlabel metal1 4094 20774 4094 20774 0 chany_bottom_out[0]
rlabel metal2 1794 36567 1794 36567 0 chany_bottom_out[10]
rlabel metal2 37490 36567 37490 36567 0 chany_bottom_out[11]
rlabel metal3 3580 1428 3580 1428 0 chany_bottom_out[12]
rlabel metal1 22172 36890 22172 36890 0 chany_bottom_out[13]
rlabel metal2 1794 17867 1794 17867 0 chany_bottom_out[14]
rlabel metal1 26910 37094 26910 37094 0 chany_bottom_out[15]
rlabel metal2 690 2064 690 2064 0 chany_bottom_out[16]
rlabel metal2 5842 1520 5842 1520 0 chany_bottom_out[17]
rlabel metal2 38226 4913 38226 4913 0 chany_bottom_out[18]
rlabel metal1 16928 2822 16928 2822 0 chany_bottom_out[1]
rlabel metal1 8878 37094 8878 37094 0 chany_bottom_out[2]
rlabel metal1 11776 37094 11776 37094 0 chany_bottom_out[3]
rlabel metal1 29808 37094 29808 37094 0 chany_bottom_out[4]
rlabel metal2 3910 1520 3910 1520 0 chany_bottom_out[5]
rlabel metal2 38226 8857 38226 8857 0 chany_bottom_out[6]
rlabel via2 38226 22491 38226 22491 0 chany_bottom_out[7]
rlabel metal1 13064 37094 13064 37094 0 chany_bottom_out[8]
rlabel metal2 38226 15181 38226 15181 0 chany_bottom_out[9]
rlabel metal1 4002 36822 4002 36822 0 chany_top_in[0]
rlabel metal2 21298 1554 21298 1554 0 chany_top_in[10]
rlabel metal2 38318 29461 38318 29461 0 chany_top_in[11]
rlabel metal2 30958 38260 30958 38260 0 chany_top_in[12]
rlabel metal2 9706 1588 9706 1588 0 chany_top_in[13]
rlabel via2 37490 11645 37490 11645 0 chany_top_in[14]
rlabel metal2 25806 1588 25806 1588 0 chany_top_in[15]
rlabel metal3 38786 748 38786 748 0 chany_top_in[16]
rlabel metal1 6256 37230 6256 37230 0 chany_top_in[17]
rlabel metal1 33028 3026 33028 3026 0 chany_top_in[18]
rlabel metal2 5198 1027 5198 1027 0 chany_top_in[1]
rlabel metal2 16146 1894 16146 1894 0 chany_top_in[2]
rlabel metal2 16698 12852 16698 12852 0 chany_top_in[3]
rlabel metal1 37352 34510 37352 34510 0 chany_top_in[4]
rlabel metal2 37490 24021 37490 24021 0 chany_top_in[5]
rlabel metal2 34822 1554 34822 1554 0 chany_top_in[6]
rlabel metal3 146 19788 146 19788 0 chany_top_in[7]
rlabel metal2 38318 13787 38318 13787 0 chany_top_in[8]
rlabel metal3 1119 25908 1119 25908 0 chany_top_in[9]
rlabel metal2 3818 13345 3818 13345 0 chany_top_out[0]
rlabel metal2 36846 37859 36846 37859 0 chany_top_out[10]
rlabel metal1 38134 2822 38134 2822 0 chany_top_out[11]
rlabel metal1 37398 36618 37398 36618 0 chany_top_out[12]
rlabel metal3 1234 27268 1234 27268 0 chany_top_out[13]
rlabel metal3 1234 29308 1234 29308 0 chany_top_out[14]
rlabel metal2 23230 1520 23230 1520 0 chany_top_out[15]
rlabel metal2 46 1044 46 1044 0 chany_top_out[16]
rlabel metal2 3818 4097 3818 4097 0 chany_top_out[17]
rlabel metal3 1234 32708 1234 32708 0 chany_top_out[18]
rlabel metal2 4002 4301 4002 4301 0 chany_top_out[1]
rlabel metal1 20056 37094 20056 37094 0 chany_top_out[2]
rlabel metal3 1234 25228 1234 25228 0 chany_top_out[3]
rlabel metal2 7130 1520 7130 1520 0 chany_top_out[4]
rlabel metal2 2622 1860 2622 1860 0 chany_top_out[5]
rlabel via2 3726 6171 3726 6171 0 chany_top_out[6]
rlabel metal1 19504 36890 19504 36890 0 chany_top_out[7]
rlabel metal2 19366 1520 19366 1520 0 chany_top_out[8]
rlabel metal1 33764 37094 33764 37094 0 chany_top_out[9]
rlabel metal1 14996 14246 14996 14246 0 clknet_0_prog_clk
rlabel metal1 1656 6834 1656 6834 0 clknet_4_0_0_prog_clk
rlabel metal1 2714 21556 2714 21556 0 clknet_4_10_0_prog_clk
rlabel metal1 1794 22542 1794 22542 0 clknet_4_11_0_prog_clk
rlabel metal2 6578 17680 6578 17680 0 clknet_4_12_0_prog_clk
rlabel metal2 9384 17646 9384 17646 0 clknet_4_13_0_prog_clk
rlabel metal1 7176 20434 7176 20434 0 clknet_4_14_0_prog_clk
rlabel metal1 7682 22678 7682 22678 0 clknet_4_15_0_prog_clk
rlabel metal2 6900 8942 6900 8942 0 clknet_4_1_0_prog_clk
rlabel metal2 2530 13600 2530 13600 0 clknet_4_2_0_prog_clk
rlabel metal1 6256 12750 6256 12750 0 clknet_4_3_0_prog_clk
rlabel metal2 9154 8942 9154 8942 0 clknet_4_4_0_prog_clk
rlabel metal1 14122 7854 14122 7854 0 clknet_4_5_0_prog_clk
rlabel metal1 9200 13294 9200 13294 0 clknet_4_6_0_prog_clk
rlabel metal2 11270 12614 11270 12614 0 clknet_4_7_0_prog_clk
rlabel metal2 2346 17442 2346 17442 0 clknet_4_8_0_prog_clk
rlabel metal1 7406 17714 7406 17714 0 clknet_4_9_0_prog_clk
rlabel metal2 38318 7701 38318 7701 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal3 1234 34068 1234 34068 0 left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal3 1717 8908 1717 8908 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 7774 2064 7774 2064 0 left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 11868 17646 11868 17646 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal1 13156 19754 13156 19754 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 23368 7854 23368 7854 0 mem_bottom_track_1.DFFR_1_.Q
rlabel via2 2346 6341 2346 6341 0 mem_bottom_track_1.DFFR_2_.Q
rlabel metal1 23828 13294 23828 13294 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal2 17986 20519 17986 20519 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 3404 5882 3404 5882 0 mem_bottom_track_1.DFFR_5_.Q
rlabel via2 3266 10115 3266 10115 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal1 2024 15062 2024 15062 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal1 9154 17782 9154 17782 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal2 12466 17969 12466 17969 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal3 17204 22780 17204 22780 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal2 6026 15827 6026 15827 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal1 5796 17714 5796 17714 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal1 3496 22066 3496 22066 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal1 2431 20026 2431 20026 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal1 4876 24106 4876 24106 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal1 6578 24242 6578 24242 0 mem_bottom_track_17.DFFR_7_.Q
rlabel metal2 9522 19550 9522 19550 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 10856 17102 10856 17102 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 20654 19720 20654 19720 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal2 13340 13124 13340 13124 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal1 29532 15470 29532 15470 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal2 18906 6596 18906 6596 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal2 20746 5032 20746 5032 0 mem_bottom_track_25.DFFR_6_.Q
rlabel metal1 7682 7446 7682 7446 0 mem_bottom_track_25.DFFR_7_.Q
rlabel metal1 10120 7378 10120 7378 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 13110 11118 13110 11118 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal2 21666 19737 21666 19737 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal2 23046 9962 23046 9962 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal3 12972 5440 12972 5440 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal2 17986 6800 17986 6800 0 mem_bottom_track_33.DFFR_5_.Q
rlabel metal2 17710 25823 17710 25823 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal3 10741 17884 10741 17884 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal2 29026 19567 29026 19567 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal1 16054 24208 16054 24208 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal1 14996 21522 14996 21522 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal1 10810 18598 10810 18598 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal1 11960 18870 11960 18870 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal1 12466 6732 12466 6732 0 mem_left_track_1.DFFR_0_.Q
rlabel metal4 17756 10948 17756 10948 0 mem_left_track_1.DFFR_1_.Q
rlabel metal1 6946 10744 6946 10744 0 mem_left_track_1.DFFR_2_.Q
rlabel metal1 8510 10642 8510 10642 0 mem_left_track_1.DFFR_3_.Q
rlabel metal1 4646 5746 4646 5746 0 mem_left_track_1.DFFR_4_.Q
rlabel metal1 5106 2618 5106 2618 0 mem_left_track_1.DFFR_5_.Q
rlabel metal1 3266 2618 3266 2618 0 mem_left_track_1.DFFR_6_.Q
rlabel metal1 1656 9622 1656 9622 0 mem_left_track_1.DFFR_7_.Q
rlabel metal1 1886 15368 1886 15368 0 mem_left_track_17.DFFR_0_.D
rlabel metal1 1702 12886 1702 12886 0 mem_left_track_17.DFFR_0_.Q
rlabel metal1 15686 18938 15686 18938 0 mem_left_track_17.DFFR_1_.Q
rlabel metal2 13110 27489 13110 27489 0 mem_left_track_17.DFFR_2_.Q
rlabel metal1 6440 13226 6440 13226 0 mem_left_track_17.DFFR_3_.Q
rlabel metal1 5290 9486 5290 9486 0 mem_left_track_17.DFFR_4_.Q
rlabel metal2 13202 24786 13202 24786 0 mem_left_track_17.DFFR_5_.Q
rlabel metal1 7084 21522 7084 21522 0 mem_left_track_17.DFFR_6_.Q
rlabel metal2 14214 25398 14214 25398 0 mem_left_track_17.DFFR_7_.Q
rlabel metal2 26450 20706 26450 20706 0 mem_left_track_25.DFFR_0_.Q
rlabel metal1 13616 20502 13616 20502 0 mem_left_track_25.DFFR_1_.Q
rlabel metal2 22862 21233 22862 21233 0 mem_left_track_25.DFFR_2_.Q
rlabel metal1 13294 22066 13294 22066 0 mem_left_track_25.DFFR_3_.Q
rlabel metal1 8648 24378 8648 24378 0 mem_left_track_25.DFFR_4_.Q
rlabel metal1 4830 23630 4830 23630 0 mem_left_track_25.DFFR_5_.Q
rlabel metal1 8004 24854 8004 24854 0 mem_left_track_25.DFFR_6_.Q
rlabel metal1 4646 15878 4646 15878 0 mem_left_track_25.DFFR_7_.Q
rlabel metal1 3450 13838 3450 13838 0 mem_left_track_33.DFFR_0_.Q
rlabel metal3 17204 8024 17204 8024 0 mem_left_track_33.DFFR_1_.Q
rlabel metal2 25576 18802 25576 18802 0 mem_left_track_33.DFFR_2_.Q
rlabel metal2 9246 8160 9246 8160 0 mem_left_track_33.DFFR_3_.Q
rlabel metal1 16928 8058 16928 8058 0 mem_left_track_33.DFFR_4_.Q
rlabel metal3 8671 19788 8671 19788 0 mem_left_track_9.DFFR_0_.Q
rlabel metal2 13662 15844 13662 15844 0 mem_left_track_9.DFFR_1_.Q
rlabel metal2 13754 15589 13754 15589 0 mem_left_track_9.DFFR_2_.Q
rlabel metal1 23690 19822 23690 19822 0 mem_left_track_9.DFFR_3_.Q
rlabel metal2 1702 11475 1702 11475 0 mem_left_track_9.DFFR_4_.Q
rlabel metal1 3358 16422 3358 16422 0 mem_left_track_9.DFFR_5_.Q
rlabel metal1 3128 14246 3128 14246 0 mem_left_track_9.DFFR_6_.Q
rlabel metal2 17250 1768 17250 1768 0 mem_right_track_0.DFFR_0_.D
rlabel metal2 6854 13719 6854 13719 0 mem_right_track_0.DFFR_0_.Q
rlabel metal2 11500 9180 11500 9180 0 mem_right_track_0.DFFR_1_.Q
rlabel metal1 9430 8568 9430 8568 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 27186 9520 27186 9520 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 15962 7174 15962 7174 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 8970 8330 8970 8330 0 mem_right_track_0.DFFR_5_.Q
rlabel metal1 11408 7990 11408 7990 0 mem_right_track_0.DFFR_6_.Q
rlabel metal3 11983 9044 11983 9044 0 mem_right_track_0.DFFR_7_.Q
rlabel metal1 4876 29138 4876 29138 0 mem_right_track_16.DFFR_0_.D
rlabel metal1 1840 23018 1840 23018 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 3358 21624 3358 21624 0 mem_right_track_16.DFFR_1_.Q
rlabel metal1 4876 21658 4876 21658 0 mem_right_track_16.DFFR_2_.Q
rlabel metal2 12558 28577 12558 28577 0 mem_right_track_16.DFFR_3_.Q
rlabel metal2 1978 23647 1978 23647 0 mem_right_track_16.DFFR_4_.Q
rlabel metal2 2530 21811 2530 21811 0 mem_right_track_16.DFFR_5_.Q
rlabel metal1 6210 19686 6210 19686 0 mem_right_track_16.DFFR_6_.Q
rlabel metal1 5704 15538 5704 15538 0 mem_right_track_16.DFFR_7_.Q
rlabel metal2 26818 18428 26818 18428 0 mem_right_track_24.DFFR_0_.Q
rlabel metal2 12926 18989 12926 18989 0 mem_right_track_24.DFFR_1_.Q
rlabel metal3 17020 14824 17020 14824 0 mem_right_track_24.DFFR_2_.Q
rlabel metal1 14444 15062 14444 15062 0 mem_right_track_24.DFFR_3_.Q
rlabel metal1 14352 24650 14352 24650 0 mem_right_track_24.DFFR_4_.Q
rlabel metal2 21850 23579 21850 23579 0 mem_right_track_24.DFFR_5_.Q
rlabel metal1 13156 22950 13156 22950 0 mem_right_track_24.DFFR_6_.Q
rlabel metal3 11500 17884 11500 17884 0 mem_right_track_24.DFFR_7_.Q
rlabel metal1 28336 13294 28336 13294 0 mem_right_track_32.DFFR_0_.Q
rlabel metal1 11178 10540 11178 10540 0 mem_right_track_32.DFFR_1_.Q
rlabel metal1 29854 13294 29854 13294 0 mem_right_track_32.DFFR_2_.Q
rlabel metal2 11178 9469 11178 9469 0 mem_right_track_32.DFFR_3_.Q
rlabel metal2 13294 15793 13294 15793 0 mem_right_track_32.DFFR_4_.Q
rlabel metal3 13064 21964 13064 21964 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 2438 17034 2438 17034 0 mem_right_track_8.DFFR_1_.Q
rlabel metal2 14122 17544 14122 17544 0 mem_right_track_8.DFFR_2_.Q
rlabel metal3 19412 18564 19412 18564 0 mem_right_track_8.DFFR_3_.Q
rlabel metal1 2714 18938 2714 18938 0 mem_right_track_8.DFFR_4_.Q
rlabel metal2 2162 23290 2162 23290 0 mem_right_track_8.DFFR_5_.Q
rlabel metal1 3450 22474 3450 22474 0 mem_right_track_8.DFFR_6_.Q
rlabel metal1 8602 14280 8602 14280 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 10718 17578 10718 17578 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 13662 19822 13662 19822 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 13754 23222 13754 23222 0 mem_top_track_0.DFFR_3_.Q
rlabel metal1 1932 10710 1932 10710 0 mem_top_track_0.DFFR_4_.Q
rlabel metal2 3910 6511 3910 6511 0 mem_top_track_0.DFFR_5_.Q
rlabel metal1 1978 13192 1978 13192 0 mem_top_track_0.DFFR_6_.Q
rlabel metal2 2714 29359 2714 29359 0 mem_top_track_0.DFFR_7_.Q
rlabel metal1 20792 4590 20792 4590 0 mem_top_track_16.DFFR_0_.D
rlabel metal2 5520 2652 5520 2652 0 mem_top_track_16.DFFR_0_.Q
rlabel via3 5451 12852 5451 12852 0 mem_top_track_16.DFFR_1_.Q
rlabel metal3 17503 18020 17503 18020 0 mem_top_track_16.DFFR_2_.Q
rlabel metal2 3818 17204 3818 17204 0 mem_top_track_16.DFFR_3_.Q
rlabel metal2 16698 3451 16698 3451 0 mem_top_track_16.DFFR_4_.Q
rlabel metal1 6302 5338 6302 5338 0 mem_top_track_16.DFFR_5_.Q
rlabel metal2 16882 5984 16882 5984 0 mem_top_track_16.DFFR_6_.Q
rlabel metal2 15410 6222 15410 6222 0 mem_top_track_16.DFFR_7_.Q
rlabel metal1 24518 21522 24518 21522 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 12650 15011 12650 15011 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 27922 13906 27922 13906 0 mem_top_track_24.DFFR_2_.Q
rlabel metal3 20332 19040 20332 19040 0 mem_top_track_24.DFFR_3_.Q
rlabel metal1 8510 17034 8510 17034 0 mem_top_track_24.DFFR_4_.Q
rlabel metal1 11178 18054 11178 18054 0 mem_top_track_24.DFFR_5_.Q
rlabel metal1 11270 15674 11270 15674 0 mem_top_track_24.DFFR_6_.Q
rlabel metal1 19642 22474 19642 22474 0 mem_top_track_24.DFFR_7_.Q
rlabel metal2 13938 26044 13938 26044 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 9384 13838 9384 13838 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 2300 5270 2300 5270 0 mem_top_track_32.DFFR_2_.Q
rlabel metal1 1886 3128 1886 3128 0 mem_top_track_32.DFFR_3_.Q
rlabel metal2 12742 3672 12742 3672 0 mem_top_track_32.DFFR_4_.Q
rlabel metal1 17342 30294 17342 30294 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 18216 24786 18216 24786 0 mem_top_track_8.DFFR_1_.Q
rlabel metal1 18492 31246 18492 31246 0 mem_top_track_8.DFFR_2_.Q
rlabel metal1 21482 24684 21482 24684 0 mem_top_track_8.DFFR_3_.Q
rlabel metal3 8878 19516 8878 19516 0 mem_top_track_8.DFFR_4_.Q
rlabel metal4 20700 19924 20700 19924 0 mem_top_track_8.DFFR_5_.Q
rlabel metal1 2024 4658 2024 4658 0 mem_top_track_8.DFFR_6_.Q
rlabel metal1 15410 18190 15410 18190 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 7130 32742 7130 32742 0 mux_bottom_track_1.INVTX1_10_.out
rlabel metal1 19826 5066 19826 5066 0 mux_bottom_track_1.INVTX1_11_.out
rlabel metal1 18216 12750 18216 12750 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal1 17802 8874 17802 8874 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 18446 22678 18446 22678 0 mux_bottom_track_1.INVTX1_3_.out
rlabel metal2 27094 24089 27094 24089 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal1 15042 9418 15042 9418 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal2 16974 16133 16974 16133 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal2 16238 5185 16238 5185 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal1 18032 28390 18032 28390 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal1 29923 22474 29923 22474 0 mux_bottom_track_1.INVTX1_9_.out
rlabel metal1 14306 18190 14306 18190 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 17802 15776 17802 15776 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 19090 21352 19090 21352 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 1978 25092 1978 25092 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 2024 32946 2024 32946 0 mux_bottom_track_1.out
rlabel metal1 14582 28186 14582 28186 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal2 19550 4063 19550 4063 0 mux_bottom_track_17.INVTX1_10_.out
rlabel metal1 9338 26894 9338 26894 0 mux_bottom_track_17.INVTX1_11_.out
rlabel via2 15410 21675 15410 21675 0 mux_bottom_track_17.INVTX1_1_.out
rlabel via2 14490 10693 14490 10693 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 5290 21454 5290 21454 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 25484 33354 25484 33354 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 15962 19754 15962 19754 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal2 16146 27642 16146 27642 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal2 10534 32028 10534 32028 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal1 9154 26282 9154 26282 0 mux_bottom_track_17.INVTX1_8_.out
rlabel metal1 7912 20978 7912 20978 0 mux_bottom_track_17.INVTX1_9_.out
rlabel metal2 9246 20723 9246 20723 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 19550 27948 19550 27948 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 8740 20842 8740 20842 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 11684 33966 11684 33966 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 11408 34170 11408 34170 0 mux_bottom_track_17.out
rlabel metal2 27278 26010 27278 26010 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal1 28612 21454 28612 21454 0 mux_bottom_track_25.INVTX1_10_.out
rlabel metal1 18722 31790 18722 31790 0 mux_bottom_track_25.INVTX1_11_.out
rlabel metal1 26588 24718 26588 24718 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal1 21482 27506 21482 27506 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal1 17894 21590 17894 21590 0 mux_bottom_track_25.INVTX1_3_.out
rlabel metal1 26772 17102 26772 17102 0 mux_bottom_track_25.INVTX1_4_.out
rlabel metal1 25208 13838 25208 13838 0 mux_bottom_track_25.INVTX1_5_.out
rlabel metal1 22402 18802 22402 18802 0 mux_bottom_track_25.INVTX1_6_.out
rlabel metal1 29486 12682 29486 12682 0 mux_bottom_track_25.INVTX1_7_.out
rlabel metal1 26266 20978 26266 20978 0 mux_bottom_track_25.INVTX1_8_.out
rlabel metal2 22494 19890 22494 19890 0 mux_bottom_track_25.INVTX1_9_.out
rlabel metal1 15226 13158 15226 13158 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 23138 14484 23138 14484 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 23966 27982 23966 27982 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 21666 4114 21666 4114 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 20286 4080 20286 4080 0 mux_bottom_track_25.out
rlabel metal2 25898 14399 25898 14399 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal1 24426 17850 24426 17850 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal2 16606 12716 16606 12716 0 mux_bottom_track_33.INVTX1_2_.out
rlabel metal1 21459 7310 21459 7310 0 mux_bottom_track_33.INVTX1_3_.out
rlabel metal2 29946 19618 29946 19618 0 mux_bottom_track_33.INVTX1_4_.out
rlabel metal2 20424 28628 20424 28628 0 mux_bottom_track_33.INVTX1_5_.out
rlabel metal1 23460 12682 23460 12682 0 mux_bottom_track_33.INVTX1_6_.out
rlabel metal2 29118 19244 29118 19244 0 mux_bottom_track_33.INVTX1_7_.out
rlabel metal1 25392 14382 25392 14382 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal3 24633 18292 24633 18292 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 25714 11662 25714 11662 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 19297 7990 19297 7990 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 20194 3026 20194 3026 0 mux_bottom_track_33.out
rlabel metal1 16974 16626 16974 16626 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 29762 17102 29762 17102 0 mux_bottom_track_9.INVTX1_10_.out
rlabel metal1 14812 27370 14812 27370 0 mux_bottom_track_9.INVTX1_11_.out
rlabel metal1 27922 16116 27922 16116 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 24380 20230 24380 20230 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 20102 22066 20102 22066 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal2 21390 30532 21390 30532 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal1 27600 32742 27600 32742 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal2 24702 23596 24702 23596 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal1 28612 16014 28612 16014 0 mux_bottom_track_9.INVTX1_7_.out
rlabel metal1 20516 27506 20516 27506 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal1 13202 26418 13202 26418 0 mux_bottom_track_9.INVTX1_9_.out
rlabel metal1 25898 16490 25898 16490 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 21942 21420 21942 21420 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 17526 25024 17526 25024 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 25438 29036 25438 29036 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 27002 29818 27002 29818 0 mux_bottom_track_9.out
rlabel metal1 24702 7752 24702 7752 0 mux_left_track_1.INVTX1_10_.out
rlabel metal2 20746 4318 20746 4318 0 mux_left_track_1.INVTX1_11_.out
rlabel metal2 20838 5185 20838 5185 0 mux_left_track_1.INVTX1_1_.out
rlabel metal2 20378 13940 20378 13940 0 mux_left_track_1.INVTX1_7_.out
rlabel metal1 23506 15062 23506 15062 0 mux_left_track_1.INVTX1_8_.out
rlabel metal1 21896 13362 21896 13362 0 mux_left_track_1.INVTX1_9_.out
rlabel metal1 6072 19210 6072 19210 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 20516 17578 20516 17578 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 17986 7225 17986 7225 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 4830 31926 4830 31926 0 mux_left_track_1.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 1886 31824 1886 31824 0 mux_left_track_1.out
rlabel metal1 6348 29070 6348 29070 0 mux_left_track_17.INVTX1_10_.out
rlabel via2 30406 12971 30406 12971 0 mux_left_track_17.INVTX1_11_.out
rlabel metal2 27094 12920 27094 12920 0 mux_left_track_17.INVTX1_2_.out
rlabel metal2 9522 9996 9522 9996 0 mux_left_track_17.INVTX1_7_.out
rlabel metal1 4048 30158 4048 30158 0 mux_left_track_17.INVTX1_8_.out
rlabel metal2 18906 29376 18906 29376 0 mux_left_track_17.INVTX1_9_.out
rlabel metal3 15778 19516 15778 19516 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 6854 21199 6854 21199 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 19550 24684 19550 24684 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 22402 33966 22402 33966 0 mux_left_track_17.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 23690 33660 23690 33660 0 mux_left_track_17.out
rlabel metal2 25990 21862 25990 21862 0 mux_left_track_25.INVTX1_10_.out
rlabel metal1 8556 29070 8556 29070 0 mux_left_track_25.INVTX1_11_.out
rlabel metal2 32062 27642 32062 27642 0 mux_left_track_25.INVTX1_2_.out
rlabel metal2 28382 16150 28382 16150 0 mux_left_track_25.INVTX1_7_.out
rlabel metal1 29670 16150 29670 16150 0 mux_left_track_25.INVTX1_8_.out
rlabel metal2 12742 29954 12742 29954 0 mux_left_track_25.INVTX1_9_.out
rlabel metal2 21390 27149 21390 27149 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 16146 17748 16146 17748 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 27048 27982 27048 27982 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 13110 30702 13110 30702 0 mux_left_track_25.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 10810 36142 10810 36142 0 mux_left_track_25.out
rlabel metal1 2254 18190 2254 18190 0 mux_left_track_33.INVTX1_1_.out
rlabel metal1 21666 6222 21666 6222 0 mux_left_track_33.INVTX1_5_.out
rlabel metal1 19642 18360 19642 18360 0 mux_left_track_33.INVTX1_6_.out
rlabel metal2 22770 7072 22770 7072 0 mux_left_track_33.INVTX1_7_.out
rlabel metal2 16514 14212 16514 14212 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 21390 7667 21390 7667 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 17112 12886 17112 12886 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal3 18377 6732 18377 6732 0 mux_left_track_33.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 18354 3468 18354 3468 0 mux_left_track_33.out
rlabel metal1 22172 25330 22172 25330 0 mux_left_track_9.INVTX1_10_.out
rlabel metal1 18676 3706 18676 3706 0 mux_left_track_9.INVTX1_11_.out
rlabel metal2 27278 7854 27278 7854 0 mux_left_track_9.INVTX1_3_.out
rlabel metal1 20148 23154 20148 23154 0 mux_left_track_9.INVTX1_7_.out
rlabel metal2 29854 17680 29854 17680 0 mux_left_track_9.INVTX1_8_.out
rlabel metal1 16376 22542 16376 22542 0 mux_left_track_9.INVTX1_9_.out
rlabel metal1 26818 19414 26818 19414 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 17526 24106 17526 24106 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 14306 17816 14306 17816 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 5474 36720 5474 36720 0 mux_left_track_9.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 5566 36346 5566 36346 0 mux_left_track_9.out
rlabel metal1 28612 32198 28612 32198 0 mux_right_track_0.INVTX1_4_.out
rlabel metal2 16560 15538 16560 15538 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 28198 16439 28198 16439 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 20562 19040 20562 19040 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 33994 11696 33994 11696 0 mux_right_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 34086 12036 34086 12036 0 mux_right_track_0.out
rlabel metal2 30774 27506 30774 27506 0 mux_right_track_16.INVTX1_4_.out
rlabel metal1 5290 19754 5290 19754 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 5934 25296 5934 25296 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 4094 26452 4094 26452 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 6256 28118 6256 28118 0 mux_right_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 6578 31110 6578 31110 0 mux_right_track_16.out
rlabel metal1 25024 7446 25024 7446 0 mux_right_track_24.INVTX1_4_.out
rlabel metal1 28428 25942 28428 25942 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 29210 13940 29210 13940 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 25300 22066 25300 22066 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 30866 24752 30866 24752 0 mux_right_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 34822 31790 34822 31790 0 mux_right_track_24.out
rlabel metal1 25346 18190 25346 18190 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 25208 10574 25208 10574 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 28198 18632 28198 18632 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 26174 28492 26174 28492 0 mux_right_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 27324 33966 27324 33966 0 mux_right_track_32.out
rlabel metal1 24150 33898 24150 33898 0 mux_right_track_8.INVTX1_4_.out
rlabel metal1 18722 16490 18722 16490 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 12466 26962 12466 26962 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 21390 25534 21390 25534 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 12880 21454 12880 21454 0 mux_right_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 5428 30226 5428 30226 0 mux_right_track_8.out
rlabel metal1 6785 34510 6785 34510 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 22862 23018 22862 23018 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 14904 9622 14904 9622 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 17986 20842 17986 20842 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 21390 4607 21390 4607 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 24150 4284 24150 4284 0 mux_top_track_0.out
rlabel metal1 24656 6630 24656 6630 0 mux_top_track_16.INVTX1_0_.out
rlabel metal1 16882 13770 16882 13770 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 19826 25398 19826 25398 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal2 8418 26554 8418 26554 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 17618 5372 17618 5372 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 18768 2346 18768 2346 0 mux_top_track_16.out
rlabel metal1 23276 4182 23276 4182 0 mux_top_track_24.INVTX1_0_.out
rlabel metal1 24242 18156 24242 18156 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 30176 15606 30176 15606 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel via1 28842 19397 28842 19397 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 31878 34578 31878 34578 0 mux_top_track_24.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal1 35328 34578 35328 34578 0 mux_top_track_24.out
rlabel metal1 17710 12206 17710 12206 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 18400 17646 18400 17646 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 7314 22508 7314 22508 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 15824 23018 15824 23018 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 21022 3468 21022 3468 0 mux_top_track_32.out
rlabel metal1 12098 34918 12098 34918 0 mux_top_track_8.INVTX1_0_.out
rlabel metal2 15410 27200 15410 27200 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 22402 24752 22402 24752 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 15456 27370 15456 27370 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 14674 19414 14674 19414 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_3_out
rlabel metal2 21482 3230 21482 3230 0 mux_top_track_8.out
rlabel metal1 9062 37162 9062 37162 0 net1
rlabel metal1 20194 5202 20194 5202 0 net10
rlabel metal1 32338 2380 32338 2380 0 net100
rlabel metal2 20746 2618 20746 2618 0 net101
rlabel metal1 33810 21862 33810 21862 0 net102
rlabel metal1 18170 3128 18170 3128 0 net103
rlabel metal2 1610 28492 1610 28492 0 net104
rlabel metal1 37628 5882 37628 5882 0 net105
rlabel metal1 22218 2380 22218 2380 0 net106
rlabel metal2 1702 17204 1702 17204 0 net107
rlabel metal1 2852 37230 2852 37230 0 net108
rlabel metal1 3864 36346 3864 36346 0 net109
rlabel metal1 1932 21454 1932 21454 0 net11
rlabel metal1 29624 2074 29624 2074 0 net110
rlabel metal1 36156 37230 36156 37230 0 net111
rlabel metal1 38042 26384 38042 26384 0 net112
rlabel metal1 24058 33626 24058 33626 0 net113
rlabel metal1 25921 36618 25921 36618 0 net114
rlabel metal1 37260 12818 37260 12818 0 net115
rlabel metal2 38042 5134 38042 5134 0 net116
rlabel metal1 23368 36754 23368 36754 0 net117
rlabel metal1 38042 35632 38042 35632 0 net118
rlabel metal1 37812 19482 37812 19482 0 net119
rlabel metal2 19458 3366 19458 3366 0 net12
rlabel metal2 23966 3196 23966 3196 0 net120
rlabel metal2 10994 2431 10994 2431 0 net121
rlabel metal1 27738 37230 27738 37230 0 net122
rlabel metal1 23598 36618 23598 36618 0 net123
rlabel metal2 11730 35972 11730 35972 0 net124
rlabel via2 37674 25211 37674 25211 0 net125
rlabel metal2 16422 19040 16422 19040 0 net126
rlabel metal1 12374 2516 12374 2516 0 net127
rlabel metal1 1610 30192 1610 30192 0 net128
rlabel metal1 29210 36618 29210 36618 0 net129
rlabel metal2 3174 36380 3174 36380 0 net13
rlabel metal2 16054 9809 16054 9809 0 net130
rlabel metal1 37168 2482 37168 2482 0 net131
rlabel metal1 3312 32334 3312 32334 0 net132
rlabel metal4 6992 12420 6992 12420 0 net133
rlabel metal1 1748 33014 1748 33014 0 net134
rlabel metal1 2254 36074 2254 36074 0 net135
rlabel metal1 37306 36108 37306 36108 0 net136
rlabel metal1 20102 4012 20102 4012 0 net137
rlabel metal2 22402 36550 22402 36550 0 net138
rlabel metal1 1610 17136 1610 17136 0 net139
rlabel metal2 37536 11084 37536 11084 0 net14
rlabel metal1 26726 37230 26726 37230 0 net140
rlabel metal1 18906 2856 18906 2856 0 net141
rlabel metal1 6325 2414 6325 2414 0 net142
rlabel metal1 35236 5202 35236 5202 0 net143
rlabel metal1 17480 3026 17480 3026 0 net144
rlabel metal3 8855 36516 8855 36516 0 net145
rlabel metal2 16146 33762 16146 33762 0 net146
rlabel metal1 28704 34714 28704 34714 0 net147
rlabel via2 4646 2533 4646 2533 0 net148
rlabel metal1 37950 14790 37950 14790 0 net149
rlabel metal1 18078 37094 18078 37094 0 net15
rlabel metal1 36984 16218 36984 16218 0 net150
rlabel metal1 12374 35802 12374 35802 0 net151
rlabel metal2 37398 15028 37398 15028 0 net152
rlabel metal4 16100 6596 16100 6596 0 net153
rlabel metal1 36662 36720 36662 36720 0 net154
rlabel metal1 37812 3026 37812 3026 0 net155
rlabel metal2 35926 35734 35926 35734 0 net156
rlabel metal1 1610 27506 1610 27506 0 net157
rlabel metal1 1610 29682 1610 29682 0 net158
rlabel metal2 23322 2465 23322 2465 0 net159
rlabel metal2 38226 28798 38226 28798 0 net16
rlabel metal1 20838 2924 20838 2924 0 net160
rlabel via3 2093 30396 2093 30396 0 net161
rlabel metal2 2254 32640 2254 32640 0 net162
rlabel metal1 4646 4454 4646 4454 0 net163
rlabel metal1 20010 37230 20010 37230 0 net164
rlabel metal1 1610 26384 1610 26384 0 net165
rlabel metal2 10902 2601 10902 2601 0 net166
rlabel metal2 6578 2975 6578 2975 0 net167
rlabel metal2 23138 5950 23138 5950 0 net168
rlabel metal1 19964 31450 19964 31450 0 net169
rlabel metal1 6026 36890 6026 36890 0 net17
rlabel metal1 18032 2618 18032 2618 0 net170
rlabel metal1 23897 36074 23897 36074 0 net171
rlabel metal1 1840 24718 1840 24718 0 net172
rlabel metal1 18078 4590 18078 4590 0 net173
rlabel metal1 17158 3570 17158 3570 0 net174
rlabel metal2 27738 26656 27738 26656 0 net175
rlabel metal1 30866 12274 30866 12274 0 net176
rlabel metal1 7084 27982 7084 27982 0 net177
rlabel metal1 5566 27982 5566 27982 0 net178
rlabel metal2 30590 23902 30590 23902 0 net179
rlabel metal1 18538 36550 18538 36550 0 net18
rlabel metal2 12926 17629 12926 17629 0 net180
rlabel metal1 24564 29206 24564 29206 0 net181
rlabel metal2 11730 31212 11730 31212 0 net182
rlabel metal2 6578 1972 6578 1972 0 net183
rlabel via3 4899 19788 4899 19788 0 net184
rlabel metal1 8648 30294 8648 30294 0 net185
rlabel metal1 19182 30158 19182 30158 0 net186
rlabel metal2 12466 30464 12466 30464 0 net187
rlabel metal1 13340 21454 13340 21454 0 net188
rlabel metal1 29026 14008 29026 14008 0 net189
rlabel metal1 22954 37196 22954 37196 0 net19
rlabel metal1 27692 15130 27692 15130 0 net190
rlabel metal1 16560 14450 16560 14450 0 net191
rlabel metal1 36570 3638 36570 3638 0 net2
rlabel metal1 28290 2550 28290 2550 0 net20
rlabel metal2 37582 23698 37582 23698 0 net21
rlabel metal1 5428 37162 5428 37162 0 net22
rlabel metal2 9430 28900 9430 28900 0 net23
rlabel metal2 3726 15606 3726 15606 0 net24
rlabel metal3 6233 8092 6233 8092 0 net25
rlabel metal3 20148 3400 20148 3400 0 net26
rlabel metal2 36202 34442 36202 34442 0 net27
rlabel metal2 15226 1938 15226 1938 0 net28
rlabel metal1 23460 2482 23460 2482 0 net29
rlabel metal2 9154 2142 9154 2142 0 net3
rlabel metal1 33994 21998 33994 21998 0 net30
rlabel metal1 37007 21862 37007 21862 0 net31
rlabel metal2 37674 32470 37674 32470 0 net32
rlabel metal1 19918 37434 19918 37434 0 net33
rlabel metal2 31510 19516 31510 19516 0 net34
rlabel metal2 10626 34485 10626 34485 0 net35
rlabel metal1 1380 4114 1380 4114 0 net36
rlabel metal1 14674 37094 14674 37094 0 net37
rlabel metal1 37582 27506 37582 27506 0 net38
rlabel metal1 26312 2550 26312 2550 0 net39
rlabel metal1 29348 8466 29348 8466 0 net4
rlabel metal2 36570 31246 36570 31246 0 net40
rlabel metal2 34546 34476 34546 34476 0 net41
rlabel metal1 22402 36618 22402 36618 0 net42
rlabel metal2 31326 4420 31326 4420 0 net43
rlabel metal1 35880 16762 35880 16762 0 net44
rlabel metal2 37766 7854 37766 7854 0 net45
rlabel metal1 5106 32198 5106 32198 0 net46
rlabel metal1 13110 36618 13110 36618 0 net47
rlabel metal2 30406 2329 30406 2329 0 net48
rlabel metal1 37099 33354 37099 33354 0 net49
rlabel metal1 36823 17170 36823 17170 0 net5
rlabel metal2 24610 5508 24610 5508 0 net50
rlabel metal1 2024 35598 2024 35598 0 net51
rlabel metal1 37766 29036 37766 29036 0 net52
rlabel metal1 36294 3706 36294 3706 0 net53
rlabel metal1 20792 26962 20792 26962 0 net54
rlabel metal1 2530 33354 2530 33354 0 net55
rlabel metal2 34546 18122 34546 18122 0 net56
rlabel metal2 37766 2210 37766 2210 0 net57
rlabel metal1 20562 6290 20562 6290 0 net58
rlabel via2 38226 21675 38226 21675 0 net59
rlabel metal1 9476 37434 9476 37434 0 net6
rlabel metal2 5198 29512 5198 29512 0 net60
rlabel metal1 18814 24038 18814 24038 0 net61
rlabel metal2 20930 37026 20930 37026 0 net62
rlabel metal1 4830 36618 4830 36618 0 net63
rlabel metal1 23598 2550 23598 2550 0 net64
rlabel metal2 37030 29002 37030 29002 0 net65
rlabel metal1 23552 36142 23552 36142 0 net66
rlabel metal2 10074 2244 10074 2244 0 net67
rlabel metal1 37766 11628 37766 11628 0 net68
rlabel metal1 26036 2618 26036 2618 0 net69
rlabel metal1 24610 19788 24610 19788 0 net7
rlabel metal2 21896 3638 21896 3638 0 net70
rlabel metal2 20194 36623 20194 36623 0 net71
rlabel metal2 30406 4964 30406 4964 0 net72
rlabel metal2 5290 2601 5290 2601 0 net73
rlabel metal2 16330 3111 16330 3111 0 net74
rlabel metal1 23138 5202 23138 5202 0 net75
rlabel metal2 37766 30532 37766 30532 0 net76
rlabel metal1 37904 14994 37904 14994 0 net77
rlabel metal1 36018 16082 36018 16082 0 net78
rlabel metal1 3128 33286 3128 33286 0 net79
rlabel metal1 35604 3162 35604 3162 0 net8
rlabel metal1 37398 14382 37398 14382 0 net80
rlabel metal1 2438 32198 2438 32198 0 net81
rlabel metal1 33166 12818 33166 12818 0 net82
rlabel metal1 3726 34714 3726 34714 0 net83
rlabel metal1 22678 4624 22678 4624 0 net84
rlabel metal1 20102 3604 20102 3604 0 net85
rlabel metal2 19090 4165 19090 4165 0 net86
rlabel metal1 37007 26826 37007 26826 0 net87
rlabel metal2 22862 5304 22862 5304 0 net88
rlabel metal1 28842 36550 28842 36550 0 net89
rlabel metal1 38042 36550 38042 36550 0 net9
rlabel metal1 24702 33966 24702 33966 0 net90
rlabel metal1 3220 36006 3220 36006 0 net91
rlabel metal1 8648 36550 8648 36550 0 net92
rlabel metal1 26864 3162 26864 3162 0 net93
rlabel metal1 24564 3162 24564 3162 0 net94
rlabel metal2 25346 35173 25346 35173 0 net95
rlabel metal1 2760 31926 2760 31926 0 net96
rlabel metal1 34891 4590 34891 4590 0 net97
rlabel metal1 37674 35054 37674 35054 0 net98
rlabel metal2 5750 36788 5750 36788 0 net99
rlabel metal2 14214 2200 14214 2200 0 pReset
rlabel metal2 14306 13736 14306 13736 0 prog_clk
rlabel metal2 38318 26775 38318 26775 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 21942 1894 21942 1894 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal1 29164 36754 29164 36754 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 28842 37196 28842 37196 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal1 2530 36176 2530 36176 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 6624 36754 6624 36754 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_
rlabel metal1 27876 3026 27876 3026 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 2898 7701 2898 7701 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
