magic
tech sky130A
magscale 1 2
timestamp 1674174822
<< viali >>
rect 12541 37417 12575 37451
rect 17969 37417 18003 37451
rect 32505 37417 32539 37451
rect 13553 37349 13587 37383
rect 14565 37349 14599 37383
rect 28549 37349 28583 37383
rect 2053 37281 2087 37315
rect 4261 37281 4295 37315
rect 9137 37281 9171 37315
rect 23029 37281 23063 37315
rect 25789 37281 25823 37315
rect 30297 37281 30331 37315
rect 37473 37281 37507 37315
rect 2329 37213 2363 37247
rect 4077 37213 4111 37247
rect 5457 37213 5491 37247
rect 6745 37213 6779 37247
rect 7389 37213 7423 37247
rect 8585 37213 8619 37247
rect 9413 37213 9447 37247
rect 10425 37213 10459 37247
rect 11713 37213 11747 37247
rect 12449 37213 12483 37247
rect 13737 37213 13771 37247
rect 14381 37213 14415 37247
rect 15209 37213 15243 37247
rect 16037 37213 16071 37247
rect 16865 37213 16899 37247
rect 18153 37213 18187 37247
rect 18613 37213 18647 37247
rect 20085 37213 20119 37247
rect 22005 37213 22039 37247
rect 22845 37213 22879 37247
rect 23489 37213 23523 37247
rect 24777 37213 24811 37247
rect 26065 37213 26099 37247
rect 27169 37213 27203 37247
rect 28089 37213 28123 37247
rect 28733 37213 28767 37247
rect 30021 37213 30055 37247
rect 32321 37213 32355 37247
rect 33057 37213 33091 37247
rect 34897 37213 34931 37247
rect 36185 37213 36219 37247
rect 37749 37213 37783 37247
rect 5273 37077 5307 37111
rect 6561 37077 6595 37111
rect 7205 37077 7239 37111
rect 8401 37077 8435 37111
rect 10609 37077 10643 37111
rect 11805 37077 11839 37111
rect 15025 37077 15059 37111
rect 16221 37077 16255 37111
rect 17049 37077 17083 37111
rect 18797 37077 18831 37111
rect 20269 37077 20303 37111
rect 22201 37077 22235 37111
rect 23673 37077 23707 37111
rect 24593 37077 24627 37111
rect 27353 37077 27387 37111
rect 27905 37077 27939 37111
rect 31769 37077 31803 37111
rect 33241 37077 33275 37111
rect 35081 37077 35115 37111
rect 36369 37077 36403 37111
rect 3985 36873 4019 36907
rect 37657 36873 37691 36907
rect 1777 36805 1811 36839
rect 7481 36805 7515 36839
rect 11805 36805 11839 36839
rect 13645 36805 13679 36839
rect 17969 36805 18003 36839
rect 25053 36805 25087 36839
rect 30113 36805 30147 36839
rect 34437 36805 34471 36839
rect 36737 36805 36771 36839
rect 3341 36737 3375 36771
rect 4169 36737 4203 36771
rect 4813 36737 4847 36771
rect 7389 36737 7423 36771
rect 8217 36737 8251 36771
rect 8677 36737 8711 36771
rect 9321 36737 9355 36771
rect 9965 36737 9999 36771
rect 10609 36737 10643 36771
rect 12817 36737 12851 36771
rect 14841 36737 14875 36771
rect 15761 36737 15795 36771
rect 32505 36737 32539 36771
rect 33149 36737 33183 36771
rect 37473 36737 37507 36771
rect 1685 36669 1719 36703
rect 2697 36669 2731 36703
rect 13553 36669 13587 36703
rect 15853 36669 15887 36703
rect 17693 36669 17727 36703
rect 22569 36669 22603 36703
rect 22845 36669 22879 36703
rect 24777 36669 24811 36703
rect 27537 36669 27571 36703
rect 27813 36669 27847 36703
rect 29837 36669 29871 36703
rect 34161 36669 34195 36703
rect 4905 36601 4939 36635
rect 8033 36601 8067 36635
rect 8769 36601 8803 36635
rect 14105 36601 14139 36635
rect 14657 36601 14691 36635
rect 26525 36601 26559 36635
rect 29285 36601 29319 36635
rect 3157 36533 3191 36567
rect 9413 36533 9447 36567
rect 10057 36533 10091 36567
rect 10701 36533 10735 36567
rect 11897 36533 11931 36567
rect 12909 36533 12943 36567
rect 19441 36533 19475 36567
rect 24317 36533 24351 36567
rect 31585 36533 31619 36567
rect 32321 36533 32355 36567
rect 32965 36533 32999 36567
rect 35909 36533 35943 36567
rect 36829 36533 36863 36567
rect 8493 36329 8527 36363
rect 26617 36329 26651 36363
rect 37381 36329 37415 36363
rect 7849 36261 7883 36295
rect 29745 36261 29779 36295
rect 36093 36261 36127 36295
rect 1593 36193 1627 36227
rect 12909 36193 12943 36227
rect 14749 36193 14783 36227
rect 15945 36193 15979 36227
rect 20729 36193 20763 36227
rect 23765 36193 23799 36227
rect 24869 36193 24903 36227
rect 25145 36193 25179 36227
rect 27813 36193 27847 36227
rect 4169 36125 4203 36159
rect 6745 36125 6779 36159
rect 7757 36125 7791 36159
rect 8401 36125 8435 36159
rect 9597 36125 9631 36159
rect 10333 36125 10367 36159
rect 10977 36125 11011 36159
rect 11621 36125 11655 36159
rect 13093 36125 13127 36159
rect 27077 36125 27111 36159
rect 27721 36125 27755 36159
rect 28357 36135 28391 36169
rect 29193 36125 29227 36159
rect 29929 36125 29963 36159
rect 30941 36125 30975 36159
rect 34897 36125 34931 36159
rect 35909 36125 35943 36159
rect 36645 36125 36679 36159
rect 36921 36125 36955 36159
rect 37565 36125 37599 36159
rect 38025 36125 38059 36159
rect 1777 36057 1811 36091
rect 3433 36057 3467 36091
rect 14473 36057 14507 36091
rect 14565 36057 14599 36091
rect 16221 36057 16255 36091
rect 17969 36057 18003 36091
rect 21005 36057 21039 36091
rect 22937 36057 22971 36091
rect 27169 36057 27203 36091
rect 31217 36057 31251 36091
rect 3985 35989 4019 36023
rect 6837 35989 6871 36023
rect 9689 35989 9723 36023
rect 10425 35989 10459 36023
rect 11069 35989 11103 36023
rect 11713 35989 11747 36023
rect 13553 35989 13587 36023
rect 22477 35989 22511 36023
rect 28457 35989 28491 36023
rect 29009 35989 29043 36023
rect 32689 35989 32723 36023
rect 34989 35989 35023 36023
rect 38209 35989 38243 36023
rect 2421 35785 2455 35819
rect 14473 35785 14507 35819
rect 30205 35785 30239 35819
rect 3065 35717 3099 35751
rect 3157 35717 3191 35751
rect 6653 35717 6687 35751
rect 11906 35717 11940 35751
rect 15393 35717 15427 35751
rect 16313 35717 16347 35751
rect 33517 35717 33551 35751
rect 1593 35649 1627 35683
rect 2329 35649 2363 35683
rect 6561 35649 6595 35683
rect 8309 35649 8343 35683
rect 10609 35649 10643 35683
rect 16865 35649 16899 35683
rect 22293 35649 22327 35683
rect 30389 35649 30423 35683
rect 36277 35649 36311 35683
rect 38025 35649 38059 35683
rect 3709 35581 3743 35615
rect 9505 35581 9539 35615
rect 9689 35581 9723 35615
rect 11805 35581 11839 35615
rect 12817 35581 12851 35615
rect 13277 35581 13311 35615
rect 15301 35581 15335 35615
rect 17141 35581 17175 35615
rect 19349 35581 19383 35615
rect 19625 35581 19659 35615
rect 21097 35581 21131 35615
rect 22569 35581 22603 35615
rect 27169 35581 27203 35615
rect 27353 35581 27387 35615
rect 27629 35581 27663 35615
rect 33241 35581 33275 35615
rect 35633 35581 35667 35615
rect 1777 35513 1811 35547
rect 10701 35513 10735 35547
rect 8401 35445 8435 35479
rect 10149 35445 10183 35479
rect 18613 35445 18647 35479
rect 24041 35445 24075 35479
rect 34989 35445 35023 35479
rect 36369 35445 36403 35479
rect 38209 35445 38243 35479
rect 1593 35241 1627 35275
rect 38209 35241 38243 35275
rect 2237 35173 2271 35207
rect 37381 35173 37415 35207
rect 10609 35105 10643 35139
rect 11069 35105 11103 35139
rect 13093 35105 13127 35139
rect 15393 35105 15427 35139
rect 18705 35105 18739 35139
rect 20453 35105 20487 35139
rect 23029 35105 23063 35139
rect 30205 35105 30239 35139
rect 32321 35105 32355 35139
rect 1777 35037 1811 35071
rect 2421 35037 2455 35071
rect 4353 35037 4387 35071
rect 6469 35037 6503 35071
rect 8401 35037 8435 35071
rect 10425 35037 10459 35071
rect 14289 35037 14323 35071
rect 17233 35037 17267 35071
rect 22937 35037 22971 35071
rect 34897 35037 34931 35071
rect 37565 35037 37599 35071
rect 38025 35037 38059 35071
rect 9321 34969 9355 35003
rect 9413 34969 9447 35003
rect 9965 34969 9999 35003
rect 13185 34969 13219 35003
rect 13737 34969 13771 35003
rect 15577 34969 15611 35003
rect 17969 34969 18003 35003
rect 20729 34969 20763 35003
rect 30297 34969 30331 35003
rect 31217 34969 31251 35003
rect 32597 34969 32631 35003
rect 34345 34969 34379 35003
rect 35173 34969 35207 35003
rect 36921 34969 36955 35003
rect 4445 34901 4479 34935
rect 6561 34901 6595 34935
rect 8493 34901 8527 34935
rect 14381 34901 14415 34935
rect 22201 34901 22235 34935
rect 2421 34697 2455 34731
rect 4813 34697 4847 34731
rect 10977 34697 11011 34731
rect 20269 34697 20303 34731
rect 24317 34697 24351 34731
rect 31493 34697 31527 34731
rect 34069 34697 34103 34731
rect 3985 34629 4019 34663
rect 9505 34629 9539 34663
rect 11805 34629 11839 34663
rect 13185 34629 13219 34663
rect 13737 34629 13771 34663
rect 14828 34629 14862 34663
rect 18797 34629 18831 34663
rect 20913 34629 20947 34663
rect 30757 34629 30791 34663
rect 35725 34629 35759 34663
rect 35817 34629 35851 34663
rect 1593 34561 1627 34595
rect 2329 34561 2363 34595
rect 3893 34561 3927 34595
rect 4997 34561 5031 34595
rect 8217 34561 8251 34595
rect 8309 34561 8343 34595
rect 10885 34561 10919 34595
rect 11713 34561 11747 34595
rect 14565 34561 14599 34595
rect 18521 34561 18555 34595
rect 20821 34561 20855 34595
rect 22569 34561 22603 34595
rect 27169 34561 27203 34595
rect 30021 34561 30055 34595
rect 31401 34561 31435 34595
rect 32321 34561 32355 34595
rect 38025 34561 38059 34595
rect 9413 34493 9447 34527
rect 10425 34493 10459 34527
rect 13093 34493 13127 34527
rect 22845 34493 22879 34527
rect 29193 34493 29227 34527
rect 36185 34493 36219 34527
rect 1777 34357 1811 34391
rect 16313 34357 16347 34391
rect 27432 34357 27466 34391
rect 32584 34357 32618 34391
rect 38209 34357 38243 34391
rect 13277 34153 13311 34187
rect 14381 34153 14415 34187
rect 25513 34153 25547 34187
rect 30021 34153 30055 34187
rect 34161 34153 34195 34187
rect 15393 34017 15427 34051
rect 19625 34017 19659 34051
rect 19901 34017 19935 34051
rect 31401 34017 31435 34051
rect 34897 34017 34931 34051
rect 36645 34017 36679 34051
rect 2145 33949 2179 33983
rect 2789 33949 2823 33983
rect 9137 33949 9171 33983
rect 11345 33949 11379 33983
rect 11989 33949 12023 33983
rect 13185 33949 13219 33983
rect 14565 33949 14599 33983
rect 22201 33949 22235 33983
rect 25421 33949 25455 33983
rect 29929 33949 29963 33983
rect 34069 33949 34103 33983
rect 11437 33881 11471 33915
rect 15669 33881 15703 33915
rect 22477 33881 22511 33915
rect 27445 33881 27479 33915
rect 27537 33881 27571 33915
rect 28457 33881 28491 33915
rect 31677 33881 31711 33915
rect 35173 33881 35207 33915
rect 1961 33813 1995 33847
rect 2881 33813 2915 33847
rect 9229 33813 9263 33847
rect 12081 33813 12115 33847
rect 17141 33813 17175 33847
rect 21373 33813 21407 33847
rect 23949 33813 23983 33847
rect 33149 33813 33183 33847
rect 11805 33609 11839 33643
rect 18613 33609 18647 33643
rect 21005 33609 21039 33643
rect 24961 33609 24995 33643
rect 35265 33609 35299 33643
rect 4537 33541 4571 33575
rect 8033 33541 8067 33575
rect 8125 33541 8159 33575
rect 10425 33541 10459 33575
rect 19533 33541 19567 33575
rect 25697 33541 25731 33575
rect 33793 33541 33827 33575
rect 36001 33541 36035 33575
rect 8677 33473 8711 33507
rect 9137 33473 9171 33507
rect 11713 33473 11747 33507
rect 12357 33473 12391 33507
rect 13461 33473 13495 33507
rect 14197 33473 14231 33507
rect 16865 33473 16899 33507
rect 19257 33473 19291 33507
rect 28457 33473 28491 33507
rect 30941 33473 30975 33507
rect 32965 33473 32999 33507
rect 35173 33473 35207 33507
rect 4445 33405 4479 33439
rect 5365 33405 5399 33439
rect 10333 33405 10367 33439
rect 10609 33405 10643 33439
rect 12449 33405 12483 33439
rect 17141 33405 17175 33439
rect 23213 33405 23247 33439
rect 23489 33405 23523 33439
rect 25605 33405 25639 33439
rect 26249 33405 26283 33439
rect 28733 33405 28767 33439
rect 30481 33405 30515 33439
rect 35909 33405 35943 33439
rect 36185 33405 36219 33439
rect 9229 33269 9263 33303
rect 13277 33269 13311 33303
rect 14289 33269 14323 33303
rect 31033 33269 31067 33303
rect 9229 33065 9263 33099
rect 10333 33065 10367 33099
rect 22569 32997 22603 33031
rect 25053 32997 25087 33031
rect 13737 32929 13771 32963
rect 20821 32929 20855 32963
rect 25973 32929 26007 32963
rect 27537 32929 27571 32963
rect 28457 32929 28491 32963
rect 1593 32861 1627 32895
rect 7389 32861 7423 32895
rect 9137 32861 9171 32895
rect 10241 32861 10275 32895
rect 10885 32861 10919 32895
rect 11529 32861 11563 32895
rect 11621 32861 11655 32895
rect 14841 32861 14875 32895
rect 24961 32861 24995 32895
rect 27353 32861 27387 32895
rect 37473 32861 37507 32895
rect 37749 32861 37783 32895
rect 10977 32793 11011 32827
rect 12725 32793 12759 32827
rect 12817 32793 12851 32827
rect 21097 32793 21131 32827
rect 1777 32725 1811 32759
rect 7481 32725 7515 32759
rect 14933 32725 14967 32759
rect 10333 32521 10367 32555
rect 11805 32521 11839 32555
rect 38117 32521 38151 32555
rect 7297 32453 7331 32487
rect 7849 32453 7883 32487
rect 17141 32453 17175 32487
rect 19993 32453 20027 32487
rect 1593 32385 1627 32419
rect 10241 32385 10275 32419
rect 11713 32385 11747 32419
rect 12357 32385 12391 32419
rect 13645 32385 13679 32419
rect 16865 32385 16899 32419
rect 23121 32385 23155 32419
rect 38301 32385 38335 32419
rect 7205 32317 7239 32351
rect 19717 32317 19751 32351
rect 23857 32317 23891 32351
rect 24777 32317 24811 32351
rect 25053 32317 25087 32351
rect 12449 32249 12483 32283
rect 1777 32181 1811 32215
rect 13737 32181 13771 32215
rect 18613 32181 18647 32215
rect 21465 32181 21499 32215
rect 26525 32181 26559 32215
rect 9229 31977 9263 32011
rect 24685 31977 24719 32011
rect 26985 31977 27019 32011
rect 36185 31977 36219 32011
rect 16865 31909 16899 31943
rect 24041 31909 24075 31943
rect 11161 31841 11195 31875
rect 12173 31841 12207 31875
rect 12725 31841 12759 31875
rect 13369 31841 13403 31875
rect 15393 31841 15427 31875
rect 19441 31841 19475 31875
rect 19717 31841 19751 31875
rect 21189 31841 21223 31875
rect 22569 31841 22603 31875
rect 32321 31841 32355 31875
rect 9137 31773 9171 31807
rect 9781 31773 9815 31807
rect 9873 31773 9907 31807
rect 15117 31773 15151 31807
rect 22293 31773 22327 31807
rect 24593 31773 24627 31807
rect 26893 31773 26927 31807
rect 27537 31773 27571 31807
rect 27629 31773 27663 31807
rect 32045 31773 32079 31807
rect 34069 31773 34103 31807
rect 36093 31773 36127 31807
rect 11253 31705 11287 31739
rect 12817 31705 12851 31739
rect 4261 31433 4295 31467
rect 6653 31433 6687 31467
rect 11805 31433 11839 31467
rect 8125 31365 8159 31399
rect 8217 31365 8251 31399
rect 9965 31365 9999 31399
rect 13369 31365 13403 31399
rect 4169 31297 4203 31331
rect 6561 31297 6595 31331
rect 9229 31297 9263 31331
rect 9873 31297 9907 31331
rect 10517 31297 10551 31331
rect 11713 31297 11747 31331
rect 15025 31297 15059 31331
rect 18613 31297 18647 31331
rect 35725 31297 35759 31331
rect 13277 31229 13311 31263
rect 14105 31229 14139 31263
rect 15117 31229 15151 31263
rect 18889 31229 18923 31263
rect 33517 31229 33551 31263
rect 33793 31229 33827 31263
rect 8677 31161 8711 31195
rect 9321 31093 9355 31127
rect 10609 31093 10643 31127
rect 20361 31093 20395 31127
rect 35265 31093 35299 31127
rect 35817 31093 35851 31127
rect 24856 30889 24890 30923
rect 31020 30889 31054 30923
rect 14289 30821 14323 30855
rect 9505 30753 9539 30787
rect 10701 30753 10735 30787
rect 11713 30753 11747 30787
rect 13461 30753 13495 30787
rect 15209 30753 15243 30787
rect 17233 30753 17267 30787
rect 18705 30753 18739 30787
rect 19625 30753 19659 30787
rect 21833 30753 21867 30787
rect 23857 30753 23891 30787
rect 24593 30753 24627 30787
rect 30757 30753 30791 30787
rect 34161 30753 34195 30787
rect 36277 30753 36311 30787
rect 36461 30753 36495 30787
rect 37289 30753 37323 30787
rect 1593 30685 1627 30719
rect 12173 30685 12207 30719
rect 14473 30685 14507 30719
rect 17969 30685 18003 30719
rect 33425 30685 33459 30719
rect 9597 30617 9631 30651
rect 10149 30617 10183 30651
rect 10793 30617 10827 30651
rect 13093 30617 13127 30651
rect 13185 30617 13219 30651
rect 15485 30617 15519 30651
rect 19901 30617 19935 30651
rect 22109 30617 22143 30651
rect 26617 30617 26651 30651
rect 32781 30617 32815 30651
rect 1777 30549 1811 30583
rect 12265 30549 12299 30583
rect 21373 30549 21407 30583
rect 9229 30345 9263 30379
rect 10506 30277 10540 30311
rect 10609 30277 10643 30311
rect 11897 30277 11931 30311
rect 13461 30277 13495 30311
rect 9137 30209 9171 30243
rect 9781 30209 9815 30243
rect 13369 30209 13403 30243
rect 14565 30209 14599 30243
rect 18705 30209 18739 30243
rect 29101 30209 29135 30243
rect 38301 30209 38335 30243
rect 9873 30141 9907 30175
rect 11805 30141 11839 30175
rect 12449 30141 12483 30175
rect 14841 30141 14875 30175
rect 18981 30141 19015 30175
rect 29837 30141 29871 30175
rect 34989 30141 35023 30175
rect 35265 30141 35299 30175
rect 11069 30073 11103 30107
rect 16313 30005 16347 30039
rect 20453 30005 20487 30039
rect 36737 30005 36771 30039
rect 38117 30005 38151 30039
rect 11529 29801 11563 29835
rect 14841 29801 14875 29835
rect 33977 29801 34011 29835
rect 10885 29733 10919 29767
rect 12265 29665 12299 29699
rect 15669 29665 15703 29699
rect 29745 29665 29779 29699
rect 31769 29665 31803 29699
rect 32229 29665 32263 29699
rect 34897 29665 34931 29699
rect 1593 29597 1627 29631
rect 10793 29597 10827 29631
rect 11437 29597 11471 29631
rect 14749 29597 14783 29631
rect 15393 29597 15427 29631
rect 17417 29597 17451 29631
rect 20637 29597 20671 29631
rect 27445 29597 27479 29631
rect 4077 29529 4111 29563
rect 12357 29529 12391 29563
rect 13277 29529 13311 29563
rect 20913 29529 20947 29563
rect 22661 29529 22695 29563
rect 25697 29529 25731 29563
rect 30021 29529 30055 29563
rect 32505 29529 32539 29563
rect 35173 29529 35207 29563
rect 36921 29529 36955 29563
rect 38117 29529 38151 29563
rect 1777 29461 1811 29495
rect 4169 29461 4203 29495
rect 38209 29461 38243 29495
rect 4721 29257 4755 29291
rect 11805 29257 11839 29291
rect 9689 29189 9723 29223
rect 9781 29189 9815 29223
rect 13185 29189 13219 29223
rect 14105 29189 14139 29223
rect 20545 29189 20579 29223
rect 4905 29121 4939 29155
rect 11713 29121 11747 29155
rect 14565 29121 14599 29155
rect 16865 29121 16899 29155
rect 22017 29121 22051 29155
rect 27261 29121 27295 29155
rect 32781 29121 32815 29155
rect 38301 29121 38335 29155
rect 1593 29053 1627 29087
rect 1869 29053 1903 29087
rect 10701 29053 10735 29087
rect 13093 29053 13127 29087
rect 17693 29053 17727 29087
rect 18337 29053 18371 29087
rect 21281 29053 21315 29087
rect 34529 29053 34563 29087
rect 14657 28985 14691 29019
rect 22109 28985 22143 29019
rect 29009 28985 29043 29019
rect 38117 28985 38151 29019
rect 18594 28917 18628 28951
rect 20085 28917 20119 28951
rect 27518 28917 27552 28951
rect 33044 28917 33078 28951
rect 6929 28713 6963 28747
rect 11253 28713 11287 28747
rect 8493 28645 8527 28679
rect 7665 28577 7699 28611
rect 10057 28577 10091 28611
rect 12081 28577 12115 28611
rect 12449 28577 12483 28611
rect 16221 28577 16255 28611
rect 32505 28577 32539 28611
rect 4537 28509 4571 28543
rect 5181 28509 5215 28543
rect 6837 28509 6871 28543
rect 7573 28509 7607 28543
rect 11161 28509 11195 28543
rect 13553 28509 13587 28543
rect 20361 28509 20395 28543
rect 8309 28441 8343 28475
rect 10149 28441 10183 28475
rect 10701 28441 10735 28475
rect 12173 28441 12207 28475
rect 16497 28441 16531 28475
rect 20637 28441 20671 28475
rect 32781 28441 32815 28475
rect 4353 28373 4387 28407
rect 4997 28373 5031 28407
rect 13645 28373 13679 28407
rect 17969 28373 18003 28407
rect 22109 28373 22143 28407
rect 34253 28373 34287 28407
rect 13001 28101 13035 28135
rect 27445 28101 27479 28135
rect 29193 28101 29227 28135
rect 33425 28101 33459 28135
rect 7757 28033 7791 28067
rect 9137 28033 9171 28067
rect 10241 28033 10275 28067
rect 11713 28033 11747 28067
rect 14565 28033 14599 28067
rect 22017 28033 22051 28067
rect 9321 27965 9355 27999
rect 12909 27965 12943 27999
rect 13369 27965 13403 27999
rect 14841 27965 14875 27999
rect 17785 27965 17819 27999
rect 18061 27965 18095 27999
rect 19809 27965 19843 27999
rect 24041 27965 24075 27999
rect 27169 27965 27203 27999
rect 33149 27965 33183 27999
rect 7849 27829 7883 27863
rect 9505 27829 9539 27863
rect 10333 27829 10367 27863
rect 11805 27829 11839 27863
rect 16313 27829 16347 27863
rect 22280 27829 22314 27863
rect 34897 27829 34931 27863
rect 15932 27625 15966 27659
rect 32854 27625 32888 27659
rect 35160 27625 35194 27659
rect 7297 27557 7331 27591
rect 8309 27557 8343 27591
rect 14381 27557 14415 27591
rect 8125 27489 8159 27523
rect 13001 27489 13035 27523
rect 13277 27489 13311 27523
rect 15669 27489 15703 27523
rect 19441 27489 19475 27523
rect 21189 27489 21223 27523
rect 28457 27489 28491 27523
rect 30113 27489 30147 27523
rect 32597 27489 32631 27523
rect 6837 27421 6871 27455
rect 7481 27421 7515 27455
rect 7941 27421 7975 27455
rect 12081 27421 12115 27455
rect 14289 27421 14323 27455
rect 26709 27421 26743 27455
rect 34897 27421 34931 27455
rect 38301 27421 38335 27455
rect 1685 27353 1719 27387
rect 1869 27353 1903 27387
rect 11437 27353 11471 27387
rect 11529 27353 11563 27387
rect 13093 27353 13127 27387
rect 19717 27353 19751 27387
rect 26985 27353 27019 27387
rect 30389 27353 30423 27387
rect 32137 27353 32171 27387
rect 6653 27285 6687 27319
rect 17417 27285 17451 27319
rect 21557 27285 21591 27319
rect 34345 27285 34379 27319
rect 36645 27285 36679 27319
rect 38117 27285 38151 27319
rect 12081 27081 12115 27115
rect 16957 27081 16991 27115
rect 21373 27081 21407 27115
rect 8493 27013 8527 27047
rect 8585 27013 8619 27047
rect 33793 27013 33827 27047
rect 7021 26945 7055 26979
rect 11989 26945 12023 26979
rect 14565 26945 14599 26979
rect 16865 26945 16899 26979
rect 18153 26945 18187 26979
rect 21281 26945 21315 26979
rect 27629 26945 27663 26979
rect 6837 26877 6871 26911
rect 9505 26877 9539 26911
rect 14841 26877 14875 26911
rect 18429 26877 18463 26911
rect 28365 26877 28399 26911
rect 29561 26877 29595 26911
rect 29837 26877 29871 26911
rect 33517 26877 33551 26911
rect 35541 26877 35575 26911
rect 7205 26809 7239 26843
rect 16313 26741 16347 26775
rect 19901 26741 19935 26775
rect 31309 26741 31343 26775
rect 1593 26537 1627 26571
rect 27813 26537 27847 26571
rect 7849 26469 7883 26503
rect 33241 26469 33275 26503
rect 38117 26469 38151 26503
rect 9229 26401 9263 26435
rect 13369 26401 13403 26435
rect 15669 26401 15703 26435
rect 15945 26401 15979 26435
rect 20729 26401 20763 26435
rect 22753 26401 22787 26435
rect 26065 26401 26099 26435
rect 31493 26401 31527 26435
rect 35633 26401 35667 26435
rect 1777 26333 1811 26367
rect 7757 26333 7791 26367
rect 9137 26333 9171 26367
rect 10885 26333 10919 26367
rect 38301 26333 38335 26367
rect 10977 26265 11011 26299
rect 12725 26265 12759 26299
rect 12817 26265 12851 26299
rect 21005 26265 21039 26299
rect 26341 26265 26375 26299
rect 31769 26265 31803 26299
rect 34897 26265 34931 26299
rect 5457 26197 5491 26231
rect 17417 26197 17451 26231
rect 11805 25993 11839 26027
rect 13829 25993 13863 26027
rect 37749 25993 37783 26027
rect 9505 25925 9539 25959
rect 10241 25925 10275 25959
rect 29653 25925 29687 25959
rect 33977 25925 34011 25959
rect 5365 25857 5399 25891
rect 7481 25857 7515 25891
rect 9413 25857 9447 25891
rect 11713 25857 11747 25891
rect 13737 25857 13771 25891
rect 27169 25857 27203 25891
rect 29377 25857 29411 25891
rect 33701 25857 33735 25891
rect 37933 25857 37967 25891
rect 5549 25789 5583 25823
rect 8769 25789 8803 25823
rect 10149 25789 10183 25823
rect 10793 25789 10827 25823
rect 19625 25789 19659 25823
rect 19901 25789 19935 25823
rect 22937 25789 22971 25823
rect 23213 25789 23247 25823
rect 24685 25789 24719 25823
rect 27445 25789 27479 25823
rect 35725 25789 35759 25823
rect 6009 25653 6043 25687
rect 7573 25653 7607 25687
rect 21373 25653 21407 25687
rect 28917 25653 28951 25687
rect 31125 25653 31159 25687
rect 7941 25449 7975 25483
rect 17049 25449 17083 25483
rect 22372 25449 22406 25483
rect 26893 25449 26927 25483
rect 32321 25449 32355 25483
rect 37197 25449 37231 25483
rect 4905 25313 4939 25347
rect 7297 25313 7331 25347
rect 9229 25313 9263 25347
rect 25145 25313 25179 25347
rect 30573 25313 30607 25347
rect 35173 25313 35207 25347
rect 5089 25245 5123 25279
rect 7481 25245 7515 25279
rect 10425 25245 10459 25279
rect 14657 25245 14691 25279
rect 15301 25245 15335 25279
rect 17693 25245 17727 25279
rect 22098 25245 22132 25279
rect 34897 25245 34931 25279
rect 37105 25245 37139 25279
rect 38025 25245 38059 25279
rect 9321 25177 9355 25211
rect 9873 25177 9907 25211
rect 15577 25177 15611 25211
rect 18429 25177 18463 25211
rect 25421 25177 25455 25211
rect 30849 25177 30883 25211
rect 5549 25109 5583 25143
rect 10517 25109 10551 25143
rect 14749 25109 14783 25143
rect 23857 25109 23891 25143
rect 36645 25109 36679 25143
rect 38209 25109 38243 25143
rect 5273 24905 5307 24939
rect 10241 24837 10275 24871
rect 12173 24837 12207 24871
rect 22845 24837 22879 24871
rect 1593 24769 1627 24803
rect 4077 24769 4111 24803
rect 4721 24769 4755 24803
rect 5181 24769 5215 24803
rect 5825 24769 5859 24803
rect 6837 24769 6871 24803
rect 7021 24769 7055 24803
rect 7941 24769 7975 24803
rect 9413 24769 9447 24803
rect 9505 24769 9539 24803
rect 13185 24769 13219 24803
rect 18153 24769 18187 24803
rect 22017 24769 22051 24803
rect 10149 24701 10183 24735
rect 11161 24701 11195 24735
rect 12081 24701 12115 24735
rect 13277 24701 13311 24735
rect 18429 24701 18463 24735
rect 28273 24701 28307 24735
rect 28549 24701 28583 24735
rect 33333 24701 33367 24735
rect 33609 24701 33643 24735
rect 35357 24701 35391 24735
rect 3893 24633 3927 24667
rect 4537 24633 4571 24667
rect 7205 24633 7239 24667
rect 12633 24633 12667 24667
rect 1777 24565 1811 24599
rect 5917 24565 5951 24599
rect 8033 24565 8067 24599
rect 19901 24565 19935 24599
rect 30021 24565 30055 24599
rect 16024 24361 16058 24395
rect 21189 24361 21223 24395
rect 1869 24225 1903 24259
rect 6837 24225 6871 24259
rect 12449 24225 12483 24259
rect 19441 24225 19475 24259
rect 34161 24225 34195 24259
rect 34897 24225 34931 24259
rect 35173 24225 35207 24259
rect 1593 24157 1627 24191
rect 7297 24157 7331 24191
rect 9781 24157 9815 24191
rect 13277 24157 13311 24191
rect 15761 24157 15795 24191
rect 28273 24157 28307 24191
rect 29745 24157 29779 24191
rect 33425 24157 33459 24191
rect 38301 24157 38335 24191
rect 6193 24089 6227 24123
rect 6285 24089 6319 24123
rect 7389 24089 7423 24123
rect 12173 24089 12207 24123
rect 12265 24089 12299 24123
rect 17785 24089 17819 24123
rect 19717 24089 19751 24123
rect 29009 24089 29043 24123
rect 30021 24089 30055 24123
rect 9873 24021 9907 24055
rect 13369 24021 13403 24055
rect 31493 24021 31527 24055
rect 36645 24021 36679 24055
rect 38117 24021 38151 24055
rect 10517 23817 10551 23851
rect 12909 23817 12943 23851
rect 18613 23817 18647 23851
rect 34069 23817 34103 23851
rect 8309 23749 8343 23783
rect 9965 23749 9999 23783
rect 21465 23749 21499 23783
rect 23949 23749 23983 23783
rect 5549 23681 5583 23715
rect 6745 23681 6779 23715
rect 10425 23681 10459 23715
rect 12817 23681 12851 23715
rect 14565 23681 14599 23715
rect 16865 23681 16899 23715
rect 23673 23681 23707 23715
rect 34529 23681 34563 23715
rect 8125 23613 8159 23647
rect 14841 23613 14875 23647
rect 19441 23613 19475 23647
rect 19717 23613 19751 23647
rect 25697 23613 25731 23647
rect 28641 23613 28675 23647
rect 28917 23613 28951 23647
rect 32321 23613 32355 23647
rect 32597 23613 32631 23647
rect 34805 23613 34839 23647
rect 6561 23545 6595 23579
rect 16313 23545 16347 23579
rect 5641 23477 5675 23511
rect 17128 23477 17162 23511
rect 30389 23477 30423 23511
rect 36277 23477 36311 23511
rect 16773 23273 16807 23307
rect 37841 23273 37875 23307
rect 33701 23205 33735 23239
rect 9689 23137 9723 23171
rect 10333 23137 10367 23171
rect 15025 23137 15059 23171
rect 19809 23137 19843 23171
rect 21833 23137 21867 23171
rect 22293 23137 22327 23171
rect 24041 23137 24075 23171
rect 26065 23137 26099 23171
rect 29745 23137 29779 23171
rect 31493 23137 31527 23171
rect 32229 23137 32263 23171
rect 34897 23137 34931 23171
rect 35173 23137 35207 23171
rect 36921 23137 36955 23171
rect 8401 23069 8435 23103
rect 11345 23069 11379 23103
rect 12449 23069 12483 23103
rect 13093 23069 13127 23103
rect 25789 23069 25823 23103
rect 31953 23069 31987 23103
rect 38025 23069 38059 23103
rect 9781 23001 9815 23035
rect 13185 23001 13219 23035
rect 15301 23001 15335 23035
rect 20085 23001 20119 23035
rect 22569 23001 22603 23035
rect 27813 23001 27847 23035
rect 30021 23001 30055 23035
rect 8493 22933 8527 22967
rect 11437 22933 11471 22967
rect 12541 22933 12575 22967
rect 1593 22729 1627 22763
rect 13001 22729 13035 22763
rect 22109 22729 22143 22763
rect 36737 22729 36771 22763
rect 9413 22661 9447 22695
rect 11897 22661 11931 22695
rect 19717 22661 19751 22695
rect 27445 22661 27479 22695
rect 1777 22593 1811 22627
rect 10793 22593 10827 22627
rect 12909 22593 12943 22627
rect 17693 22593 17727 22627
rect 22017 22593 22051 22627
rect 22661 22593 22695 22627
rect 24685 22593 24719 22627
rect 27169 22593 27203 22627
rect 32781 22593 32815 22627
rect 34989 22593 35023 22627
rect 38025 22593 38059 22627
rect 4537 22525 4571 22559
rect 9321 22525 9355 22559
rect 10333 22525 10367 22559
rect 11805 22525 11839 22559
rect 12081 22525 12115 22559
rect 17969 22525 18003 22559
rect 22937 22525 22971 22559
rect 28917 22525 28951 22559
rect 33057 22525 33091 22559
rect 35265 22525 35299 22559
rect 38209 22457 38243 22491
rect 10885 22389 10919 22423
rect 34529 22389 34563 22423
rect 18705 22185 18739 22219
rect 25770 22185 25804 22219
rect 36829 22185 36863 22219
rect 4445 22049 4479 22083
rect 9873 22049 9907 22083
rect 12817 22049 12851 22083
rect 16221 22049 16255 22083
rect 20729 22049 20763 22083
rect 22201 22049 22235 22083
rect 23029 22049 23063 22083
rect 25513 22049 25547 22083
rect 31033 22049 31067 22083
rect 37473 22049 37507 22083
rect 4629 21981 4663 22015
rect 8401 21981 8435 22015
rect 16129 21981 16163 22015
rect 18637 21981 18671 22015
rect 20637 21981 20671 22015
rect 22753 21981 22787 22015
rect 36737 21981 36771 22015
rect 37381 21981 37415 22015
rect 38025 21981 38059 22015
rect 9229 21913 9263 21947
rect 9321 21913 9355 21947
rect 12357 21913 12391 21947
rect 12449 21913 12483 21947
rect 14657 21913 14691 21947
rect 14749 21913 14783 21947
rect 15669 21913 15703 21947
rect 21373 21913 21407 21947
rect 31309 21913 31343 21947
rect 34989 21913 35023 21947
rect 35081 21913 35115 21947
rect 36001 21913 36035 21947
rect 5089 21845 5123 21879
rect 8493 21845 8527 21879
rect 27261 21845 27295 21879
rect 32781 21845 32815 21879
rect 38209 21845 38243 21879
rect 4813 21641 4847 21675
rect 5457 21641 5491 21675
rect 25053 21641 25087 21675
rect 30481 21641 30515 21675
rect 31677 21641 31711 21675
rect 35725 21641 35759 21675
rect 36645 21641 36679 21675
rect 37565 21641 37599 21675
rect 9229 21573 9263 21607
rect 13185 21573 13219 21607
rect 17785 21573 17819 21607
rect 21281 21573 21315 21607
rect 33333 21573 33367 21607
rect 38209 21573 38243 21607
rect 1685 21505 1719 21539
rect 2513 21505 2547 21539
rect 4997 21505 5031 21539
rect 5641 21505 5675 21539
rect 7665 21505 7699 21539
rect 10609 21505 10643 21539
rect 12357 21505 12391 21539
rect 13093 21505 13127 21539
rect 16865 21505 16899 21539
rect 17693 21505 17727 21539
rect 21005 21505 21039 21539
rect 22017 21505 22051 21539
rect 24961 21505 24995 21539
rect 25605 21505 25639 21539
rect 30389 21505 30423 21539
rect 31585 21505 31619 21539
rect 34713 21505 34747 21539
rect 35633 21505 35667 21539
rect 36553 21505 36587 21539
rect 37473 21505 37507 21539
rect 38117 21505 38151 21539
rect 8401 21437 8435 21471
rect 9137 21437 9171 21471
rect 10149 21437 10183 21471
rect 22845 21437 22879 21471
rect 33241 21437 33275 21471
rect 33517 21437 33551 21471
rect 1869 21369 1903 21403
rect 7757 21369 7791 21403
rect 2329 21301 2363 21335
rect 10701 21301 10735 21335
rect 12449 21301 12483 21335
rect 16957 21301 16991 21335
rect 25697 21301 25731 21335
rect 34713 21301 34747 21335
rect 1777 21097 1811 21131
rect 18153 21097 18187 21131
rect 19533 21097 19567 21131
rect 21189 21097 21223 21131
rect 29009 21097 29043 21131
rect 29837 21097 29871 21131
rect 30757 21097 30791 21131
rect 32045 21097 32079 21131
rect 34161 21097 34195 21131
rect 36553 21097 36587 21131
rect 37841 21097 37875 21131
rect 23397 21029 23431 21063
rect 37197 21029 37231 21063
rect 8125 20961 8159 20995
rect 10333 20961 10367 20995
rect 11345 20961 11379 20995
rect 15209 20961 15243 20995
rect 15393 20961 15427 20995
rect 22109 20961 22143 20995
rect 31401 20961 31435 20995
rect 35265 20961 35299 20995
rect 11253 20893 11287 20927
rect 12173 20893 12207 20927
rect 13093 20893 13127 20927
rect 13553 20893 13587 20927
rect 14565 20893 14599 20927
rect 14657 20893 14691 20927
rect 18061 20893 18095 20927
rect 18705 20893 18739 20927
rect 19441 20893 19475 20927
rect 21373 20893 21407 20927
rect 21833 20893 21867 20927
rect 23305 20893 23339 20927
rect 26249 20893 26283 20927
rect 27169 20893 27203 20927
rect 28917 20893 28951 20927
rect 29745 20893 29779 20927
rect 30665 20893 30699 20927
rect 31309 20893 31343 20927
rect 31953 20893 31987 20927
rect 34345 20893 34379 20927
rect 36461 20893 36495 20927
rect 37105 20893 37139 20927
rect 37749 20893 37783 20927
rect 1685 20825 1719 20859
rect 7481 20825 7515 20859
rect 7573 20825 7607 20859
rect 9781 20825 9815 20859
rect 9873 20825 9907 20859
rect 13645 20825 13679 20859
rect 17049 20825 17083 20859
rect 24685 20825 24719 20859
rect 24777 20825 24811 20859
rect 25697 20825 25731 20859
rect 26525 20825 26559 20859
rect 32689 20825 32723 20859
rect 32781 20825 32815 20859
rect 33333 20825 33367 20859
rect 34989 20825 35023 20859
rect 35081 20825 35115 20859
rect 12265 20757 12299 20791
rect 12909 20757 12943 20791
rect 18797 20757 18831 20791
rect 27261 20757 27295 20791
rect 1777 20553 1811 20587
rect 12357 20553 12391 20587
rect 17509 20553 17543 20587
rect 18889 20553 18923 20587
rect 25789 20553 25823 20587
rect 29193 20553 29227 20587
rect 31125 20553 31159 20587
rect 33057 20553 33091 20587
rect 35725 20553 35759 20587
rect 36369 20553 36403 20587
rect 37565 20553 37599 20587
rect 38209 20553 38243 20587
rect 6745 20485 6779 20519
rect 13461 20485 13495 20519
rect 15301 20485 15335 20519
rect 15393 20485 15427 20519
rect 22937 20485 22971 20519
rect 23029 20485 23063 20519
rect 23949 20485 23983 20519
rect 26433 20485 26467 20519
rect 28549 20485 28583 20519
rect 29837 20485 29871 20519
rect 32413 20485 32447 20519
rect 34529 20485 34563 20519
rect 34621 20485 34655 20519
rect 1961 20417 1995 20451
rect 8033 20417 8067 20451
rect 10241 20417 10275 20451
rect 10425 20417 10459 20451
rect 12265 20417 12299 20451
rect 17417 20417 17451 20451
rect 18153 20417 18187 20451
rect 18797 20417 18831 20451
rect 24777 20417 24811 20451
rect 25697 20417 25731 20451
rect 26341 20417 26375 20451
rect 27169 20417 27203 20451
rect 28457 20417 28491 20451
rect 29101 20417 29135 20451
rect 29745 20417 29779 20451
rect 30389 20417 30423 20451
rect 31033 20417 31067 20451
rect 32321 20417 32355 20451
rect 32965 20417 32999 20451
rect 33609 20417 33643 20451
rect 35633 20417 35667 20451
rect 36277 20417 36311 20451
rect 37473 20417 37507 20451
rect 38117 20417 38151 20451
rect 6653 20349 6687 20383
rect 7297 20349 7331 20383
rect 9597 20349 9631 20383
rect 13369 20349 13403 20383
rect 14381 20349 14415 20383
rect 15577 20349 15611 20383
rect 25053 20349 25087 20383
rect 27445 20349 27479 20383
rect 10885 20281 10919 20315
rect 18245 20281 18279 20315
rect 35081 20281 35115 20315
rect 8125 20213 8159 20247
rect 30481 20213 30515 20247
rect 33701 20213 33735 20247
rect 6653 20009 6687 20043
rect 10241 20009 10275 20043
rect 14657 20009 14691 20043
rect 16773 20009 16807 20043
rect 17417 20009 17451 20043
rect 22753 20009 22787 20043
rect 27629 20009 27663 20043
rect 28917 20009 28951 20043
rect 31401 20009 31435 20043
rect 32045 20009 32079 20043
rect 33793 20009 33827 20043
rect 36185 20009 36219 20043
rect 36829 20009 36863 20043
rect 38025 20009 38059 20043
rect 8401 19941 8435 19975
rect 21373 19941 21407 19975
rect 28273 19941 28307 19975
rect 37473 19941 37507 19975
rect 13277 19873 13311 19907
rect 20821 19873 20855 19907
rect 23673 19873 23707 19907
rect 25421 19873 25455 19907
rect 29837 19873 29871 19907
rect 30481 19873 30515 19907
rect 6837 19805 6871 19839
rect 7297 19805 7331 19839
rect 8585 19805 8619 19839
rect 9597 19805 9631 19839
rect 9781 19805 9815 19839
rect 11345 19805 11379 19839
rect 14565 19805 14599 19839
rect 15209 19805 15243 19839
rect 16037 19805 16071 19839
rect 16681 19805 16715 19839
rect 17325 19805 17359 19839
rect 22661 19805 22695 19839
rect 25145 19805 25179 19839
rect 26617 19805 26651 19839
rect 26893 19805 26927 19839
rect 27537 19805 27571 19839
rect 28181 19805 28215 19839
rect 28825 19805 28859 19839
rect 31309 19805 31343 19839
rect 31953 19805 31987 19839
rect 32621 19815 32655 19849
rect 33701 19805 33735 19839
rect 36093 19805 36127 19839
rect 36737 19805 36771 19839
rect 37381 19805 37415 19839
rect 38209 19805 38243 19839
rect 11897 19737 11931 19771
rect 13001 19737 13035 19771
rect 13093 19737 13127 19771
rect 20913 19737 20947 19771
rect 23397 19737 23431 19771
rect 23489 19737 23523 19771
rect 29929 19737 29963 19771
rect 32689 19737 32723 19771
rect 34989 19737 35023 19771
rect 35081 19737 35115 19771
rect 35633 19737 35667 19771
rect 7389 19669 7423 19703
rect 11161 19669 11195 19703
rect 11989 19669 12023 19703
rect 15301 19669 15335 19703
rect 16129 19669 16163 19703
rect 1593 19465 1627 19499
rect 7481 19465 7515 19499
rect 12173 19465 12207 19499
rect 14197 19465 14231 19499
rect 16957 19465 16991 19499
rect 17693 19465 17727 19499
rect 18981 19465 19015 19499
rect 20269 19465 20303 19499
rect 20913 19465 20947 19499
rect 24593 19465 24627 19499
rect 25513 19465 25547 19499
rect 26157 19465 26191 19499
rect 27905 19465 27939 19499
rect 32413 19465 32447 19499
rect 33241 19465 33275 19499
rect 34713 19465 34747 19499
rect 36185 19465 36219 19499
rect 36829 19465 36863 19499
rect 8769 19397 8803 19431
rect 10149 19397 10183 19431
rect 10241 19397 10275 19431
rect 12909 19397 12943 19431
rect 15393 19397 15427 19431
rect 16313 19397 16347 19431
rect 33885 19397 33919 19431
rect 35357 19397 35391 19431
rect 1777 19329 1811 19363
rect 7665 19329 7699 19363
rect 12081 19329 12115 19363
rect 14105 19329 14139 19363
rect 16865 19329 16899 19363
rect 17601 19329 17635 19363
rect 18889 19329 18923 19363
rect 20177 19329 20211 19363
rect 20821 19329 20855 19363
rect 22017 19329 22051 19363
rect 23581 19329 23615 19363
rect 24501 19329 24535 19363
rect 25421 19329 25455 19363
rect 26065 19329 26099 19363
rect 27169 19329 27203 19363
rect 27261 19329 27295 19363
rect 27813 19329 27847 19363
rect 28549 19329 28583 19363
rect 30849 19329 30883 19363
rect 32321 19329 32355 19363
rect 33149 19329 33183 19363
rect 33793 19329 33827 19363
rect 34621 19329 34655 19363
rect 35265 19329 35299 19363
rect 36093 19329 36127 19363
rect 36737 19329 36771 19363
rect 38025 19329 38059 19363
rect 8677 19261 8711 19295
rect 9137 19261 9171 19295
rect 11161 19261 11195 19295
rect 12817 19261 12851 19295
rect 15301 19261 15335 19295
rect 23857 19261 23891 19295
rect 28733 19261 28767 19295
rect 29009 19261 29043 19295
rect 13369 19193 13403 19227
rect 22109 19125 22143 19159
rect 30941 19125 30975 19159
rect 38209 19125 38243 19159
rect 15577 18921 15611 18955
rect 18337 18921 18371 18955
rect 23673 18921 23707 18955
rect 26341 18921 26375 18955
rect 30481 18921 30515 18955
rect 31585 18921 31619 18955
rect 34161 18921 34195 18955
rect 35725 18921 35759 18955
rect 36369 18921 36403 18955
rect 10977 18853 11011 18887
rect 33241 18853 33275 18887
rect 9597 18785 9631 18819
rect 10425 18785 10459 18819
rect 12173 18785 12207 18819
rect 19441 18785 19475 18819
rect 21281 18785 21315 18819
rect 21833 18785 21867 18819
rect 24685 18785 24719 18819
rect 27997 18785 28031 18819
rect 37841 18785 37875 18819
rect 8217 18717 8251 18751
rect 14657 18717 14691 18751
rect 15485 18717 15519 18751
rect 16129 18717 16163 18751
rect 18245 18717 18279 18751
rect 23581 18717 23615 18751
rect 24593 18717 24627 18751
rect 25237 18717 25271 18751
rect 26249 18717 26283 18751
rect 28457 18717 28491 18751
rect 29745 18717 29779 18751
rect 30389 18717 30423 18751
rect 31485 18717 31519 18751
rect 33149 18717 33183 18751
rect 34069 18717 34103 18751
rect 34989 18717 35023 18751
rect 35633 18717 35667 18751
rect 36277 18717 36311 18751
rect 10517 18649 10551 18683
rect 12265 18649 12299 18683
rect 13185 18649 13219 18683
rect 14749 18649 14783 18683
rect 19625 18649 19659 18683
rect 21925 18649 21959 18683
rect 22845 18649 22879 18683
rect 25329 18649 25363 18683
rect 26985 18649 27019 18683
rect 27077 18649 27111 18683
rect 28733 18649 28767 18683
rect 37289 18649 37323 18683
rect 37381 18649 37415 18683
rect 8309 18581 8343 18615
rect 16221 18581 16255 18615
rect 29837 18581 29871 18615
rect 35081 18581 35115 18615
rect 7665 18377 7699 18411
rect 9045 18377 9079 18411
rect 10241 18377 10275 18411
rect 22477 18377 22511 18411
rect 24409 18377 24443 18411
rect 26065 18377 26099 18411
rect 27445 18377 27479 18411
rect 28733 18377 28767 18411
rect 29377 18377 29411 18411
rect 33609 18377 33643 18411
rect 36829 18377 36863 18411
rect 37933 18377 37967 18411
rect 12357 18309 12391 18343
rect 13921 18309 13955 18343
rect 23765 18309 23799 18343
rect 28089 18309 28123 18343
rect 31217 18309 31251 18343
rect 32505 18309 32539 18343
rect 35081 18309 35115 18343
rect 7573 18241 7607 18275
rect 8585 18241 8619 18275
rect 9229 18241 9263 18275
rect 10149 18241 10183 18275
rect 10793 18241 10827 18275
rect 14565 18241 14599 18275
rect 19441 18241 19475 18275
rect 22385 18241 22419 18275
rect 23029 18241 23063 18275
rect 23673 18241 23707 18275
rect 24317 18241 24351 18275
rect 25145 18241 25179 18275
rect 25973 18241 26007 18275
rect 27353 18241 27387 18275
rect 27997 18241 28031 18275
rect 28641 18241 28675 18275
rect 29285 18241 29319 18275
rect 33517 18241 33551 18275
rect 34437 18241 34471 18275
rect 34989 18241 35023 18275
rect 35817 18241 35851 18275
rect 36737 18241 36771 18275
rect 37841 18241 37875 18275
rect 1593 18173 1627 18207
rect 1869 18173 1903 18207
rect 12265 18173 12299 18207
rect 13277 18173 13311 18207
rect 31125 18173 31159 18207
rect 31401 18173 31435 18207
rect 32413 18173 32447 18207
rect 8401 18105 8435 18139
rect 25237 18105 25271 18139
rect 32965 18105 32999 18139
rect 35633 18105 35667 18139
rect 10885 18037 10919 18071
rect 14013 18037 14047 18071
rect 14657 18037 14691 18071
rect 19257 18037 19291 18071
rect 23121 18037 23155 18071
rect 34437 18037 34471 18071
rect 25789 17833 25823 17867
rect 27997 17833 28031 17867
rect 28641 17833 28675 17867
rect 37933 17833 37967 17867
rect 37289 17765 37323 17799
rect 9689 17697 9723 17731
rect 11069 17697 11103 17731
rect 13093 17697 13127 17731
rect 23765 17697 23799 17731
rect 30389 17697 30423 17731
rect 35909 17697 35943 17731
rect 8309 17629 8343 17663
rect 14289 17629 14323 17663
rect 18705 17629 18739 17663
rect 19625 17629 19659 17663
rect 23029 17629 23063 17663
rect 23673 17629 23707 17663
rect 25697 17629 25731 17663
rect 27905 17629 27939 17663
rect 28549 17629 28583 17663
rect 31309 17629 31343 17663
rect 32873 17629 32907 17663
rect 33517 17629 33551 17663
rect 34161 17629 34195 17663
rect 34897 17629 34931 17663
rect 37197 17629 37231 17663
rect 37841 17629 37875 17663
rect 9229 17561 9263 17595
rect 9321 17561 9355 17595
rect 11161 17561 11195 17595
rect 12081 17561 12115 17595
rect 13185 17561 13219 17595
rect 13737 17561 13771 17595
rect 26433 17561 26467 17595
rect 26525 17561 26559 17595
rect 27445 17561 27479 17595
rect 29837 17561 29871 17595
rect 29929 17561 29963 17595
rect 34253 17561 34287 17595
rect 35081 17561 35115 17595
rect 8401 17493 8435 17527
rect 14381 17493 14415 17527
rect 18797 17493 18831 17527
rect 19441 17493 19475 17527
rect 23121 17493 23155 17527
rect 31401 17493 31435 17527
rect 32965 17493 32999 17527
rect 33609 17493 33643 17527
rect 17785 17289 17819 17323
rect 19349 17289 19383 17323
rect 27261 17289 27295 17323
rect 29193 17289 29227 17323
rect 32321 17289 32355 17323
rect 8861 17221 8895 17255
rect 20085 17221 20119 17255
rect 20637 17221 20671 17255
rect 22937 17221 22971 17255
rect 23029 17221 23063 17255
rect 23949 17221 23983 17255
rect 30665 17221 30699 17255
rect 33517 17221 33551 17255
rect 35357 17221 35391 17255
rect 36829 17221 36863 17255
rect 1777 17153 1811 17187
rect 17693 17153 17727 17187
rect 19257 17153 19291 17187
rect 22017 17153 22051 17187
rect 27169 17153 27203 17187
rect 29101 17153 29135 17187
rect 29837 17153 29871 17187
rect 32505 17153 32539 17187
rect 36737 17153 36771 17187
rect 38025 17153 38059 17187
rect 8769 17085 8803 17119
rect 9137 17085 9171 17119
rect 19993 17085 20027 17119
rect 30573 17085 30607 17119
rect 31217 17085 31251 17119
rect 33425 17085 33459 17119
rect 34069 17085 34103 17119
rect 35265 17085 35299 17119
rect 36093 17085 36127 17119
rect 38209 17017 38243 17051
rect 1593 16949 1627 16983
rect 22109 16949 22143 16983
rect 29929 16949 29963 16983
rect 35265 16745 35299 16779
rect 25973 16609 26007 16643
rect 26433 16609 26467 16643
rect 30205 16609 30239 16643
rect 30849 16609 30883 16643
rect 31769 16609 31803 16643
rect 33333 16609 33367 16643
rect 20545 16541 20579 16575
rect 21181 16551 21215 16585
rect 23213 16541 23247 16575
rect 25329 16541 25363 16575
rect 28273 16541 28307 16575
rect 28917 16541 28951 16575
rect 35173 16541 35207 16575
rect 36001 16541 36035 16575
rect 36461 16541 36495 16575
rect 37297 16541 37331 16575
rect 37749 16541 37783 16575
rect 37841 16541 37875 16575
rect 20637 16473 20671 16507
rect 25421 16473 25455 16507
rect 26157 16473 26191 16507
rect 30297 16473 30331 16507
rect 31861 16473 31895 16507
rect 32781 16473 32815 16507
rect 33425 16473 33459 16507
rect 34345 16473 34379 16507
rect 36553 16473 36587 16507
rect 21281 16405 21315 16439
rect 23305 16405 23339 16439
rect 28365 16405 28399 16439
rect 29009 16405 29043 16439
rect 35817 16405 35851 16439
rect 37105 16405 37139 16439
rect 30941 16201 30975 16235
rect 31493 16201 31527 16235
rect 36829 16201 36863 16235
rect 17049 16133 17083 16167
rect 18521 16133 18555 16167
rect 19073 16133 19107 16167
rect 25329 16133 25363 16167
rect 27813 16133 27847 16167
rect 28365 16133 28399 16167
rect 29469 16133 29503 16167
rect 32505 16133 32539 16167
rect 34437 16133 34471 16167
rect 36185 16133 36219 16167
rect 1593 16065 1627 16099
rect 6745 16065 6779 16099
rect 7941 16065 7975 16099
rect 23121 16065 23155 16099
rect 23765 16065 23799 16099
rect 30849 16065 30883 16099
rect 31677 16065 31711 16099
rect 33517 16065 33551 16099
rect 35449 16065 35483 16099
rect 36093 16065 36127 16099
rect 36737 16065 36771 16099
rect 38025 16065 38059 16099
rect 8033 15997 8067 16031
rect 16957 15997 16991 16031
rect 18429 15997 18463 16031
rect 20821 15997 20855 16031
rect 21005 15997 21039 16031
rect 25237 15997 25271 16031
rect 26249 15997 26283 16031
rect 27721 15997 27755 16031
rect 29377 15997 29411 16031
rect 30297 15997 30331 16031
rect 32413 15997 32447 16031
rect 33057 15997 33091 16031
rect 34345 15997 34379 16031
rect 34989 15997 35023 16031
rect 6561 15929 6595 15963
rect 17509 15929 17543 15963
rect 23857 15929 23891 15963
rect 35541 15929 35575 15963
rect 1777 15861 1811 15895
rect 21189 15861 21223 15895
rect 23213 15861 23247 15895
rect 33609 15861 33643 15895
rect 38209 15861 38243 15895
rect 26249 15657 26283 15691
rect 27905 15657 27939 15691
rect 31033 15657 31067 15691
rect 11345 15521 11379 15555
rect 33977 15521 34011 15555
rect 37013 15521 37047 15555
rect 37841 15521 37875 15555
rect 6837 15453 6871 15487
rect 15921 15453 15955 15487
rect 20545 15453 20579 15487
rect 22477 15453 22511 15487
rect 22661 15453 22695 15487
rect 23605 15463 23639 15497
rect 24593 15453 24627 15487
rect 25513 15453 25547 15487
rect 26157 15453 26191 15487
rect 27261 15453 27295 15487
rect 27445 15453 27479 15487
rect 29929 15453 29963 15487
rect 30389 15453 30423 15487
rect 31217 15453 31251 15487
rect 31677 15453 31711 15487
rect 32321 15453 32355 15487
rect 32965 15453 32999 15487
rect 33057 15453 33091 15487
rect 34897 15453 34931 15487
rect 35725 15453 35759 15487
rect 10333 15385 10367 15419
rect 10425 15385 10459 15419
rect 28457 15385 28491 15419
rect 28549 15385 28583 15419
rect 29101 15385 29135 15419
rect 33701 15385 33735 15419
rect 33793 15385 33827 15419
rect 34989 15385 35023 15419
rect 36369 15385 36403 15419
rect 36461 15385 36495 15419
rect 37565 15385 37599 15419
rect 37657 15385 37691 15419
rect 6653 15317 6687 15351
rect 15761 15317 15795 15351
rect 20637 15317 20671 15351
rect 23121 15317 23155 15351
rect 23673 15317 23707 15351
rect 24685 15317 24719 15351
rect 25605 15317 25639 15351
rect 29745 15317 29779 15351
rect 30481 15317 30515 15351
rect 31769 15317 31803 15351
rect 32413 15317 32447 15351
rect 35541 15317 35575 15351
rect 8125 15113 8159 15147
rect 13645 15113 13679 15147
rect 16129 15113 16163 15147
rect 20177 15113 20211 15147
rect 26433 15113 26467 15147
rect 29561 15113 29595 15147
rect 35909 15113 35943 15147
rect 14381 15045 14415 15079
rect 14933 15045 14967 15079
rect 16957 15045 16991 15079
rect 30849 15045 30883 15079
rect 38301 15045 38335 15079
rect 8033 14977 8067 15011
rect 9781 14977 9815 15011
rect 13553 14977 13587 15011
rect 16313 14977 16347 15011
rect 20085 14977 20119 15011
rect 22201 14977 22235 15011
rect 23581 14977 23615 15011
rect 25053 14977 25087 15011
rect 26617 14977 26651 15011
rect 27169 14977 27203 15011
rect 27261 14977 27295 15011
rect 29009 14977 29043 15011
rect 29469 14977 29503 15011
rect 32321 14977 32355 15011
rect 32965 14977 32999 15011
rect 34161 14977 34195 15011
rect 35265 14977 35299 15011
rect 36093 14977 36127 15011
rect 36737 14977 36771 15011
rect 38117 14977 38151 15011
rect 14289 14909 14323 14943
rect 22293 14909 22327 14943
rect 23397 14909 23431 14943
rect 28365 14909 28399 14943
rect 28549 14909 28583 14943
rect 30757 14909 30791 14943
rect 31033 14909 31067 14943
rect 34345 14909 34379 14943
rect 36829 14909 36863 14943
rect 17141 14841 17175 14875
rect 33057 14841 33091 14875
rect 9873 14773 9907 14807
rect 24041 14773 24075 14807
rect 25145 14773 25179 14807
rect 32413 14773 32447 14807
rect 34529 14773 34563 14807
rect 1593 14569 1627 14603
rect 17693 14569 17727 14603
rect 20913 14569 20947 14603
rect 29837 14569 29871 14603
rect 33333 14569 33367 14603
rect 34253 14569 34287 14603
rect 34989 14501 35023 14535
rect 16037 14433 16071 14467
rect 17049 14433 17083 14467
rect 21557 14433 21591 14467
rect 32873 14433 32907 14467
rect 36553 14433 36587 14467
rect 37473 14433 37507 14467
rect 1777 14365 1811 14399
rect 9137 14365 9171 14399
rect 12265 14365 12299 14399
rect 14933 14365 14967 14399
rect 15025 14365 15059 14399
rect 20637 14365 20671 14399
rect 23029 14365 23063 14399
rect 23673 14365 23707 14399
rect 24593 14365 24627 14399
rect 29009 14365 29043 14399
rect 29745 14365 29779 14399
rect 31585 14365 31619 14399
rect 32689 14365 32723 14399
rect 34161 14365 34195 14399
rect 34897 14365 34931 14399
rect 36461 14365 36495 14399
rect 16129 14297 16163 14331
rect 17601 14297 17635 14331
rect 21649 14297 21683 14331
rect 22569 14297 22603 14331
rect 27537 14297 27571 14331
rect 27629 14297 27663 14331
rect 28549 14297 28583 14331
rect 30481 14297 30515 14331
rect 30573 14297 30607 14331
rect 31125 14297 31159 14331
rect 35817 14297 35851 14331
rect 37197 14297 37231 14331
rect 37289 14297 37323 14331
rect 9229 14229 9263 14263
rect 12357 14229 12391 14263
rect 23121 14229 23155 14263
rect 23765 14229 23799 14263
rect 24685 14229 24719 14263
rect 29101 14229 29135 14263
rect 31677 14229 31711 14263
rect 9321 14025 9355 14059
rect 14933 14025 14967 14059
rect 30205 14025 30239 14059
rect 32413 14025 32447 14059
rect 33793 14025 33827 14059
rect 34529 14025 34563 14059
rect 11897 13957 11931 13991
rect 17877 13957 17911 13991
rect 20637 13957 20671 13991
rect 22201 13957 22235 13991
rect 24777 13957 24811 13991
rect 28273 13957 28307 13991
rect 28825 13957 28859 13991
rect 35817 13957 35851 13991
rect 1593 13889 1627 13923
rect 8861 13889 8895 13923
rect 14289 13889 14323 13923
rect 18889 13889 18923 13923
rect 23581 13889 23615 13923
rect 29469 13889 29503 13923
rect 30113 13889 30147 13923
rect 31217 13889 31251 13923
rect 32597 13889 32631 13923
rect 33977 13889 34011 13923
rect 34713 13889 34747 13923
rect 38025 13889 38059 13923
rect 8677 13821 8711 13855
rect 11805 13821 11839 13855
rect 12081 13821 12115 13855
rect 14473 13821 14507 13855
rect 17785 13821 17819 13855
rect 18429 13821 18463 13855
rect 19993 13821 20027 13855
rect 20177 13821 20211 13855
rect 21281 13821 21315 13855
rect 22109 13821 22143 13855
rect 23121 13821 23155 13855
rect 23673 13821 23707 13855
rect 24685 13821 24719 13855
rect 24961 13821 24995 13855
rect 28181 13821 28215 13855
rect 31033 13821 31067 13855
rect 35725 13821 35759 13855
rect 36001 13821 36035 13855
rect 1777 13685 1811 13719
rect 18981 13685 19015 13719
rect 29285 13685 29319 13719
rect 31401 13685 31435 13719
rect 38209 13685 38243 13719
rect 14749 13481 14783 13515
rect 30389 13481 30423 13515
rect 34161 13481 34195 13515
rect 38209 13481 38243 13515
rect 23305 13413 23339 13447
rect 24593 13413 24627 13447
rect 28917 13413 28951 13447
rect 37565 13413 37599 13447
rect 10793 13345 10827 13379
rect 11069 13345 11103 13379
rect 16957 13345 16991 13379
rect 17233 13345 17267 13379
rect 19993 13345 20027 13379
rect 26341 13345 26375 13379
rect 26525 13345 26559 13379
rect 28733 13345 28767 13379
rect 29929 13345 29963 13379
rect 31217 13345 31251 13379
rect 31401 13345 31435 13379
rect 32413 13345 32447 13379
rect 14933 13277 14967 13311
rect 21557 13277 21591 13311
rect 22661 13277 22695 13311
rect 23489 13277 23523 13311
rect 24777 13277 24811 13311
rect 27905 13277 27939 13311
rect 28549 13277 28583 13311
rect 29745 13277 29779 13311
rect 32321 13277 32355 13311
rect 32965 13277 32999 13311
rect 34069 13277 34103 13311
rect 35081 13277 35115 13311
rect 38117 13277 38151 13311
rect 10885 13209 10919 13243
rect 17049 13209 17083 13243
rect 33057 13209 33091 13243
rect 37013 13209 37047 13243
rect 37105 13209 37139 13243
rect 21649 13141 21683 13175
rect 22753 13141 22787 13175
rect 26985 13141 27019 13175
rect 27997 13141 28031 13175
rect 31861 13141 31895 13175
rect 34897 13141 34931 13175
rect 35541 13141 35575 13175
rect 36185 13141 36219 13175
rect 28089 12937 28123 12971
rect 32597 12937 32631 12971
rect 33333 12937 33367 12971
rect 10609 12869 10643 12903
rect 12265 12869 12299 12903
rect 18337 12869 18371 12903
rect 23673 12869 23707 12903
rect 24225 12869 24259 12903
rect 25053 12869 25087 12903
rect 31585 12869 31619 12903
rect 34897 12869 34931 12903
rect 36185 12869 36219 12903
rect 36277 12869 36311 12903
rect 1593 12801 1627 12835
rect 4261 12801 4295 12835
rect 10517 12801 10551 12835
rect 12173 12801 12207 12835
rect 15025 12801 15059 12835
rect 19901 12801 19935 12835
rect 22201 12801 22235 12835
rect 25605 12801 25639 12835
rect 28273 12801 28307 12835
rect 29285 12801 29319 12835
rect 31401 12801 31435 12835
rect 32781 12801 32815 12835
rect 33241 12801 33275 12835
rect 34069 12801 34103 12835
rect 38025 12801 38059 12835
rect 18245 12733 18279 12767
rect 18889 12733 18923 12767
rect 22017 12733 22051 12767
rect 23581 12733 23615 12767
rect 24961 12733 24995 12767
rect 29101 12733 29135 12767
rect 30205 12733 30239 12767
rect 30389 12733 30423 12767
rect 34805 12733 34839 12767
rect 36461 12733 36495 12767
rect 14841 12665 14875 12699
rect 19717 12665 19751 12699
rect 22385 12665 22419 12699
rect 30849 12665 30883 12699
rect 35357 12665 35391 12699
rect 1777 12597 1811 12631
rect 4077 12597 4111 12631
rect 29469 12597 29503 12631
rect 34161 12597 34195 12631
rect 38209 12597 38243 12631
rect 4905 12393 4939 12427
rect 14381 12393 14415 12427
rect 19717 12393 19751 12427
rect 33885 12393 33919 12427
rect 37749 12393 37783 12427
rect 23949 12257 23983 12291
rect 29837 12257 29871 12291
rect 30481 12257 30515 12291
rect 31309 12257 31343 12291
rect 34989 12257 35023 12291
rect 35633 12257 35667 12291
rect 37013 12257 37047 12291
rect 4813 12189 4847 12223
rect 14289 12189 14323 12223
rect 19901 12189 19935 12223
rect 20361 12189 20395 12223
rect 32321 12189 32355 12223
rect 33425 12189 33459 12223
rect 34069 12189 34103 12223
rect 36921 12189 36955 12223
rect 37657 12189 37691 12223
rect 22937 12121 22971 12155
rect 23029 12121 23063 12155
rect 24685 12121 24719 12155
rect 24777 12121 24811 12155
rect 25697 12121 25731 12155
rect 29906 12121 29940 12155
rect 31033 12121 31067 12155
rect 31125 12121 31159 12155
rect 35081 12121 35115 12155
rect 20453 12053 20487 12087
rect 32137 12053 32171 12087
rect 33241 12053 33275 12087
rect 36093 12053 36127 12087
rect 12633 11849 12667 11883
rect 16221 11849 16255 11883
rect 29653 11849 29687 11883
rect 32965 11849 32999 11883
rect 36553 11849 36587 11883
rect 16957 11781 16991 11815
rect 17693 11781 17727 11815
rect 18613 11781 18647 11815
rect 20085 11781 20119 11815
rect 21005 11781 21039 11815
rect 25421 11781 25455 11815
rect 30849 11781 30883 11815
rect 31769 11781 31803 11815
rect 6929 11713 6963 11747
rect 12541 11713 12575 11747
rect 16129 11713 16163 11747
rect 16865 11713 16899 11747
rect 22017 11713 22051 11747
rect 22661 11713 22695 11747
rect 26433 11713 26467 11747
rect 29561 11713 29595 11747
rect 32321 11713 32355 11747
rect 33149 11713 33183 11747
rect 34805 11713 34839 11747
rect 35817 11713 35851 11747
rect 36461 11713 36495 11747
rect 37749 11713 37783 11747
rect 17601 11645 17635 11679
rect 19993 11645 20027 11679
rect 25329 11645 25363 11679
rect 30757 11645 30791 11679
rect 34621 11645 34655 11679
rect 35909 11645 35943 11679
rect 25881 11577 25915 11611
rect 34989 11577 35023 11611
rect 6745 11509 6779 11543
rect 22109 11509 22143 11543
rect 22753 11509 22787 11543
rect 26525 11509 26559 11543
rect 32413 11509 32447 11543
rect 37841 11509 37875 11543
rect 1777 11305 1811 11339
rect 9689 11305 9723 11339
rect 10793 11305 10827 11339
rect 19993 11305 20027 11339
rect 22293 11305 22327 11339
rect 29929 11305 29963 11339
rect 30757 11305 30791 11339
rect 7389 11237 7423 11271
rect 18429 11237 18463 11271
rect 21465 11237 21499 11271
rect 35541 11237 35575 11271
rect 6561 11169 6595 11203
rect 9321 11169 9355 11203
rect 21281 11169 21315 11203
rect 31309 11169 31343 11203
rect 37841 11169 37875 11203
rect 6469 11101 6503 11135
rect 7573 11101 7607 11135
rect 9137 11101 9171 11135
rect 10701 11101 10735 11135
rect 13277 11101 13311 11135
rect 15853 11101 15887 11135
rect 18337 11101 18371 11135
rect 21097 11101 21131 11135
rect 22201 11101 22235 11135
rect 30113 11101 30147 11135
rect 30665 11101 30699 11135
rect 34897 11101 34931 11135
rect 34989 11101 35023 11135
rect 35725 11101 35759 11135
rect 36829 11101 36863 11135
rect 1685 11033 1719 11067
rect 13461 11033 13495 11067
rect 19901 11033 19935 11067
rect 37013 11033 37047 11067
rect 37565 11033 37599 11067
rect 37657 11033 37691 11067
rect 15945 10965 15979 10999
rect 28917 10965 28951 10999
rect 1593 10761 1627 10795
rect 9137 10761 9171 10795
rect 20085 10761 20119 10795
rect 29561 10761 29595 10795
rect 36001 10761 36035 10795
rect 38209 10761 38243 10795
rect 27353 10693 27387 10727
rect 27905 10693 27939 10727
rect 1777 10625 1811 10659
rect 9045 10625 9079 10659
rect 14565 10625 14599 10659
rect 15209 10625 15243 10659
rect 15393 10625 15427 10659
rect 19993 10625 20027 10659
rect 22201 10625 22235 10659
rect 24133 10625 24167 10659
rect 28917 10625 28951 10659
rect 30021 10625 30055 10659
rect 36185 10625 36219 10659
rect 36921 10625 36955 10659
rect 38025 10625 38059 10659
rect 27261 10557 27295 10591
rect 29101 10557 29135 10591
rect 30113 10489 30147 10523
rect 14657 10421 14691 10455
rect 15853 10421 15887 10455
rect 22293 10421 22327 10455
rect 24225 10421 24259 10455
rect 36737 10421 36771 10455
rect 16129 10217 16163 10251
rect 27353 10217 27387 10251
rect 30481 10217 30515 10251
rect 36737 10217 36771 10251
rect 38209 10217 38243 10251
rect 25237 10149 25271 10183
rect 22569 10081 22603 10115
rect 24593 10081 24627 10115
rect 2237 10013 2271 10047
rect 12449 10013 12483 10047
rect 12633 10013 12667 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 17785 10013 17819 10047
rect 21465 10013 21499 10047
rect 24777 10013 24811 10047
rect 27261 10013 27295 10047
rect 30389 10013 30423 10047
rect 36921 10013 36955 10047
rect 37565 10013 37599 10047
rect 38025 10013 38059 10047
rect 22661 9945 22695 9979
rect 23581 9945 23615 9979
rect 2237 9877 2271 9911
rect 13093 9877 13127 9911
rect 17877 9877 17911 9911
rect 21557 9877 21591 9911
rect 37381 9877 37415 9911
rect 12449 9673 12483 9707
rect 13185 9673 13219 9707
rect 15761 9673 15795 9707
rect 29193 9673 29227 9707
rect 17049 9605 17083 9639
rect 21005 9605 21039 9639
rect 23489 9605 23523 9639
rect 24961 9605 24995 9639
rect 2053 9537 2087 9571
rect 13093 9537 13127 9571
rect 14657 9537 14691 9571
rect 15301 9537 15335 9571
rect 19901 9537 19935 9571
rect 22661 9537 22695 9571
rect 24869 9537 24903 9571
rect 29377 9537 29411 9571
rect 37933 9537 37967 9571
rect 16957 9469 16991 9503
rect 20361 9469 20395 9503
rect 20545 9469 20579 9503
rect 23397 9469 23431 9503
rect 14473 9401 14507 9435
rect 15117 9401 15151 9435
rect 17509 9401 17543 9435
rect 23949 9401 23983 9435
rect 37749 9401 37783 9435
rect 1869 9333 1903 9367
rect 19717 9333 19751 9367
rect 22753 9333 22787 9367
rect 14933 9129 14967 9163
rect 20177 9129 20211 9163
rect 22385 9129 22419 9163
rect 14473 8993 14507 9027
rect 25329 8993 25363 9027
rect 30573 8993 30607 9027
rect 37565 8993 37599 9027
rect 1593 8925 1627 8959
rect 14289 8925 14323 8959
rect 20361 8925 20395 8959
rect 22293 8925 22327 8959
rect 22937 8925 22971 8959
rect 27169 8925 27203 8959
rect 32965 8925 32999 8959
rect 23213 8857 23247 8891
rect 24685 8857 24719 8891
rect 24777 8857 24811 8891
rect 30113 8857 30147 8891
rect 30205 8857 30239 8891
rect 1777 8789 1811 8823
rect 27261 8789 27295 8823
rect 32781 8789 32815 8823
rect 10425 8585 10459 8619
rect 28917 8585 28951 8619
rect 30113 8585 30147 8619
rect 38117 8585 38151 8619
rect 22201 8517 22235 8551
rect 22753 8517 22787 8551
rect 27721 8517 27755 8551
rect 28273 8517 28307 8551
rect 10333 8449 10367 8483
rect 26433 8449 26467 8483
rect 29101 8449 29135 8483
rect 38301 8449 38335 8483
rect 21281 8381 21315 8415
rect 22109 8381 22143 8415
rect 27629 8381 27663 8415
rect 26525 8245 26559 8279
rect 1593 8041 1627 8075
rect 8309 8041 8343 8075
rect 31861 8041 31895 8075
rect 27721 7973 27755 8007
rect 31585 7973 31619 8007
rect 37749 7905 37783 7939
rect 1777 7837 1811 7871
rect 8217 7837 8251 7871
rect 21741 7837 21775 7871
rect 21833 7837 21867 7871
rect 23397 7837 23431 7871
rect 27721 7837 27755 7871
rect 32413 7837 32447 7871
rect 37473 7837 37507 7871
rect 31401 7769 31435 7803
rect 23213 7701 23247 7735
rect 32229 7701 32263 7735
rect 26617 7497 26651 7531
rect 38117 7497 38151 7531
rect 1777 7361 1811 7395
rect 20453 7361 20487 7395
rect 23765 7361 23799 7395
rect 25973 7361 26007 7395
rect 26157 7361 26191 7395
rect 38301 7361 38335 7395
rect 1593 7157 1627 7191
rect 20269 7157 20303 7191
rect 23581 7157 23615 7191
rect 9229 6817 9263 6851
rect 24041 6817 24075 6851
rect 31493 6817 31527 6851
rect 9137 6749 9171 6783
rect 23397 6749 23431 6783
rect 23581 6749 23615 6783
rect 24777 6749 24811 6783
rect 29745 6749 29779 6783
rect 30481 6681 30515 6715
rect 30573 6681 30607 6715
rect 24593 6613 24627 6647
rect 29837 6613 29871 6647
rect 14933 6273 14967 6307
rect 24501 6273 24535 6307
rect 30481 6273 30515 6307
rect 15025 6069 15059 6103
rect 24593 6069 24627 6103
rect 30297 6069 30331 6103
rect 1593 5865 1627 5899
rect 1777 5661 1811 5695
rect 26341 5661 26375 5695
rect 38025 5661 38059 5695
rect 37657 5593 37691 5627
rect 26157 5525 26191 5559
rect 38209 5525 38243 5559
rect 22661 5321 22695 5355
rect 23949 5321 23983 5355
rect 29469 5321 29503 5355
rect 22569 5185 22603 5219
rect 23857 5185 23891 5219
rect 29377 5185 29411 5219
rect 37749 4641 37783 4675
rect 1593 4573 1627 4607
rect 2237 4573 2271 4607
rect 37473 4573 37507 4607
rect 1777 4437 1811 4471
rect 38025 4097 38059 4131
rect 37841 3893 37875 3927
rect 36737 3689 36771 3723
rect 1593 3485 1627 3519
rect 36921 3485 36955 3519
rect 37565 3485 37599 3519
rect 38025 3485 38059 3519
rect 1777 3349 1811 3383
rect 37381 3349 37415 3383
rect 38209 3349 38243 3383
rect 2329 3145 2363 3179
rect 3985 3145 4019 3179
rect 22661 3145 22695 3179
rect 35265 3145 35299 3179
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3157 3009 3191 3043
rect 4169 3009 4203 3043
rect 5549 3009 5583 3043
rect 13277 3009 13311 3043
rect 17049 3009 17083 3043
rect 22845 3009 22879 3043
rect 30389 3009 30423 3043
rect 35449 3009 35483 3043
rect 35909 3009 35943 3043
rect 36001 3009 36035 3043
rect 36921 3009 36955 3043
rect 38025 3009 38059 3043
rect 2973 2873 3007 2907
rect 13093 2873 13127 2907
rect 16865 2873 16899 2907
rect 36737 2873 36771 2907
rect 1777 2805 1811 2839
rect 5365 2805 5399 2839
rect 30573 2805 30607 2839
rect 38209 2805 38243 2839
rect 10425 2601 10459 2635
rect 11713 2601 11747 2635
rect 14289 2601 14323 2635
rect 18153 2601 18187 2635
rect 19441 2601 19475 2635
rect 22017 2601 22051 2635
rect 24593 2601 24627 2635
rect 27169 2601 27203 2635
rect 2973 2533 3007 2567
rect 7297 2533 7331 2567
rect 9781 2533 9815 2567
rect 20085 2533 20119 2567
rect 13185 2465 13219 2499
rect 15209 2465 15243 2499
rect 17141 2465 17175 2499
rect 31217 2465 31251 2499
rect 32597 2465 32631 2499
rect 2053 2397 2087 2431
rect 2789 2397 2823 2431
rect 3985 2397 4019 2431
rect 5273 2397 5307 2431
rect 6561 2397 6595 2431
rect 7481 2397 7515 2431
rect 9321 2397 9355 2431
rect 9965 2397 9999 2431
rect 10609 2397 10643 2431
rect 11897 2397 11931 2431
rect 12909 2397 12943 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 16865 2397 16899 2431
rect 18337 2397 18371 2431
rect 19625 2397 19659 2431
rect 20269 2397 20303 2431
rect 22201 2397 22235 2431
rect 23213 2397 23247 2431
rect 23489 2397 23523 2431
rect 24777 2397 24811 2431
rect 26065 2397 26099 2431
rect 27353 2397 27387 2431
rect 27813 2397 27847 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 32321 2397 32355 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 35909 2397 35943 2431
rect 36645 2397 36679 2431
rect 37473 2397 37507 2431
rect 38025 2397 38059 2431
rect 2237 2261 2271 2295
rect 4169 2261 4203 2295
rect 5457 2261 5491 2295
rect 6745 2261 6779 2295
rect 9137 2261 9171 2295
rect 25881 2261 25915 2295
rect 27997 2261 28031 2295
rect 29929 2261 29963 2295
rect 33793 2261 33827 2295
rect 35081 2261 35115 2295
rect 36093 2261 36127 2295
rect 36829 2261 36863 2295
rect 37657 2261 37691 2295
<< metal1 >>
rect 2866 38292 2872 38344
rect 2924 38332 2930 38344
rect 4614 38332 4620 38344
rect 2924 38304 4620 38332
rect 2924 38292 2930 38304
rect 4614 38292 4620 38304
rect 4672 38292 4678 38344
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 12529 37451 12587 37457
rect 12529 37417 12541 37451
rect 12575 37448 12587 37451
rect 14734 37448 14740 37460
rect 12575 37420 14740 37448
rect 12575 37417 12587 37420
rect 12529 37411 12587 37417
rect 14734 37408 14740 37420
rect 14792 37408 14798 37460
rect 17770 37408 17776 37460
rect 17828 37448 17834 37460
rect 17957 37451 18015 37457
rect 17957 37448 17969 37451
rect 17828 37420 17969 37448
rect 17828 37408 17834 37420
rect 17957 37417 17969 37420
rect 18003 37417 18015 37451
rect 17957 37411 18015 37417
rect 30926 37408 30932 37460
rect 30984 37448 30990 37460
rect 32493 37451 32551 37457
rect 32493 37448 32505 37451
rect 30984 37420 32505 37448
rect 30984 37408 30990 37420
rect 32493 37417 32505 37420
rect 32539 37417 32551 37451
rect 32493 37411 32551 37417
rect 13541 37383 13599 37389
rect 13541 37349 13553 37383
rect 13587 37349 13599 37383
rect 13541 37343 13599 37349
rect 14553 37383 14611 37389
rect 14553 37349 14565 37383
rect 14599 37380 14611 37383
rect 17862 37380 17868 37392
rect 14599 37352 17868 37380
rect 14599 37349 14611 37352
rect 14553 37343 14611 37349
rect 1946 37272 1952 37324
rect 2004 37312 2010 37324
rect 2041 37315 2099 37321
rect 2041 37312 2053 37315
rect 2004 37284 2053 37312
rect 2004 37272 2010 37284
rect 2041 37281 2053 37284
rect 2087 37281 2099 37315
rect 2041 37275 2099 37281
rect 4249 37315 4307 37321
rect 4249 37281 4261 37315
rect 4295 37312 4307 37315
rect 4890 37312 4896 37324
rect 4295 37284 4896 37312
rect 4295 37281 4307 37284
rect 4249 37275 4307 37281
rect 4890 37272 4896 37284
rect 4948 37272 4954 37324
rect 8386 37272 8392 37324
rect 8444 37312 8450 37324
rect 9125 37315 9183 37321
rect 9125 37312 9137 37315
rect 8444 37284 9137 37312
rect 8444 37272 8450 37284
rect 9125 37281 9137 37284
rect 9171 37281 9183 37315
rect 13556 37312 13584 37343
rect 17862 37340 17868 37352
rect 17920 37340 17926 37392
rect 18138 37340 18144 37392
rect 18196 37380 18202 37392
rect 18966 37380 18972 37392
rect 18196 37352 18972 37380
rect 18196 37340 18202 37352
rect 18966 37340 18972 37352
rect 19024 37340 19030 37392
rect 28166 37340 28172 37392
rect 28224 37380 28230 37392
rect 28537 37383 28595 37389
rect 28537 37380 28549 37383
rect 28224 37352 28549 37380
rect 28224 37340 28230 37352
rect 28537 37349 28549 37352
rect 28583 37349 28595 37383
rect 28537 37343 28595 37349
rect 9125 37275 9183 37281
rect 11624 37284 12572 37312
rect 13556 37284 19334 37312
rect 2130 37204 2136 37256
rect 2188 37244 2194 37256
rect 2317 37247 2375 37253
rect 2317 37244 2329 37247
rect 2188 37216 2329 37244
rect 2188 37204 2194 37216
rect 2317 37213 2329 37216
rect 2363 37213 2375 37247
rect 2317 37207 2375 37213
rect 3418 37204 3424 37256
rect 3476 37244 3482 37256
rect 4065 37247 4123 37253
rect 4065 37244 4077 37247
rect 3476 37216 4077 37244
rect 3476 37204 3482 37216
rect 4065 37213 4077 37216
rect 4111 37213 4123 37247
rect 4065 37207 4123 37213
rect 5166 37204 5172 37256
rect 5224 37244 5230 37256
rect 5445 37247 5503 37253
rect 5445 37244 5457 37247
rect 5224 37216 5457 37244
rect 5224 37204 5230 37216
rect 5445 37213 5457 37216
rect 5491 37213 5503 37247
rect 5445 37207 5503 37213
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 6733 37247 6791 37253
rect 6733 37244 6745 37247
rect 5868 37216 6745 37244
rect 5868 37204 5874 37216
rect 6733 37213 6745 37216
rect 6779 37213 6791 37247
rect 6733 37207 6791 37213
rect 7098 37204 7104 37256
rect 7156 37244 7162 37256
rect 7377 37247 7435 37253
rect 7377 37244 7389 37247
rect 7156 37216 7389 37244
rect 7156 37204 7162 37216
rect 7377 37213 7389 37216
rect 7423 37213 7435 37247
rect 7377 37207 7435 37213
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37244 8631 37247
rect 9030 37244 9036 37256
rect 8619 37216 9036 37244
rect 8619 37213 8631 37216
rect 8573 37207 8631 37213
rect 9030 37204 9036 37216
rect 9088 37204 9094 37256
rect 9401 37247 9459 37253
rect 9401 37213 9413 37247
rect 9447 37244 9459 37247
rect 9490 37244 9496 37256
rect 9447 37216 9496 37244
rect 9447 37213 9459 37216
rect 9401 37207 9459 37213
rect 9490 37204 9496 37216
rect 9548 37204 9554 37256
rect 10413 37247 10471 37253
rect 10413 37213 10425 37247
rect 10459 37244 10471 37247
rect 11624 37244 11652 37284
rect 10459 37216 11652 37244
rect 11701 37247 11759 37253
rect 10459 37213 10471 37216
rect 10413 37207 10471 37213
rect 11701 37213 11713 37247
rect 11747 37213 11759 37247
rect 11701 37207 11759 37213
rect 8110 37136 8116 37188
rect 8168 37176 8174 37188
rect 10042 37176 10048 37188
rect 8168 37148 10048 37176
rect 8168 37136 8174 37148
rect 10042 37136 10048 37148
rect 10100 37136 10106 37188
rect 11054 37176 11060 37188
rect 10244 37148 11060 37176
rect 5261 37111 5319 37117
rect 5261 37077 5273 37111
rect 5307 37108 5319 37111
rect 6362 37108 6368 37120
rect 5307 37080 6368 37108
rect 5307 37077 5319 37080
rect 5261 37071 5319 37077
rect 6362 37068 6368 37080
rect 6420 37068 6426 37120
rect 6549 37111 6607 37117
rect 6549 37077 6561 37111
rect 6595 37108 6607 37111
rect 6638 37108 6644 37120
rect 6595 37080 6644 37108
rect 6595 37077 6607 37080
rect 6549 37071 6607 37077
rect 6638 37068 6644 37080
rect 6696 37068 6702 37120
rect 7190 37108 7196 37120
rect 7151 37080 7196 37108
rect 7190 37068 7196 37080
rect 7248 37068 7254 37120
rect 8389 37111 8447 37117
rect 8389 37077 8401 37111
rect 8435 37108 8447 37111
rect 9122 37108 9128 37120
rect 8435 37080 9128 37108
rect 8435 37077 8447 37080
rect 8389 37071 8447 37077
rect 9122 37068 9128 37080
rect 9180 37068 9186 37120
rect 9766 37068 9772 37120
rect 9824 37108 9830 37120
rect 10244 37108 10272 37148
rect 11054 37136 11060 37148
rect 11112 37136 11118 37188
rect 11716 37176 11744 37207
rect 12250 37204 12256 37256
rect 12308 37244 12314 37256
rect 12437 37247 12495 37253
rect 12437 37244 12449 37247
rect 12308 37216 12449 37244
rect 12308 37204 12314 37216
rect 12437 37213 12449 37216
rect 12483 37213 12495 37247
rect 12544 37244 12572 37284
rect 13630 37244 13636 37256
rect 12544 37216 13636 37244
rect 12437 37207 12495 37213
rect 13630 37204 13636 37216
rect 13688 37204 13694 37256
rect 13725 37247 13783 37253
rect 13725 37213 13737 37247
rect 13771 37213 13783 37247
rect 13725 37207 13783 37213
rect 13740 37176 13768 37207
rect 13814 37204 13820 37256
rect 13872 37244 13878 37256
rect 14369 37247 14427 37253
rect 14369 37244 14381 37247
rect 13872 37216 14381 37244
rect 13872 37204 13878 37216
rect 14369 37213 14381 37216
rect 14415 37213 14427 37247
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 14369 37207 14427 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 15286 37204 15292 37256
rect 15344 37244 15350 37256
rect 16025 37247 16083 37253
rect 16025 37244 16037 37247
rect 15344 37216 16037 37244
rect 15344 37204 15350 37216
rect 16025 37213 16037 37216
rect 16071 37213 16083 37247
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16025 37207 16083 37213
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 18141 37247 18199 37253
rect 18141 37213 18153 37247
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 15930 37176 15936 37188
rect 11716 37148 12434 37176
rect 13740 37148 15936 37176
rect 9824 37080 10272 37108
rect 9824 37068 9830 37080
rect 10318 37068 10324 37120
rect 10376 37108 10382 37120
rect 10597 37111 10655 37117
rect 10597 37108 10609 37111
rect 10376 37080 10609 37108
rect 10376 37068 10382 37080
rect 10597 37077 10609 37080
rect 10643 37077 10655 37111
rect 10597 37071 10655 37077
rect 11330 37068 11336 37120
rect 11388 37108 11394 37120
rect 11793 37111 11851 37117
rect 11793 37108 11805 37111
rect 11388 37080 11805 37108
rect 11388 37068 11394 37080
rect 11793 37077 11805 37080
rect 11839 37077 11851 37111
rect 12406 37108 12434 37148
rect 15930 37136 15936 37148
rect 15988 37136 15994 37188
rect 18156 37176 18184 37207
rect 18230 37204 18236 37256
rect 18288 37244 18294 37256
rect 18601 37247 18659 37253
rect 18601 37244 18613 37247
rect 18288 37216 18613 37244
rect 18288 37204 18294 37216
rect 18601 37213 18613 37216
rect 18647 37213 18659 37247
rect 19306 37244 19334 37284
rect 22738 37272 22744 37324
rect 22796 37312 22802 37324
rect 23017 37315 23075 37321
rect 23017 37312 23029 37315
rect 22796 37284 23029 37312
rect 22796 37272 22802 37284
rect 23017 37281 23029 37284
rect 23063 37281 23075 37315
rect 25774 37312 25780 37324
rect 25735 37284 25780 37312
rect 23017 37275 23075 37281
rect 25774 37272 25780 37284
rect 25832 37272 25838 37324
rect 28000 37284 28304 37312
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 19306 37216 20085 37244
rect 18601 37207 18659 37213
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 20073 37207 20131 37213
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 21993 37247 22051 37253
rect 21993 37244 22005 37247
rect 20588 37216 22005 37244
rect 20588 37204 20594 37216
rect 21993 37213 22005 37216
rect 22039 37213 22051 37247
rect 21993 37207 22051 37213
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22612 37216 22845 37244
rect 22612 37204 22618 37216
rect 22833 37213 22845 37216
rect 22879 37213 22891 37247
rect 23474 37244 23480 37256
rect 23435 37216 23480 37244
rect 22833 37207 22891 37213
rect 23474 37204 23480 37216
rect 23532 37204 23538 37256
rect 24486 37204 24492 37256
rect 24544 37244 24550 37256
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 24544 37216 24777 37244
rect 24544 37204 24550 37216
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 26050 37244 26056 37256
rect 26011 37216 26056 37244
rect 24765 37207 24823 37213
rect 26050 37204 26056 37216
rect 26108 37204 26114 37256
rect 27157 37247 27215 37253
rect 27157 37213 27169 37247
rect 27203 37244 27215 37247
rect 27203 37216 27476 37244
rect 27203 37213 27215 37216
rect 27157 37207 27215 37213
rect 18322 37176 18328 37188
rect 18156 37148 18328 37176
rect 18322 37136 18328 37148
rect 18380 37136 18386 37188
rect 18874 37136 18880 37188
rect 18932 37176 18938 37188
rect 18932 37148 24624 37176
rect 18932 37136 18938 37148
rect 14918 37108 14924 37120
rect 12406 37080 14924 37108
rect 11793 37071 11851 37077
rect 14918 37068 14924 37080
rect 14976 37068 14982 37120
rect 15010 37068 15016 37120
rect 15068 37108 15074 37120
rect 15068 37080 15113 37108
rect 15068 37068 15074 37080
rect 16114 37068 16120 37120
rect 16172 37108 16178 37120
rect 16209 37111 16267 37117
rect 16209 37108 16221 37111
rect 16172 37080 16221 37108
rect 16172 37068 16178 37080
rect 16209 37077 16221 37080
rect 16255 37077 16267 37111
rect 16209 37071 16267 37077
rect 16758 37068 16764 37120
rect 16816 37108 16822 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 16816 37080 17049 37108
rect 16816 37068 16822 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 18785 37111 18843 37117
rect 18785 37077 18797 37111
rect 18831 37108 18843 37111
rect 19334 37108 19340 37120
rect 18831 37080 19340 37108
rect 18831 37077 18843 37080
rect 18785 37071 18843 37077
rect 19334 37068 19340 37080
rect 19392 37068 19398 37120
rect 19978 37068 19984 37120
rect 20036 37108 20042 37120
rect 20257 37111 20315 37117
rect 20257 37108 20269 37111
rect 20036 37080 20269 37108
rect 20036 37068 20042 37080
rect 20257 37077 20269 37080
rect 20303 37077 20315 37111
rect 20257 37071 20315 37077
rect 21266 37068 21272 37120
rect 21324 37108 21330 37120
rect 22189 37111 22247 37117
rect 22189 37108 22201 37111
rect 21324 37080 22201 37108
rect 21324 37068 21330 37080
rect 22189 37077 22201 37080
rect 22235 37077 22247 37111
rect 22189 37071 22247 37077
rect 23198 37068 23204 37120
rect 23256 37108 23262 37120
rect 24596 37117 24624 37148
rect 23661 37111 23719 37117
rect 23661 37108 23673 37111
rect 23256 37080 23673 37108
rect 23256 37068 23262 37080
rect 23661 37077 23673 37080
rect 23707 37077 23719 37111
rect 23661 37071 23719 37077
rect 24581 37111 24639 37117
rect 24581 37077 24593 37111
rect 24627 37077 24639 37111
rect 24581 37071 24639 37077
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27341 37111 27399 37117
rect 27341 37108 27353 37111
rect 26476 37080 27353 37108
rect 26476 37068 26482 37080
rect 27341 37077 27353 37080
rect 27387 37077 27399 37111
rect 27448 37108 27476 37216
rect 27706 37204 27712 37256
rect 27764 37244 27770 37256
rect 28000 37244 28028 37284
rect 27764 37216 28028 37244
rect 27764 37204 27770 37216
rect 28074 37204 28080 37256
rect 28132 37244 28138 37256
rect 28276 37244 28304 37284
rect 29086 37272 29092 37324
rect 29144 37312 29150 37324
rect 30285 37315 30343 37321
rect 30285 37312 30297 37315
rect 29144 37284 30297 37312
rect 29144 37272 29150 37284
rect 30285 37281 30297 37284
rect 30331 37281 30343 37315
rect 37461 37315 37519 37321
rect 30285 37275 30343 37281
rect 31312 37284 33640 37312
rect 31312 37256 31340 37284
rect 28721 37247 28779 37253
rect 28721 37244 28733 37247
rect 28132 37216 28177 37244
rect 28276 37216 28733 37244
rect 28132 37204 28138 37216
rect 28721 37213 28733 37216
rect 28767 37213 28779 37247
rect 28721 37207 28779 37213
rect 30009 37247 30067 37253
rect 30009 37213 30021 37247
rect 30055 37213 30067 37247
rect 30009 37207 30067 37213
rect 27522 37136 27528 37188
rect 27580 37176 27586 37188
rect 30024 37176 30052 37207
rect 31294 37204 31300 37256
rect 31352 37204 31358 37256
rect 31570 37204 31576 37256
rect 31628 37244 31634 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 31628 37216 32321 37244
rect 31628 37204 31634 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 32309 37207 32367 37213
rect 32950 37204 32956 37256
rect 33008 37244 33014 37256
rect 33045 37247 33103 37253
rect 33045 37244 33057 37247
rect 33008 37216 33057 37244
rect 33008 37204 33014 37216
rect 33045 37213 33057 37216
rect 33091 37213 33103 37247
rect 33045 37207 33103 37213
rect 27580 37148 28028 37176
rect 27580 37136 27586 37148
rect 27893 37111 27951 37117
rect 27893 37108 27905 37111
rect 27448 37080 27905 37108
rect 27341 37071 27399 37077
rect 27893 37077 27905 37080
rect 27939 37077 27951 37111
rect 28000 37108 28028 37148
rect 28276 37148 30052 37176
rect 28276 37108 28304 37148
rect 28000 37080 28304 37108
rect 30024 37108 30052 37148
rect 30374 37136 30380 37188
rect 30432 37176 30438 37188
rect 30432 37148 30696 37176
rect 30432 37136 30438 37148
rect 30466 37108 30472 37120
rect 30024 37080 30472 37108
rect 27893 37071 27951 37077
rect 30466 37068 30472 37080
rect 30524 37068 30530 37120
rect 30668 37108 30696 37148
rect 30742 37136 30748 37188
rect 30800 37136 30806 37188
rect 33502 37176 33508 37188
rect 33060 37148 33508 37176
rect 31662 37108 31668 37120
rect 30668 37080 31668 37108
rect 31662 37068 31668 37080
rect 31720 37068 31726 37120
rect 31757 37111 31815 37117
rect 31757 37077 31769 37111
rect 31803 37108 31815 37111
rect 33060 37108 33088 37148
rect 33502 37136 33508 37148
rect 33560 37136 33566 37188
rect 33612 37176 33640 37284
rect 37461 37281 37473 37315
rect 37507 37312 37519 37315
rect 38654 37312 38660 37324
rect 37507 37284 38660 37312
rect 37507 37281 37519 37284
rect 37461 37275 37519 37281
rect 38654 37272 38660 37284
rect 38712 37272 38718 37324
rect 33686 37204 33692 37256
rect 33744 37244 33750 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 33744 37216 34897 37244
rect 33744 37204 33750 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 36170 37244 36176 37256
rect 36131 37216 36176 37244
rect 34885 37207 34943 37213
rect 36170 37204 36176 37216
rect 36228 37204 36234 37256
rect 37737 37247 37795 37253
rect 37737 37213 37749 37247
rect 37783 37213 37795 37247
rect 37737 37207 37795 37213
rect 37752 37176 37780 37207
rect 33612 37148 37780 37176
rect 31803 37080 33088 37108
rect 31803 37077 31815 37080
rect 31757 37071 31815 37077
rect 33134 37068 33140 37120
rect 33192 37108 33198 37120
rect 33229 37111 33287 37117
rect 33229 37108 33241 37111
rect 33192 37080 33241 37108
rect 33192 37068 33198 37080
rect 33229 37077 33241 37080
rect 33275 37077 33287 37111
rect 33229 37071 33287 37077
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 35069 37111 35127 37117
rect 35069 37108 35081 37111
rect 34572 37080 35081 37108
rect 34572 37068 34578 37080
rect 35069 37077 35081 37080
rect 35115 37077 35127 37111
rect 35069 37071 35127 37077
rect 36078 37068 36084 37120
rect 36136 37108 36142 37120
rect 36357 37111 36415 37117
rect 36357 37108 36369 37111
rect 36136 37080 36369 37108
rect 36136 37068 36142 37080
rect 36357 37077 36369 37080
rect 36403 37077 36415 37111
rect 36357 37071 36415 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 3973 36907 4031 36913
rect 3973 36873 3985 36907
rect 4019 36904 4031 36907
rect 4019 36876 14872 36904
rect 4019 36873 4031 36876
rect 3973 36867 4031 36873
rect 1765 36839 1823 36845
rect 1765 36805 1777 36839
rect 1811 36836 1823 36839
rect 2222 36836 2228 36848
rect 1811 36808 2228 36836
rect 1811 36805 1823 36808
rect 1765 36799 1823 36805
rect 2222 36796 2228 36808
rect 2280 36796 2286 36848
rect 7469 36839 7527 36845
rect 7469 36805 7481 36839
rect 7515 36836 7527 36839
rect 9766 36836 9772 36848
rect 7515 36808 9772 36836
rect 7515 36805 7527 36808
rect 7469 36799 7527 36805
rect 9766 36796 9772 36808
rect 9824 36796 9830 36848
rect 9858 36796 9864 36848
rect 9916 36836 9922 36848
rect 9916 36808 9988 36836
rect 9916 36796 9922 36808
rect 2774 36728 2780 36780
rect 2832 36768 2838 36780
rect 3329 36771 3387 36777
rect 3329 36768 3341 36771
rect 2832 36740 3341 36768
rect 2832 36728 2838 36740
rect 3329 36737 3341 36740
rect 3375 36737 3387 36771
rect 4154 36768 4160 36780
rect 4115 36740 4160 36768
rect 3329 36731 3387 36737
rect 4154 36728 4160 36740
rect 4212 36728 4218 36780
rect 4801 36771 4859 36777
rect 4801 36737 4813 36771
rect 4847 36768 4859 36771
rect 7190 36768 7196 36780
rect 4847 36740 7196 36768
rect 4847 36737 4859 36740
rect 4801 36731 4859 36737
rect 7190 36728 7196 36740
rect 7248 36728 7254 36780
rect 7377 36771 7435 36777
rect 7377 36737 7389 36771
rect 7423 36768 7435 36771
rect 8110 36768 8116 36780
rect 7423 36740 8116 36768
rect 7423 36737 7435 36740
rect 7377 36731 7435 36737
rect 8110 36728 8116 36740
rect 8168 36728 8174 36780
rect 8205 36771 8263 36777
rect 8205 36737 8217 36771
rect 8251 36768 8263 36771
rect 8478 36768 8484 36780
rect 8251 36740 8484 36768
rect 8251 36737 8263 36740
rect 8205 36731 8263 36737
rect 8478 36728 8484 36740
rect 8536 36728 8542 36780
rect 8662 36768 8668 36780
rect 8623 36740 8668 36768
rect 8662 36728 8668 36740
rect 8720 36728 8726 36780
rect 9309 36771 9367 36777
rect 9309 36737 9321 36771
rect 9355 36768 9367 36771
rect 9674 36768 9680 36780
rect 9355 36740 9680 36768
rect 9355 36737 9367 36740
rect 9309 36731 9367 36737
rect 9674 36728 9680 36740
rect 9732 36728 9738 36780
rect 9960 36777 9988 36808
rect 11606 36796 11612 36848
rect 11664 36836 11670 36848
rect 11793 36839 11851 36845
rect 11793 36836 11805 36839
rect 11664 36808 11805 36836
rect 11664 36796 11670 36808
rect 11793 36805 11805 36808
rect 11839 36805 11851 36839
rect 11793 36799 11851 36805
rect 9953 36771 10011 36777
rect 9953 36737 9965 36771
rect 9999 36737 10011 36771
rect 10594 36768 10600 36780
rect 10555 36740 10600 36768
rect 9953 36731 10011 36737
rect 10594 36728 10600 36740
rect 10652 36728 10658 36780
rect 12618 36768 12624 36780
rect 10704 36740 12624 36768
rect 1673 36703 1731 36709
rect 1673 36700 1685 36703
rect 1596 36672 1685 36700
rect 1596 36644 1624 36672
rect 1673 36669 1685 36672
rect 1719 36669 1731 36703
rect 1673 36663 1731 36669
rect 2685 36703 2743 36709
rect 2685 36669 2697 36703
rect 2731 36700 2743 36703
rect 10704 36700 10732 36740
rect 12618 36728 12624 36740
rect 12676 36728 12682 36780
rect 12820 36777 12848 36876
rect 13633 36839 13691 36845
rect 13633 36805 13645 36839
rect 13679 36836 13691 36839
rect 13679 36808 14780 36836
rect 13679 36805 13691 36808
rect 13633 36799 13691 36805
rect 12805 36771 12863 36777
rect 12805 36737 12817 36771
rect 12851 36737 12863 36771
rect 12805 36731 12863 36737
rect 2731 36672 10732 36700
rect 2731 36669 2743 36672
rect 2685 36663 2743 36669
rect 11054 36660 11060 36712
rect 11112 36700 11118 36712
rect 11112 36672 12112 36700
rect 11112 36660 11118 36672
rect 1578 36592 1584 36644
rect 1636 36592 1642 36644
rect 4893 36635 4951 36641
rect 4893 36601 4905 36635
rect 4939 36632 4951 36635
rect 8018 36632 8024 36644
rect 4939 36604 7880 36632
rect 7979 36604 8024 36632
rect 4939 36601 4951 36604
rect 4893 36595 4951 36601
rect 2774 36524 2780 36576
rect 2832 36564 2838 36576
rect 3145 36567 3203 36573
rect 3145 36564 3157 36567
rect 2832 36536 3157 36564
rect 2832 36524 2838 36536
rect 3145 36533 3157 36536
rect 3191 36533 3203 36567
rect 7852 36564 7880 36604
rect 8018 36592 8024 36604
rect 8076 36592 8082 36644
rect 8757 36635 8815 36641
rect 8757 36601 8769 36635
rect 8803 36632 8815 36635
rect 11974 36632 11980 36644
rect 8803 36604 11980 36632
rect 8803 36601 8815 36604
rect 8757 36595 8815 36601
rect 11974 36592 11980 36604
rect 12032 36592 12038 36644
rect 12084 36632 12112 36672
rect 12158 36660 12164 36712
rect 12216 36700 12222 36712
rect 13541 36703 13599 36709
rect 13541 36700 13553 36703
rect 12216 36672 13553 36700
rect 12216 36660 12222 36672
rect 13541 36669 13553 36672
rect 13587 36669 13599 36703
rect 13541 36663 13599 36669
rect 13630 36660 13636 36712
rect 13688 36700 13694 36712
rect 14752 36700 14780 36808
rect 14844 36777 14872 36876
rect 14918 36864 14924 36916
rect 14976 36904 14982 36916
rect 17770 36904 17776 36916
rect 14976 36876 17776 36904
rect 14976 36864 14982 36876
rect 17770 36864 17776 36876
rect 17828 36864 17834 36916
rect 18046 36864 18052 36916
rect 18104 36864 18110 36916
rect 26602 36904 26608 36916
rect 22066 36876 26608 36904
rect 15654 36796 15660 36848
rect 15712 36836 15718 36848
rect 17862 36836 17868 36848
rect 15712 36808 17868 36836
rect 15712 36796 15718 36808
rect 17862 36796 17868 36808
rect 17920 36796 17926 36848
rect 17957 36839 18015 36845
rect 17957 36805 17969 36839
rect 18003 36836 18015 36839
rect 18064 36836 18092 36864
rect 18003 36808 18092 36836
rect 18003 36805 18015 36808
rect 17957 36799 18015 36805
rect 18414 36796 18420 36848
rect 18472 36796 18478 36848
rect 14829 36771 14887 36777
rect 14829 36737 14841 36771
rect 14875 36737 14887 36771
rect 15746 36768 15752 36780
rect 15707 36740 15752 36768
rect 14829 36731 14887 36737
rect 15746 36728 15752 36740
rect 15804 36728 15810 36780
rect 15841 36703 15899 36709
rect 15841 36700 15853 36703
rect 13688 36672 14688 36700
rect 14752 36672 15853 36700
rect 13688 36660 13694 36672
rect 12250 36632 12256 36644
rect 12084 36604 12256 36632
rect 12250 36592 12256 36604
rect 12308 36592 12314 36644
rect 12986 36592 12992 36644
rect 13044 36632 13050 36644
rect 14093 36635 14151 36641
rect 13044 36604 13308 36632
rect 13044 36592 13050 36604
rect 9306 36564 9312 36576
rect 7852 36536 9312 36564
rect 3145 36527 3203 36533
rect 9306 36524 9312 36536
rect 9364 36524 9370 36576
rect 9398 36524 9404 36576
rect 9456 36564 9462 36576
rect 10045 36567 10103 36573
rect 9456 36536 9501 36564
rect 9456 36524 9462 36536
rect 10045 36533 10057 36567
rect 10091 36564 10103 36567
rect 10502 36564 10508 36576
rect 10091 36536 10508 36564
rect 10091 36533 10103 36536
rect 10045 36527 10103 36533
rect 10502 36524 10508 36536
rect 10560 36524 10566 36576
rect 10689 36567 10747 36573
rect 10689 36533 10701 36567
rect 10735 36564 10747 36567
rect 11422 36564 11428 36576
rect 10735 36536 11428 36564
rect 10735 36533 10747 36536
rect 10689 36527 10747 36533
rect 11422 36524 11428 36536
rect 11480 36524 11486 36576
rect 11606 36524 11612 36576
rect 11664 36564 11670 36576
rect 11885 36567 11943 36573
rect 11885 36564 11897 36567
rect 11664 36536 11897 36564
rect 11664 36524 11670 36536
rect 11885 36533 11897 36536
rect 11931 36533 11943 36567
rect 11885 36527 11943 36533
rect 12897 36567 12955 36573
rect 12897 36533 12909 36567
rect 12943 36564 12955 36567
rect 13170 36564 13176 36576
rect 12943 36536 13176 36564
rect 12943 36533 12955 36536
rect 12897 36527 12955 36533
rect 13170 36524 13176 36536
rect 13228 36524 13234 36576
rect 13280 36564 13308 36604
rect 14093 36601 14105 36635
rect 14139 36632 14151 36635
rect 14366 36632 14372 36644
rect 14139 36604 14372 36632
rect 14139 36601 14151 36604
rect 14093 36595 14151 36601
rect 14366 36592 14372 36604
rect 14424 36592 14430 36644
rect 14660 36641 14688 36672
rect 15841 36669 15853 36672
rect 15887 36669 15899 36703
rect 15841 36663 15899 36669
rect 16850 36660 16856 36712
rect 16908 36700 16914 36712
rect 17681 36703 17739 36709
rect 17681 36700 17693 36703
rect 16908 36672 17693 36700
rect 16908 36660 16914 36672
rect 17681 36669 17693 36672
rect 17727 36669 17739 36703
rect 17681 36663 17739 36669
rect 14645 36635 14703 36641
rect 14645 36601 14657 36635
rect 14691 36601 14703 36635
rect 22066 36632 22094 36876
rect 24670 36836 24676 36848
rect 24058 36808 24676 36836
rect 24670 36796 24676 36808
rect 24728 36796 24734 36848
rect 25056 36845 25084 36876
rect 26602 36864 26608 36876
rect 26660 36864 26666 36916
rect 27080 36876 29132 36904
rect 25041 36839 25099 36845
rect 25041 36805 25053 36839
rect 25087 36805 25099 36839
rect 25041 36799 25099 36805
rect 25498 36796 25504 36848
rect 25556 36796 25562 36848
rect 22554 36700 22560 36712
rect 22515 36672 22560 36700
rect 22554 36660 22560 36672
rect 22612 36660 22618 36712
rect 22833 36703 22891 36709
rect 22833 36669 22845 36703
rect 22879 36700 22891 36703
rect 24762 36700 24768 36712
rect 22879 36672 23980 36700
rect 24723 36672 24768 36700
rect 22879 36669 22891 36672
rect 22833 36663 22891 36669
rect 23952 36644 23980 36672
rect 24762 36660 24768 36672
rect 24820 36660 24826 36712
rect 27080 36700 27108 36876
rect 28258 36796 28264 36848
rect 28316 36796 28322 36848
rect 29104 36836 29132 36876
rect 29638 36864 29644 36916
rect 29696 36904 29702 36916
rect 29696 36876 31432 36904
rect 29696 36864 29702 36876
rect 30101 36839 30159 36845
rect 30101 36836 30113 36839
rect 29104 36808 30113 36836
rect 30101 36805 30113 36808
rect 30147 36836 30159 36839
rect 30374 36836 30380 36848
rect 30147 36808 30380 36836
rect 30147 36805 30159 36808
rect 30101 36799 30159 36805
rect 30374 36796 30380 36808
rect 30432 36796 30438 36848
rect 30558 36796 30564 36848
rect 30616 36796 30622 36848
rect 31404 36768 31432 36876
rect 31662 36864 31668 36916
rect 31720 36904 31726 36916
rect 32490 36904 32496 36916
rect 31720 36876 32496 36904
rect 31720 36864 31726 36876
rect 32490 36864 32496 36876
rect 32548 36864 32554 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37645 36907 37703 36913
rect 37645 36904 37657 36907
rect 37424 36876 37657 36904
rect 37424 36864 37430 36876
rect 37645 36873 37657 36876
rect 37691 36873 37703 36907
rect 37645 36867 37703 36873
rect 32214 36796 32220 36848
rect 32272 36836 32278 36848
rect 32272 36808 33180 36836
rect 32272 36796 32278 36808
rect 33152 36777 33180 36808
rect 34054 36796 34060 36848
rect 34112 36836 34118 36848
rect 34425 36839 34483 36845
rect 34425 36836 34437 36839
rect 34112 36808 34437 36836
rect 34112 36796 34118 36808
rect 34425 36805 34437 36808
rect 34471 36805 34483 36839
rect 36538 36836 36544 36848
rect 35650 36808 36544 36836
rect 34425 36799 34483 36805
rect 36538 36796 36544 36808
rect 36596 36796 36602 36848
rect 36722 36836 36728 36848
rect 36683 36808 36728 36836
rect 36722 36796 36728 36808
rect 36780 36796 36786 36848
rect 32493 36771 32551 36777
rect 32493 36768 32505 36771
rect 31404 36740 32505 36768
rect 32493 36737 32505 36740
rect 32539 36737 32551 36771
rect 32493 36731 32551 36737
rect 33137 36771 33195 36777
rect 33137 36737 33149 36771
rect 33183 36737 33195 36771
rect 37458 36768 37464 36780
rect 37419 36740 37464 36768
rect 33137 36731 33195 36737
rect 37458 36728 37464 36740
rect 37516 36728 37522 36780
rect 24872 36672 27108 36700
rect 14645 36595 14703 36601
rect 18984 36604 22094 36632
rect 18984 36564 19012 36604
rect 23934 36592 23940 36644
rect 23992 36592 23998 36644
rect 24578 36592 24584 36644
rect 24636 36632 24642 36644
rect 24872 36632 24900 36672
rect 27154 36660 27160 36712
rect 27212 36700 27218 36712
rect 27522 36700 27528 36712
rect 27212 36672 27528 36700
rect 27212 36660 27218 36672
rect 27522 36660 27528 36672
rect 27580 36660 27586 36712
rect 27798 36700 27804 36712
rect 27632 36672 27804 36700
rect 24636 36604 24900 36632
rect 26513 36635 26571 36641
rect 24636 36592 24642 36604
rect 26513 36601 26525 36635
rect 26559 36632 26571 36635
rect 27632 36632 27660 36672
rect 27798 36660 27804 36672
rect 27856 36660 27862 36712
rect 29822 36660 29828 36712
rect 29880 36700 29886 36712
rect 34149 36703 34207 36709
rect 34149 36700 34161 36703
rect 29880 36672 29925 36700
rect 31128 36672 34161 36700
rect 29880 36660 29886 36672
rect 26559 36604 27660 36632
rect 26559 36601 26571 36604
rect 26513 36595 26571 36601
rect 28810 36592 28816 36644
rect 28868 36632 28874 36644
rect 29273 36635 29331 36641
rect 29273 36632 29285 36635
rect 28868 36604 29285 36632
rect 28868 36592 28874 36604
rect 29273 36601 29285 36604
rect 29319 36601 29331 36635
rect 29273 36595 29331 36601
rect 19426 36564 19432 36576
rect 13280 36536 19012 36564
rect 19387 36536 19432 36564
rect 19426 36524 19432 36536
rect 19484 36524 19490 36576
rect 20254 36524 20260 36576
rect 20312 36564 20318 36576
rect 24305 36567 24363 36573
rect 24305 36564 24317 36567
rect 20312 36536 24317 36564
rect 20312 36524 20318 36536
rect 24305 36533 24317 36536
rect 24351 36564 24363 36567
rect 25130 36564 25136 36576
rect 24351 36536 25136 36564
rect 24351 36533 24363 36536
rect 24305 36527 24363 36533
rect 25130 36524 25136 36536
rect 25188 36524 25194 36576
rect 25222 36524 25228 36576
rect 25280 36564 25286 36576
rect 29086 36564 29092 36576
rect 25280 36536 29092 36564
rect 25280 36524 25286 36536
rect 29086 36524 29092 36536
rect 29144 36524 29150 36576
rect 29822 36524 29828 36576
rect 29880 36564 29886 36576
rect 31128 36564 31156 36672
rect 33152 36644 33180 36672
rect 34149 36669 34161 36672
rect 34195 36669 34207 36703
rect 34149 36663 34207 36669
rect 33134 36592 33140 36644
rect 33192 36592 33198 36644
rect 29880 36536 31156 36564
rect 29880 36524 29886 36536
rect 31294 36524 31300 36576
rect 31352 36564 31358 36576
rect 31573 36567 31631 36573
rect 31573 36564 31585 36567
rect 31352 36536 31585 36564
rect 31352 36524 31358 36536
rect 31573 36533 31585 36536
rect 31619 36533 31631 36567
rect 32306 36564 32312 36576
rect 32267 36536 32312 36564
rect 31573 36527 31631 36533
rect 32306 36524 32312 36536
rect 32364 36524 32370 36576
rect 32398 36524 32404 36576
rect 32456 36564 32462 36576
rect 32953 36567 33011 36573
rect 32953 36564 32965 36567
rect 32456 36536 32965 36564
rect 32456 36524 32462 36536
rect 32953 36533 32965 36536
rect 32999 36533 33011 36567
rect 32953 36527 33011 36533
rect 35894 36524 35900 36576
rect 35952 36564 35958 36576
rect 35952 36536 35997 36564
rect 35952 36524 35958 36536
rect 36078 36524 36084 36576
rect 36136 36564 36142 36576
rect 36817 36567 36875 36573
rect 36817 36564 36829 36567
rect 36136 36536 36829 36564
rect 36136 36524 36142 36536
rect 36817 36533 36829 36536
rect 36863 36533 36875 36567
rect 36817 36527 36875 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 8478 36360 8484 36372
rect 8439 36332 8484 36360
rect 8478 36320 8484 36332
rect 8536 36320 8542 36372
rect 8662 36320 8668 36372
rect 8720 36360 8726 36372
rect 9858 36360 9864 36372
rect 8720 36332 9864 36360
rect 8720 36320 8726 36332
rect 9858 36320 9864 36332
rect 9916 36360 9922 36372
rect 10594 36360 10600 36372
rect 9916 36332 10600 36360
rect 9916 36320 9922 36332
rect 10594 36320 10600 36332
rect 10652 36320 10658 36372
rect 11882 36360 11888 36372
rect 11532 36332 11888 36360
rect 7837 36295 7895 36301
rect 7837 36261 7849 36295
rect 7883 36292 7895 36295
rect 11532 36292 11560 36332
rect 11882 36320 11888 36332
rect 11940 36320 11946 36372
rect 11974 36320 11980 36372
rect 12032 36360 12038 36372
rect 12032 36332 17264 36360
rect 12032 36320 12038 36332
rect 17236 36292 17264 36332
rect 17954 36320 17960 36372
rect 18012 36360 18018 36372
rect 18012 36332 22094 36360
rect 18012 36320 18018 36332
rect 20622 36292 20628 36304
rect 7883 36264 11560 36292
rect 11624 36264 15884 36292
rect 17236 36264 20628 36292
rect 7883 36261 7895 36264
rect 7837 36255 7895 36261
rect 1578 36224 1584 36236
rect 1539 36196 1584 36224
rect 1578 36184 1584 36196
rect 1636 36184 1642 36236
rect 11514 36224 11520 36236
rect 8404 36196 11520 36224
rect 4157 36159 4215 36165
rect 4157 36125 4169 36159
rect 4203 36156 4215 36159
rect 4614 36156 4620 36168
rect 4203 36128 4620 36156
rect 4203 36125 4215 36128
rect 4157 36119 4215 36125
rect 4614 36116 4620 36128
rect 4672 36116 4678 36168
rect 6730 36156 6736 36168
rect 6691 36128 6736 36156
rect 6730 36116 6736 36128
rect 6788 36116 6794 36168
rect 8404 36165 8432 36196
rect 11514 36184 11520 36196
rect 11572 36184 11578 36236
rect 7745 36159 7803 36165
rect 7745 36125 7757 36159
rect 7791 36125 7803 36159
rect 7745 36119 7803 36125
rect 8389 36159 8447 36165
rect 8389 36125 8401 36159
rect 8435 36125 8447 36159
rect 9582 36156 9588 36168
rect 9543 36128 9588 36156
rect 8389 36119 8447 36125
rect 1762 36088 1768 36100
rect 1723 36060 1768 36088
rect 1762 36048 1768 36060
rect 1820 36048 1826 36100
rect 3421 36091 3479 36097
rect 3421 36057 3433 36091
rect 3467 36088 3479 36091
rect 5442 36088 5448 36100
rect 3467 36060 5448 36088
rect 3467 36057 3479 36060
rect 3421 36051 3479 36057
rect 5442 36048 5448 36060
rect 5500 36048 5506 36100
rect 7760 36088 7788 36119
rect 9582 36116 9588 36128
rect 9640 36116 9646 36168
rect 10321 36159 10379 36165
rect 10321 36125 10333 36159
rect 10367 36156 10379 36159
rect 10594 36156 10600 36168
rect 10367 36128 10600 36156
rect 10367 36125 10379 36128
rect 10321 36119 10379 36125
rect 10594 36116 10600 36128
rect 10652 36116 10658 36168
rect 10686 36116 10692 36168
rect 10744 36156 10750 36168
rect 11624 36165 11652 36264
rect 12897 36227 12955 36233
rect 12897 36193 12909 36227
rect 12943 36224 12955 36227
rect 13170 36224 13176 36236
rect 12943 36196 13176 36224
rect 12943 36193 12955 36196
rect 12897 36187 12955 36193
rect 13170 36184 13176 36196
rect 13228 36184 13234 36236
rect 13814 36184 13820 36236
rect 13872 36224 13878 36236
rect 14737 36227 14795 36233
rect 14737 36224 14749 36227
rect 13872 36196 14749 36224
rect 13872 36184 13878 36196
rect 14737 36193 14749 36196
rect 14783 36193 14795 36227
rect 14737 36187 14795 36193
rect 10965 36159 11023 36165
rect 10965 36156 10977 36159
rect 10744 36128 10977 36156
rect 10744 36116 10750 36128
rect 10965 36125 10977 36128
rect 11011 36125 11023 36159
rect 10965 36119 11023 36125
rect 11609 36159 11667 36165
rect 11609 36125 11621 36159
rect 11655 36125 11667 36159
rect 12986 36156 12992 36168
rect 11609 36119 11667 36125
rect 11716 36128 12992 36156
rect 11716 36088 11744 36128
rect 12986 36116 12992 36128
rect 13044 36116 13050 36168
rect 13078 36116 13084 36168
rect 13136 36156 13142 36168
rect 13136 36128 13181 36156
rect 13136 36116 13142 36128
rect 7760 36060 11744 36088
rect 11882 36048 11888 36100
rect 11940 36088 11946 36100
rect 14458 36088 14464 36100
rect 11940 36060 13676 36088
rect 14419 36060 14464 36088
rect 11940 36048 11946 36060
rect 3973 36023 4031 36029
rect 3973 35989 3985 36023
rect 4019 36020 4031 36023
rect 6730 36020 6736 36032
rect 4019 35992 6736 36020
rect 4019 35989 4031 35992
rect 3973 35983 4031 35989
rect 6730 35980 6736 35992
rect 6788 35980 6794 36032
rect 6825 36023 6883 36029
rect 6825 35989 6837 36023
rect 6871 36020 6883 36023
rect 8018 36020 8024 36032
rect 6871 35992 8024 36020
rect 6871 35989 6883 35992
rect 6825 35983 6883 35989
rect 8018 35980 8024 35992
rect 8076 35980 8082 36032
rect 9030 35980 9036 36032
rect 9088 36020 9094 36032
rect 9398 36020 9404 36032
rect 9088 35992 9404 36020
rect 9088 35980 9094 35992
rect 9398 35980 9404 35992
rect 9456 35980 9462 36032
rect 9674 36020 9680 36032
rect 9635 35992 9680 36020
rect 9674 35980 9680 35992
rect 9732 35980 9738 36032
rect 10410 36020 10416 36032
rect 10371 35992 10416 36020
rect 10410 35980 10416 35992
rect 10468 35980 10474 36032
rect 11054 36020 11060 36032
rect 11015 35992 11060 36020
rect 11054 35980 11060 35992
rect 11112 35980 11118 36032
rect 11701 36023 11759 36029
rect 11701 35989 11713 36023
rect 11747 36020 11759 36023
rect 12066 36020 12072 36032
rect 11747 35992 12072 36020
rect 11747 35989 11759 35992
rect 11701 35983 11759 35989
rect 12066 35980 12072 35992
rect 12124 35980 12130 36032
rect 13538 36020 13544 36032
rect 13499 35992 13544 36020
rect 13538 35980 13544 35992
rect 13596 35980 13602 36032
rect 13648 36020 13676 36060
rect 14458 36048 14464 36060
rect 14516 36048 14522 36100
rect 14553 36091 14611 36097
rect 14553 36057 14565 36091
rect 14599 36057 14611 36091
rect 14553 36051 14611 36057
rect 14568 36020 14596 36051
rect 13648 35992 14596 36020
rect 15856 36020 15884 36264
rect 20622 36252 20628 36264
rect 20680 36252 20686 36304
rect 22066 36292 22094 36332
rect 23474 36320 23480 36372
rect 23532 36360 23538 36372
rect 26602 36360 26608 36372
rect 23532 36332 26188 36360
rect 26563 36332 26608 36360
rect 23532 36320 23538 36332
rect 24578 36292 24584 36304
rect 22066 36264 24584 36292
rect 24578 36252 24584 36264
rect 24636 36252 24642 36304
rect 26160 36292 26188 36332
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 27062 36320 27068 36372
rect 27120 36360 27126 36372
rect 32398 36360 32404 36372
rect 27120 36332 32404 36360
rect 27120 36320 27126 36332
rect 32398 36320 32404 36332
rect 32456 36320 32462 36372
rect 32490 36320 32496 36372
rect 32548 36360 32554 36372
rect 35894 36360 35900 36372
rect 32548 36332 35900 36360
rect 32548 36320 32554 36332
rect 35894 36320 35900 36332
rect 35952 36320 35958 36372
rect 36170 36320 36176 36372
rect 36228 36360 36234 36372
rect 37369 36363 37427 36369
rect 37369 36360 37381 36363
rect 36228 36332 37381 36360
rect 36228 36320 36234 36332
rect 37369 36329 37381 36332
rect 37415 36329 37427 36363
rect 37369 36323 37427 36329
rect 29733 36295 29791 36301
rect 26160 36264 29316 36292
rect 15933 36227 15991 36233
rect 15933 36193 15945 36227
rect 15979 36224 15991 36227
rect 16850 36224 16856 36236
rect 15979 36196 16856 36224
rect 15979 36193 15991 36196
rect 15933 36187 15991 36193
rect 16850 36184 16856 36196
rect 16908 36184 16914 36236
rect 16942 36184 16948 36236
rect 17000 36224 17006 36236
rect 20530 36224 20536 36236
rect 17000 36196 20536 36224
rect 17000 36184 17006 36196
rect 20530 36184 20536 36196
rect 20588 36184 20594 36236
rect 20717 36227 20775 36233
rect 20717 36193 20729 36227
rect 20763 36224 20775 36227
rect 22278 36224 22284 36236
rect 20763 36196 22284 36224
rect 20763 36193 20775 36196
rect 20717 36187 20775 36193
rect 22278 36184 22284 36196
rect 22336 36224 22342 36236
rect 22554 36224 22560 36236
rect 22336 36196 22560 36224
rect 22336 36184 22342 36196
rect 22554 36184 22560 36196
rect 22612 36224 22618 36236
rect 23753 36227 23811 36233
rect 23753 36224 23765 36227
rect 22612 36196 23765 36224
rect 22612 36184 22618 36196
rect 23753 36193 23765 36196
rect 23799 36224 23811 36227
rect 24762 36224 24768 36236
rect 23799 36196 24768 36224
rect 23799 36193 23811 36196
rect 23753 36187 23811 36193
rect 24762 36184 24768 36196
rect 24820 36224 24826 36236
rect 24857 36227 24915 36233
rect 24857 36224 24869 36227
rect 24820 36196 24869 36224
rect 24820 36184 24826 36196
rect 24857 36193 24869 36196
rect 24903 36193 24915 36227
rect 25130 36224 25136 36236
rect 25091 36196 25136 36224
rect 24857 36187 24915 36193
rect 25130 36184 25136 36196
rect 25188 36184 25194 36236
rect 27801 36227 27859 36233
rect 27801 36193 27813 36227
rect 27847 36224 27859 36227
rect 27982 36224 27988 36236
rect 27847 36196 27988 36224
rect 27847 36193 27859 36196
rect 27801 36187 27859 36193
rect 27982 36184 27988 36196
rect 28040 36184 28046 36236
rect 28442 36184 28448 36236
rect 28500 36224 28506 36236
rect 29086 36224 29092 36236
rect 28500 36196 29092 36224
rect 28500 36184 28506 36196
rect 29086 36184 29092 36196
rect 29144 36184 29150 36236
rect 28345 36169 28403 36175
rect 17862 36116 17868 36168
rect 17920 36156 17926 36168
rect 19426 36156 19432 36168
rect 17920 36128 19432 36156
rect 17920 36116 17926 36128
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 22094 36116 22100 36168
rect 22152 36116 22158 36168
rect 26234 36116 26240 36168
rect 26292 36116 26298 36168
rect 27062 36156 27068 36168
rect 27023 36128 27068 36156
rect 27062 36116 27068 36128
rect 27120 36116 27126 36168
rect 27706 36156 27712 36168
rect 27667 36128 27712 36156
rect 27706 36116 27712 36128
rect 27764 36116 27770 36168
rect 28166 36116 28172 36168
rect 28224 36166 28230 36168
rect 28345 36166 28357 36169
rect 28224 36138 28357 36166
rect 28224 36116 28230 36138
rect 28345 36135 28357 36138
rect 28391 36135 28403 36169
rect 28345 36129 28403 36135
rect 28994 36116 29000 36168
rect 29052 36156 29058 36168
rect 29181 36159 29239 36165
rect 29181 36156 29193 36159
rect 29052 36128 29193 36156
rect 29052 36116 29058 36128
rect 29181 36125 29193 36128
rect 29227 36125 29239 36159
rect 29288 36156 29316 36264
rect 29733 36261 29745 36295
rect 29779 36261 29791 36295
rect 29733 36255 29791 36261
rect 36081 36295 36139 36301
rect 36081 36261 36093 36295
rect 36127 36292 36139 36295
rect 36262 36292 36268 36304
rect 36127 36264 36268 36292
rect 36127 36261 36139 36264
rect 36081 36255 36139 36261
rect 29748 36224 29776 36255
rect 36262 36252 36268 36264
rect 36320 36252 36326 36304
rect 33686 36224 33692 36236
rect 29748 36196 33692 36224
rect 33686 36184 33692 36196
rect 33744 36184 33750 36236
rect 29917 36159 29975 36165
rect 29917 36156 29929 36159
rect 29288 36128 29929 36156
rect 29181 36119 29239 36125
rect 29917 36125 29929 36128
rect 29963 36125 29975 36159
rect 29917 36119 29975 36125
rect 30466 36116 30472 36168
rect 30524 36156 30530 36168
rect 30929 36159 30987 36165
rect 30929 36156 30941 36159
rect 30524 36128 30941 36156
rect 30524 36116 30530 36128
rect 30929 36125 30941 36128
rect 30975 36125 30987 36159
rect 30929 36119 30987 36125
rect 33502 36116 33508 36168
rect 33560 36156 33566 36168
rect 34885 36159 34943 36165
rect 34885 36156 34897 36159
rect 33560 36128 34897 36156
rect 33560 36116 33566 36128
rect 34885 36125 34897 36128
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 35897 36159 35955 36165
rect 35897 36125 35909 36159
rect 35943 36125 35955 36159
rect 35897 36119 35955 36125
rect 16206 36088 16212 36100
rect 16167 36060 16212 36088
rect 16206 36048 16212 36060
rect 16264 36048 16270 36100
rect 16666 36048 16672 36100
rect 16724 36048 16730 36100
rect 17770 36048 17776 36100
rect 17828 36088 17834 36100
rect 17957 36091 18015 36097
rect 17957 36088 17969 36091
rect 17828 36060 17969 36088
rect 17828 36048 17834 36060
rect 17957 36057 17969 36060
rect 18003 36057 18015 36091
rect 20990 36088 20996 36100
rect 20951 36060 20996 36088
rect 17957 36051 18015 36057
rect 20990 36048 20996 36060
rect 21048 36048 21054 36100
rect 22925 36091 22983 36097
rect 22925 36057 22937 36091
rect 22971 36088 22983 36091
rect 23106 36088 23112 36100
rect 22971 36060 23112 36088
rect 22971 36057 22983 36060
rect 22925 36051 22983 36057
rect 23106 36048 23112 36060
rect 23164 36048 23170 36100
rect 24578 36048 24584 36100
rect 24636 36088 24642 36100
rect 24636 36060 25360 36088
rect 24636 36048 24642 36060
rect 22465 36023 22523 36029
rect 22465 36020 22477 36023
rect 15856 35992 22477 36020
rect 22465 35989 22477 35992
rect 22511 36020 22523 36023
rect 25222 36020 25228 36032
rect 22511 35992 25228 36020
rect 22511 35989 22523 35992
rect 22465 35983 22523 35989
rect 25222 35980 25228 35992
rect 25280 35980 25286 36032
rect 25332 36020 25360 36060
rect 26418 36048 26424 36100
rect 26476 36088 26482 36100
rect 27157 36091 27215 36097
rect 27157 36088 27169 36091
rect 26476 36060 27169 36088
rect 26476 36048 26482 36060
rect 27157 36057 27169 36060
rect 27203 36057 27215 36091
rect 27157 36051 27215 36057
rect 31110 36048 31116 36100
rect 31168 36088 31174 36100
rect 31205 36091 31263 36097
rect 31205 36088 31217 36091
rect 31168 36060 31217 36088
rect 31168 36048 31174 36060
rect 31205 36057 31217 36060
rect 31251 36057 31263 36091
rect 35250 36088 35256 36100
rect 32430 36060 35256 36088
rect 31205 36051 31263 36057
rect 35250 36048 35256 36060
rect 35308 36048 35314 36100
rect 35912 36088 35940 36119
rect 36170 36116 36176 36168
rect 36228 36156 36234 36168
rect 36633 36159 36691 36165
rect 36633 36156 36645 36159
rect 36228 36128 36645 36156
rect 36228 36116 36234 36128
rect 36633 36125 36645 36128
rect 36679 36125 36691 36159
rect 36633 36119 36691 36125
rect 36909 36159 36967 36165
rect 36909 36125 36921 36159
rect 36955 36156 36967 36159
rect 37553 36159 37611 36165
rect 37553 36156 37565 36159
rect 36955 36128 37565 36156
rect 36955 36125 36967 36128
rect 36909 36119 36967 36125
rect 37553 36125 37565 36128
rect 37599 36125 37611 36159
rect 37553 36119 37611 36125
rect 37826 36116 37832 36168
rect 37884 36156 37890 36168
rect 38013 36159 38071 36165
rect 38013 36156 38025 36159
rect 37884 36128 38025 36156
rect 37884 36116 37890 36128
rect 38013 36125 38025 36128
rect 38059 36125 38071 36159
rect 38013 36119 38071 36125
rect 37734 36088 37740 36100
rect 35912 36060 37740 36088
rect 37734 36048 37740 36060
rect 37792 36048 37798 36100
rect 28350 36020 28356 36032
rect 25332 35992 28356 36020
rect 28350 35980 28356 35992
rect 28408 35980 28414 36032
rect 28442 35980 28448 36032
rect 28500 36020 28506 36032
rect 28500 35992 28545 36020
rect 28500 35980 28506 35992
rect 28626 35980 28632 36032
rect 28684 36020 28690 36032
rect 28997 36023 29055 36029
rect 28997 36020 29009 36023
rect 28684 35992 29009 36020
rect 28684 35980 28690 35992
rect 28997 35989 29009 35992
rect 29043 35989 29055 36023
rect 28997 35983 29055 35989
rect 29178 35980 29184 36032
rect 29236 36020 29242 36032
rect 31294 36020 31300 36032
rect 29236 35992 31300 36020
rect 29236 35980 29242 35992
rect 31294 35980 31300 35992
rect 31352 35980 31358 36032
rect 32582 35980 32588 36032
rect 32640 36020 32646 36032
rect 32677 36023 32735 36029
rect 32677 36020 32689 36023
rect 32640 35992 32689 36020
rect 32640 35980 32646 35992
rect 32677 35989 32689 35992
rect 32723 35989 32735 36023
rect 32677 35983 32735 35989
rect 34977 36023 35035 36029
rect 34977 35989 34989 36023
rect 35023 36020 35035 36023
rect 35526 36020 35532 36032
rect 35023 35992 35532 36020
rect 35023 35989 35035 35992
rect 34977 35983 35035 35989
rect 35526 35980 35532 35992
rect 35584 35980 35590 36032
rect 38194 36020 38200 36032
rect 38155 35992 38200 36020
rect 38194 35980 38200 35992
rect 38252 35980 38258 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1762 35776 1768 35828
rect 1820 35816 1826 35828
rect 2409 35819 2467 35825
rect 2409 35816 2421 35819
rect 1820 35788 2421 35816
rect 1820 35776 1826 35788
rect 2409 35785 2421 35788
rect 2455 35785 2467 35819
rect 2409 35779 2467 35785
rect 8294 35776 8300 35828
rect 8352 35816 8358 35828
rect 10778 35816 10784 35828
rect 8352 35788 10784 35816
rect 8352 35776 8358 35788
rect 10778 35776 10784 35788
rect 10836 35776 10842 35828
rect 12342 35776 12348 35828
rect 12400 35816 12406 35828
rect 13078 35816 13084 35828
rect 12400 35788 13084 35816
rect 12400 35776 12406 35788
rect 13078 35776 13084 35788
rect 13136 35776 13142 35828
rect 14458 35816 14464 35828
rect 14419 35788 14464 35816
rect 14458 35776 14464 35788
rect 14516 35776 14522 35828
rect 29270 35816 29276 35828
rect 16316 35788 29276 35816
rect 3050 35748 3056 35760
rect 3011 35720 3056 35748
rect 3050 35708 3056 35720
rect 3108 35708 3114 35760
rect 3145 35751 3203 35757
rect 3145 35717 3157 35751
rect 3191 35748 3203 35751
rect 3970 35748 3976 35760
rect 3191 35720 3976 35748
rect 3191 35717 3203 35720
rect 3145 35711 3203 35717
rect 3970 35708 3976 35720
rect 4028 35708 4034 35760
rect 6641 35751 6699 35757
rect 6641 35717 6653 35751
rect 6687 35748 6699 35751
rect 9398 35748 9404 35760
rect 6687 35720 9404 35748
rect 6687 35717 6699 35720
rect 6641 35711 6699 35717
rect 9398 35708 9404 35720
rect 9456 35708 9462 35760
rect 11514 35748 11520 35760
rect 9692 35720 11520 35748
rect 1486 35640 1492 35692
rect 1544 35680 1550 35692
rect 1581 35683 1639 35689
rect 1581 35680 1593 35683
rect 1544 35652 1593 35680
rect 1544 35640 1550 35652
rect 1581 35649 1593 35652
rect 1627 35649 1639 35683
rect 2314 35680 2320 35692
rect 2275 35652 2320 35680
rect 1581 35643 1639 35649
rect 2314 35640 2320 35652
rect 2372 35640 2378 35692
rect 6546 35680 6552 35692
rect 6507 35652 6552 35680
rect 6546 35640 6552 35652
rect 6604 35640 6610 35692
rect 8297 35683 8355 35689
rect 8297 35649 8309 35683
rect 8343 35680 8355 35683
rect 8570 35680 8576 35692
rect 8343 35652 8576 35680
rect 8343 35649 8355 35652
rect 8297 35643 8355 35649
rect 8570 35640 8576 35652
rect 8628 35640 8634 35692
rect 9692 35680 9720 35720
rect 11514 35708 11520 35720
rect 11572 35708 11578 35760
rect 11882 35708 11888 35760
rect 11940 35757 11946 35760
rect 11940 35748 11952 35757
rect 11940 35720 11985 35748
rect 11940 35711 11952 35720
rect 11940 35708 11946 35711
rect 12066 35708 12072 35760
rect 12124 35748 12130 35760
rect 16316 35757 16344 35788
rect 29270 35776 29276 35788
rect 29328 35776 29334 35828
rect 30193 35819 30251 35825
rect 30193 35785 30205 35819
rect 30239 35816 30251 35819
rect 31570 35816 31576 35828
rect 30239 35788 31576 35816
rect 30239 35785 30251 35788
rect 30193 35779 30251 35785
rect 31570 35776 31576 35788
rect 31628 35776 31634 35828
rect 15381 35751 15439 35757
rect 15381 35748 15393 35751
rect 12124 35720 15393 35748
rect 12124 35708 12130 35720
rect 15381 35717 15393 35720
rect 15427 35717 15439 35751
rect 15381 35711 15439 35717
rect 16301 35751 16359 35757
rect 16301 35717 16313 35751
rect 16347 35717 16359 35751
rect 16301 35711 16359 35717
rect 17586 35708 17592 35760
rect 17644 35708 17650 35760
rect 18414 35708 18420 35760
rect 18472 35748 18478 35760
rect 19702 35748 19708 35760
rect 18472 35720 19708 35748
rect 18472 35708 18478 35720
rect 19702 35708 19708 35720
rect 19760 35708 19766 35760
rect 20070 35708 20076 35760
rect 20128 35708 20134 35760
rect 23290 35708 23296 35760
rect 23348 35708 23354 35760
rect 33502 35748 33508 35760
rect 33463 35720 33508 35748
rect 33502 35708 33508 35720
rect 33560 35708 33566 35760
rect 35618 35748 35624 35760
rect 34730 35720 35624 35748
rect 35618 35708 35624 35720
rect 35676 35708 35682 35760
rect 8680 35652 9720 35680
rect 10597 35683 10655 35689
rect 8680 35624 8708 35652
rect 10597 35649 10609 35683
rect 10643 35680 10655 35683
rect 10686 35680 10692 35692
rect 10643 35652 10692 35680
rect 10643 35649 10655 35652
rect 10597 35643 10655 35649
rect 10686 35640 10692 35652
rect 10744 35640 10750 35692
rect 11330 35640 11336 35692
rect 11388 35680 11394 35692
rect 11388 35652 11652 35680
rect 11388 35640 11394 35652
rect 3697 35615 3755 35621
rect 3697 35581 3709 35615
rect 3743 35612 3755 35615
rect 8662 35612 8668 35624
rect 3743 35584 8668 35612
rect 3743 35581 3755 35584
rect 3697 35575 3755 35581
rect 8662 35572 8668 35584
rect 8720 35572 8726 35624
rect 9398 35572 9404 35624
rect 9456 35612 9462 35624
rect 9493 35615 9551 35621
rect 9493 35612 9505 35615
rect 9456 35584 9505 35612
rect 9456 35572 9462 35584
rect 9493 35581 9505 35584
rect 9539 35581 9551 35615
rect 9493 35575 9551 35581
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 10318 35612 10324 35624
rect 9723 35584 10324 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 10318 35572 10324 35584
rect 10376 35572 10382 35624
rect 11624 35612 11652 35652
rect 12710 35640 12716 35692
rect 12768 35680 12774 35692
rect 16850 35680 16856 35692
rect 12768 35652 13400 35680
rect 16811 35652 16856 35680
rect 12768 35640 12774 35652
rect 11793 35615 11851 35621
rect 11793 35612 11805 35615
rect 11624 35584 11805 35612
rect 11793 35581 11805 35584
rect 11839 35581 11851 35615
rect 11793 35575 11851 35581
rect 12618 35572 12624 35624
rect 12676 35612 12682 35624
rect 12805 35615 12863 35621
rect 12805 35612 12817 35615
rect 12676 35584 12817 35612
rect 12676 35572 12682 35584
rect 12805 35581 12817 35584
rect 12851 35612 12863 35615
rect 12894 35612 12900 35624
rect 12851 35584 12900 35612
rect 12851 35581 12863 35584
rect 12805 35575 12863 35581
rect 12894 35572 12900 35584
rect 12952 35572 12958 35624
rect 13078 35572 13084 35624
rect 13136 35612 13142 35624
rect 13265 35615 13323 35621
rect 13265 35612 13277 35615
rect 13136 35584 13277 35612
rect 13136 35572 13142 35584
rect 13265 35581 13277 35584
rect 13311 35581 13323 35615
rect 13372 35612 13400 35652
rect 16850 35640 16856 35652
rect 16908 35640 16914 35692
rect 22278 35680 22284 35692
rect 22239 35652 22284 35680
rect 22278 35640 22284 35652
rect 22336 35640 22342 35692
rect 30377 35683 30435 35689
rect 30377 35649 30389 35683
rect 30423 35680 30435 35683
rect 31478 35680 31484 35692
rect 30423 35652 31484 35680
rect 30423 35649 30435 35652
rect 30377 35643 30435 35649
rect 31478 35640 31484 35652
rect 31536 35640 31542 35692
rect 34790 35640 34796 35692
rect 34848 35680 34854 35692
rect 36265 35683 36323 35689
rect 36265 35680 36277 35683
rect 34848 35652 36277 35680
rect 34848 35640 34854 35652
rect 36265 35649 36277 35652
rect 36311 35649 36323 35683
rect 36265 35643 36323 35649
rect 38013 35683 38071 35689
rect 38013 35649 38025 35683
rect 38059 35680 38071 35683
rect 38378 35680 38384 35692
rect 38059 35652 38384 35680
rect 38059 35649 38071 35652
rect 38013 35643 38071 35649
rect 38378 35640 38384 35652
rect 38436 35640 38442 35692
rect 15289 35615 15347 35621
rect 15289 35612 15301 35615
rect 13372 35584 15301 35612
rect 13265 35575 13323 35581
rect 15289 35581 15301 35584
rect 15335 35581 15347 35615
rect 17126 35612 17132 35624
rect 17087 35584 17132 35612
rect 15289 35575 15347 35581
rect 17126 35572 17132 35584
rect 17184 35572 17190 35624
rect 17494 35572 17500 35624
rect 17552 35612 17558 35624
rect 19334 35612 19340 35624
rect 17552 35584 18828 35612
rect 19295 35584 19340 35612
rect 17552 35572 17558 35584
rect 1765 35547 1823 35553
rect 1765 35513 1777 35547
rect 1811 35544 1823 35547
rect 2866 35544 2872 35556
rect 1811 35516 2872 35544
rect 1811 35513 1823 35516
rect 1765 35507 1823 35513
rect 2866 35504 2872 35516
rect 2924 35504 2930 35556
rect 8570 35504 8576 35556
rect 8628 35544 8634 35556
rect 10689 35547 10747 35553
rect 8628 35516 10364 35544
rect 8628 35504 8634 35516
rect 8389 35479 8447 35485
rect 8389 35445 8401 35479
rect 8435 35476 8447 35479
rect 10042 35476 10048 35488
rect 8435 35448 10048 35476
rect 8435 35445 8447 35448
rect 8389 35439 8447 35445
rect 10042 35436 10048 35448
rect 10100 35436 10106 35488
rect 10134 35436 10140 35488
rect 10192 35476 10198 35488
rect 10336 35476 10364 35516
rect 10689 35513 10701 35547
rect 10735 35544 10747 35547
rect 16666 35544 16672 35556
rect 10735 35516 16672 35544
rect 10735 35513 10747 35516
rect 10689 35507 10747 35513
rect 16666 35504 16672 35516
rect 16724 35504 16730 35556
rect 16390 35476 16396 35488
rect 10192 35448 10237 35476
rect 10336 35448 16396 35476
rect 10192 35436 10198 35448
rect 16390 35436 16396 35448
rect 16448 35436 16454 35488
rect 17218 35436 17224 35488
rect 17276 35476 17282 35488
rect 18601 35479 18659 35485
rect 18601 35476 18613 35479
rect 17276 35448 18613 35476
rect 17276 35436 17282 35448
rect 18601 35445 18613 35448
rect 18647 35445 18659 35479
rect 18800 35476 18828 35584
rect 19334 35572 19340 35584
rect 19392 35572 19398 35624
rect 19610 35612 19616 35624
rect 19571 35584 19616 35612
rect 19610 35572 19616 35584
rect 19668 35572 19674 35624
rect 19702 35572 19708 35624
rect 19760 35612 19766 35624
rect 21085 35615 21143 35621
rect 21085 35612 21097 35615
rect 19760 35584 21097 35612
rect 19760 35572 19766 35584
rect 21085 35581 21097 35584
rect 21131 35581 21143 35615
rect 21085 35575 21143 35581
rect 22557 35615 22615 35621
rect 22557 35581 22569 35615
rect 22603 35612 22615 35615
rect 23566 35612 23572 35624
rect 22603 35584 23572 35612
rect 22603 35581 22615 35584
rect 22557 35575 22615 35581
rect 23566 35572 23572 35584
rect 23624 35572 23630 35624
rect 27157 35615 27215 35621
rect 27157 35581 27169 35615
rect 27203 35581 27215 35615
rect 27338 35612 27344 35624
rect 27299 35584 27344 35612
rect 27157 35575 27215 35581
rect 27172 35544 27200 35575
rect 27338 35572 27344 35584
rect 27396 35572 27402 35624
rect 27617 35615 27675 35621
rect 27617 35612 27629 35615
rect 27540 35584 27629 35612
rect 27430 35544 27436 35556
rect 20640 35516 22094 35544
rect 20640 35476 20668 35516
rect 18800 35448 20668 35476
rect 22066 35476 22094 35516
rect 23860 35516 27108 35544
rect 27172 35516 27436 35544
rect 23860 35476 23888 35516
rect 22066 35448 23888 35476
rect 18601 35439 18659 35445
rect 23934 35436 23940 35488
rect 23992 35476 23998 35488
rect 24029 35479 24087 35485
rect 24029 35476 24041 35479
rect 23992 35448 24041 35476
rect 23992 35436 23998 35448
rect 24029 35445 24041 35448
rect 24075 35445 24087 35479
rect 27080 35476 27108 35516
rect 27430 35504 27436 35516
rect 27488 35504 27494 35556
rect 27540 35476 27568 35584
rect 27617 35581 27629 35584
rect 27663 35581 27675 35615
rect 33226 35612 33232 35624
rect 33187 35584 33232 35612
rect 27617 35575 27675 35581
rect 33226 35572 33232 35584
rect 33284 35572 33290 35624
rect 35621 35615 35679 35621
rect 35621 35581 35633 35615
rect 35667 35612 35679 35615
rect 35710 35612 35716 35624
rect 35667 35584 35716 35612
rect 35667 35581 35679 35584
rect 35621 35575 35679 35581
rect 35710 35572 35716 35584
rect 35768 35572 35774 35624
rect 28718 35476 28724 35488
rect 27080 35448 28724 35476
rect 24029 35439 24087 35445
rect 28718 35436 28724 35448
rect 28776 35436 28782 35488
rect 34698 35436 34704 35488
rect 34756 35476 34762 35488
rect 34977 35479 35035 35485
rect 34977 35476 34989 35479
rect 34756 35448 34989 35476
rect 34756 35436 34762 35448
rect 34977 35445 34989 35448
rect 35023 35445 35035 35479
rect 34977 35439 35035 35445
rect 36357 35479 36415 35485
rect 36357 35445 36369 35479
rect 36403 35476 36415 35479
rect 37550 35476 37556 35488
rect 36403 35448 37556 35476
rect 36403 35445 36415 35448
rect 36357 35439 36415 35445
rect 37550 35436 37556 35448
rect 37608 35436 37614 35488
rect 38194 35476 38200 35488
rect 38155 35448 38200 35476
rect 38194 35436 38200 35448
rect 38252 35436 38258 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1581 35275 1639 35281
rect 1581 35241 1593 35275
rect 1627 35272 1639 35275
rect 6546 35272 6552 35284
rect 1627 35244 6552 35272
rect 1627 35241 1639 35244
rect 1581 35235 1639 35241
rect 6546 35232 6552 35244
rect 6604 35232 6610 35284
rect 15378 35272 15384 35284
rect 8404 35244 15384 35272
rect 2225 35207 2283 35213
rect 2225 35173 2237 35207
rect 2271 35204 2283 35207
rect 6914 35204 6920 35216
rect 2271 35176 6920 35204
rect 2271 35173 2283 35176
rect 2225 35167 2283 35173
rect 6914 35164 6920 35176
rect 6972 35164 6978 35216
rect 658 35096 664 35148
rect 716 35136 722 35148
rect 716 35108 2452 35136
rect 716 35096 722 35108
rect 1394 35028 1400 35080
rect 1452 35068 1458 35080
rect 2424 35077 2452 35108
rect 1765 35071 1823 35077
rect 1765 35068 1777 35071
rect 1452 35040 1777 35068
rect 1452 35028 1458 35040
rect 1765 35037 1777 35040
rect 1811 35037 1823 35071
rect 1765 35031 1823 35037
rect 2409 35071 2467 35077
rect 2409 35037 2421 35071
rect 2455 35037 2467 35071
rect 2409 35031 2467 35037
rect 4341 35071 4399 35077
rect 4341 35037 4353 35071
rect 4387 35037 4399 35071
rect 6454 35068 6460 35080
rect 6415 35040 6460 35068
rect 4341 35031 4399 35037
rect 4356 35000 4384 35031
rect 6454 35028 6460 35040
rect 6512 35028 6518 35080
rect 8404 35077 8432 35244
rect 15378 35232 15384 35244
rect 15436 35232 15442 35284
rect 15562 35232 15568 35284
rect 15620 35272 15626 35284
rect 19610 35272 19616 35284
rect 15620 35244 19616 35272
rect 15620 35232 15626 35244
rect 19610 35232 19616 35244
rect 19668 35272 19674 35284
rect 21818 35272 21824 35284
rect 19668 35244 21824 35272
rect 19668 35232 19674 35244
rect 21818 35232 21824 35244
rect 21876 35232 21882 35284
rect 22186 35232 22192 35284
rect 22244 35272 22250 35284
rect 32306 35272 32312 35284
rect 22244 35244 32312 35272
rect 22244 35232 22250 35244
rect 32306 35232 32312 35244
rect 32364 35232 32370 35284
rect 35250 35232 35256 35284
rect 35308 35272 35314 35284
rect 35710 35272 35716 35284
rect 35308 35244 35716 35272
rect 35308 35232 35314 35244
rect 35710 35232 35716 35244
rect 35768 35232 35774 35284
rect 38197 35275 38255 35281
rect 38197 35241 38209 35275
rect 38243 35272 38255 35275
rect 39298 35272 39304 35284
rect 38243 35244 39304 35272
rect 38243 35241 38255 35244
rect 38197 35235 38255 35241
rect 39298 35232 39304 35244
rect 39356 35232 39362 35284
rect 10502 35204 10508 35216
rect 9140 35176 10508 35204
rect 8389 35071 8447 35077
rect 8389 35037 8401 35071
rect 8435 35037 8447 35071
rect 8389 35031 8447 35037
rect 9140 35000 9168 35176
rect 10502 35164 10508 35176
rect 10560 35164 10566 35216
rect 11330 35204 11336 35216
rect 11072 35176 11336 35204
rect 9306 35096 9312 35148
rect 9364 35136 9370 35148
rect 9364 35108 9996 35136
rect 9364 35096 9370 35108
rect 9968 35068 9996 35108
rect 10042 35096 10048 35148
rect 10100 35136 10106 35148
rect 10597 35139 10655 35145
rect 10597 35136 10609 35139
rect 10100 35108 10609 35136
rect 10100 35096 10106 35108
rect 10597 35105 10609 35108
rect 10643 35105 10655 35139
rect 10597 35099 10655 35105
rect 10870 35096 10876 35148
rect 10928 35136 10934 35148
rect 11072 35145 11100 35176
rect 11330 35164 11336 35176
rect 11388 35164 11394 35216
rect 11514 35164 11520 35216
rect 11572 35204 11578 35216
rect 11572 35176 11836 35204
rect 11572 35164 11578 35176
rect 11057 35139 11115 35145
rect 11057 35136 11069 35139
rect 10928 35108 11069 35136
rect 10928 35096 10934 35108
rect 11057 35105 11069 35108
rect 11103 35105 11115 35139
rect 11057 35099 11115 35105
rect 10413 35071 10471 35077
rect 10413 35068 10425 35071
rect 9968 35040 10425 35068
rect 10413 35037 10425 35040
rect 10459 35037 10471 35071
rect 11808 35068 11836 35176
rect 11882 35164 11888 35216
rect 11940 35204 11946 35216
rect 20070 35204 20076 35216
rect 11940 35176 20076 35204
rect 11940 35164 11946 35176
rect 20070 35164 20076 35176
rect 20128 35164 20134 35216
rect 37369 35207 37427 35213
rect 37369 35173 37381 35207
rect 37415 35173 37427 35207
rect 37369 35167 37427 35173
rect 13081 35139 13139 35145
rect 13081 35136 13093 35139
rect 12406 35108 13093 35136
rect 12406 35068 12434 35108
rect 13081 35105 13093 35108
rect 13127 35105 13139 35139
rect 13081 35099 13139 35105
rect 13170 35096 13176 35148
rect 13228 35136 13234 35148
rect 15381 35139 15439 35145
rect 15381 35136 15393 35139
rect 13228 35108 15393 35136
rect 13228 35096 13234 35108
rect 15381 35105 15393 35108
rect 15427 35105 15439 35139
rect 15381 35099 15439 35105
rect 16850 35096 16856 35148
rect 16908 35136 16914 35148
rect 18693 35139 18751 35145
rect 18693 35136 18705 35139
rect 16908 35108 18705 35136
rect 16908 35096 16914 35108
rect 18693 35105 18705 35108
rect 18739 35105 18751 35139
rect 18693 35099 18751 35105
rect 19334 35096 19340 35148
rect 19392 35136 19398 35148
rect 20441 35139 20499 35145
rect 20441 35136 20453 35139
rect 19392 35108 20453 35136
rect 19392 35096 19398 35108
rect 20441 35105 20453 35108
rect 20487 35136 20499 35139
rect 22278 35136 22284 35148
rect 20487 35108 22284 35136
rect 20487 35105 20499 35108
rect 20441 35099 20499 35105
rect 22278 35096 22284 35108
rect 22336 35096 22342 35148
rect 23017 35139 23075 35145
rect 23017 35105 23029 35139
rect 23063 35136 23075 35139
rect 23474 35136 23480 35148
rect 23063 35108 23480 35136
rect 23063 35105 23075 35108
rect 23017 35099 23075 35105
rect 23474 35096 23480 35108
rect 23532 35096 23538 35148
rect 29086 35096 29092 35148
rect 29144 35136 29150 35148
rect 30193 35139 30251 35145
rect 30193 35136 30205 35139
rect 29144 35108 30205 35136
rect 29144 35096 29150 35108
rect 30193 35105 30205 35108
rect 30239 35105 30251 35139
rect 30193 35099 30251 35105
rect 32309 35139 32367 35145
rect 32309 35105 32321 35139
rect 32355 35136 32367 35139
rect 33226 35136 33232 35148
rect 32355 35108 33232 35136
rect 32355 35105 32367 35108
rect 32309 35099 32367 35105
rect 33226 35096 33232 35108
rect 33284 35136 33290 35148
rect 37384 35136 37412 35167
rect 33284 35108 34468 35136
rect 37384 35108 38056 35136
rect 33284 35096 33290 35108
rect 34440 35080 34468 35108
rect 11808 35040 12434 35068
rect 10413 35031 10471 35037
rect 13998 35028 14004 35080
rect 14056 35068 14062 35080
rect 14277 35071 14335 35077
rect 14277 35068 14289 35071
rect 14056 35040 14289 35068
rect 14056 35028 14062 35040
rect 14277 35037 14289 35040
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 14366 35028 14372 35080
rect 14424 35068 14430 35080
rect 14642 35068 14648 35080
rect 14424 35040 14648 35068
rect 14424 35028 14430 35040
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 17221 35071 17279 35077
rect 17221 35037 17233 35071
rect 17267 35068 17279 35071
rect 17310 35068 17316 35080
rect 17267 35040 17316 35068
rect 17267 35037 17279 35040
rect 17221 35031 17279 35037
rect 17310 35028 17316 35040
rect 17368 35068 17374 35080
rect 17494 35068 17500 35080
rect 17368 35040 17500 35068
rect 17368 35028 17374 35040
rect 17494 35028 17500 35040
rect 17552 35028 17558 35080
rect 20346 35068 20352 35080
rect 17604 35040 20352 35068
rect 9306 35000 9312 35012
rect 4356 34972 9168 35000
rect 9267 34972 9312 35000
rect 9306 34960 9312 34972
rect 9364 34960 9370 35012
rect 9401 35003 9459 35009
rect 9401 34969 9413 35003
rect 9447 35000 9459 35003
rect 9674 35000 9680 35012
rect 9447 34972 9680 35000
rect 9447 34969 9459 34972
rect 9401 34963 9459 34969
rect 9674 34960 9680 34972
rect 9732 34960 9738 35012
rect 9953 35003 10011 35009
rect 9953 34969 9965 35003
rect 9999 35000 10011 35003
rect 10778 35000 10784 35012
rect 9999 34972 10784 35000
rect 9999 34969 10011 34972
rect 9953 34963 10011 34969
rect 10778 34960 10784 34972
rect 10836 35000 10842 35012
rect 12158 35000 12164 35012
rect 10836 34972 12164 35000
rect 10836 34960 10842 34972
rect 12158 34960 12164 34972
rect 12216 34960 12222 35012
rect 12250 34960 12256 35012
rect 12308 35000 12314 35012
rect 13170 35000 13176 35012
rect 12308 34972 13032 35000
rect 13131 34972 13176 35000
rect 12308 34960 12314 34972
rect 4433 34935 4491 34941
rect 4433 34901 4445 34935
rect 4479 34932 4491 34935
rect 4982 34932 4988 34944
rect 4479 34904 4988 34932
rect 4479 34901 4491 34904
rect 4433 34895 4491 34901
rect 4982 34892 4988 34904
rect 5040 34892 5046 34944
rect 6546 34932 6552 34944
rect 6507 34904 6552 34932
rect 6546 34892 6552 34904
rect 6604 34892 6610 34944
rect 8481 34935 8539 34941
rect 8481 34901 8493 34935
rect 8527 34932 8539 34935
rect 12802 34932 12808 34944
rect 8527 34904 12808 34932
rect 8527 34901 8539 34904
rect 8481 34895 8539 34901
rect 12802 34892 12808 34904
rect 12860 34892 12866 34944
rect 13004 34932 13032 34972
rect 13170 34960 13176 34972
rect 13228 34960 13234 35012
rect 13262 34960 13268 35012
rect 13320 35000 13326 35012
rect 13725 35003 13783 35009
rect 13725 35000 13737 35003
rect 13320 34972 13737 35000
rect 13320 34960 13326 34972
rect 13725 34969 13737 34972
rect 13771 34969 13783 35003
rect 15565 35003 15623 35009
rect 15565 35000 15577 35003
rect 13725 34963 13783 34969
rect 14016 34972 15577 35000
rect 14016 34932 14044 34972
rect 15565 34969 15577 34972
rect 15611 34969 15623 35003
rect 15565 34963 15623 34969
rect 13004 34904 14044 34932
rect 14369 34935 14427 34941
rect 14369 34901 14381 34935
rect 14415 34932 14427 34935
rect 14550 34932 14556 34944
rect 14415 34904 14556 34932
rect 14415 34901 14427 34904
rect 14369 34895 14427 34901
rect 14550 34892 14556 34904
rect 14608 34892 14614 34944
rect 14642 34892 14648 34944
rect 14700 34932 14706 34944
rect 17604 34932 17632 35040
rect 20346 35028 20352 35040
rect 20404 35028 20410 35080
rect 22922 35068 22928 35080
rect 22883 35040 22928 35068
rect 22922 35028 22928 35040
rect 22980 35028 22986 35080
rect 34422 35028 34428 35080
rect 34480 35068 34486 35080
rect 34885 35071 34943 35077
rect 34885 35068 34897 35071
rect 34480 35040 34897 35068
rect 34480 35028 34486 35040
rect 34885 35037 34897 35040
rect 34931 35037 34943 35071
rect 37550 35068 37556 35080
rect 37511 35040 37556 35068
rect 34885 35031 34943 35037
rect 37550 35028 37556 35040
rect 37608 35028 37614 35080
rect 38028 35077 38056 35108
rect 38013 35071 38071 35077
rect 38013 35037 38025 35071
rect 38059 35037 38071 35071
rect 38013 35031 38071 35037
rect 17957 35003 18015 35009
rect 17957 34969 17969 35003
rect 18003 34969 18015 35003
rect 17957 34963 18015 34969
rect 14700 34904 17632 34932
rect 17972 34932 18000 34963
rect 18782 34960 18788 35012
rect 18840 35000 18846 35012
rect 19978 35000 19984 35012
rect 18840 34972 19984 35000
rect 18840 34960 18846 34972
rect 19978 34960 19984 34972
rect 20036 34960 20042 35012
rect 20714 35000 20720 35012
rect 20675 34972 20720 35000
rect 20714 34960 20720 34972
rect 20772 34960 20778 35012
rect 20806 34960 20812 35012
rect 20864 35000 20870 35012
rect 23106 35000 23112 35012
rect 20864 34972 21206 35000
rect 22020 34972 23112 35000
rect 20864 34960 20870 34972
rect 22020 34932 22048 34972
rect 23106 34960 23112 34972
rect 23164 34960 23170 35012
rect 30282 34960 30288 35012
rect 30340 35000 30346 35012
rect 31202 35000 31208 35012
rect 30340 34972 30385 35000
rect 31163 34972 31208 35000
rect 30340 34960 30346 34972
rect 31202 34960 31208 34972
rect 31260 34960 31266 35012
rect 32582 35000 32588 35012
rect 32543 34972 32588 35000
rect 32582 34960 32588 34972
rect 32640 34960 32646 35012
rect 33318 34960 33324 35012
rect 33376 34960 33382 35012
rect 34333 35003 34391 35009
rect 34333 34969 34345 35003
rect 34379 35000 34391 35003
rect 34606 35000 34612 35012
rect 34379 34972 34612 35000
rect 34379 34969 34391 34972
rect 34333 34963 34391 34969
rect 34606 34960 34612 34972
rect 34664 34960 34670 35012
rect 34698 34960 34704 35012
rect 34756 35000 34762 35012
rect 35161 35003 35219 35009
rect 35161 35000 35173 35003
rect 34756 34972 35173 35000
rect 34756 34960 34762 34972
rect 35161 34969 35173 34972
rect 35207 34969 35219 35003
rect 36814 35000 36820 35012
rect 36386 34972 36820 35000
rect 35161 34963 35219 34969
rect 36814 34960 36820 34972
rect 36872 34960 36878 35012
rect 36909 35003 36967 35009
rect 36909 34969 36921 35003
rect 36955 34969 36967 35003
rect 36909 34963 36967 34969
rect 17972 34904 22048 34932
rect 14700 34892 14706 34904
rect 22094 34892 22100 34944
rect 22152 34932 22158 34944
rect 22189 34935 22247 34941
rect 22189 34932 22201 34935
rect 22152 34904 22201 34932
rect 22152 34892 22158 34904
rect 22189 34901 22201 34904
rect 22235 34901 22247 34935
rect 22189 34895 22247 34901
rect 33410 34892 33416 34944
rect 33468 34932 33474 34944
rect 36924 34932 36952 34963
rect 33468 34904 36952 34932
rect 33468 34892 33474 34904
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 2222 34688 2228 34740
rect 2280 34728 2286 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 2280 34700 2421 34728
rect 2280 34688 2286 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 4801 34731 4859 34737
rect 4801 34728 4813 34731
rect 2409 34691 2467 34697
rect 2746 34700 4813 34728
rect 2746 34660 2774 34700
rect 4801 34697 4813 34700
rect 4847 34697 4859 34731
rect 4801 34691 4859 34697
rect 5442 34688 5448 34740
rect 5500 34728 5506 34740
rect 10870 34728 10876 34740
rect 5500 34700 10876 34728
rect 5500 34688 5506 34700
rect 10870 34688 10876 34700
rect 10928 34688 10934 34740
rect 10962 34688 10968 34740
rect 11020 34728 11026 34740
rect 19426 34728 19432 34740
rect 11020 34700 11065 34728
rect 11716 34700 16160 34728
rect 11020 34688 11026 34700
rect 3970 34660 3976 34672
rect 1596 34632 2774 34660
rect 3931 34632 3976 34660
rect 1596 34601 1624 34632
rect 3970 34620 3976 34632
rect 4028 34620 4034 34672
rect 6546 34620 6552 34672
rect 6604 34660 6610 34672
rect 9493 34663 9551 34669
rect 9493 34660 9505 34663
rect 6604 34632 9505 34660
rect 6604 34620 6610 34632
rect 9493 34629 9505 34632
rect 9539 34629 9551 34663
rect 9493 34623 9551 34629
rect 10410 34620 10416 34672
rect 10468 34660 10474 34672
rect 11716 34660 11744 34700
rect 10468 34632 11744 34660
rect 11793 34663 11851 34669
rect 10468 34620 10474 34632
rect 11793 34629 11805 34663
rect 11839 34660 11851 34663
rect 11882 34660 11888 34672
rect 11839 34632 11888 34660
rect 11839 34629 11851 34632
rect 11793 34623 11851 34629
rect 11882 34620 11888 34632
rect 11940 34620 11946 34672
rect 12802 34620 12808 34672
rect 12860 34660 12866 34672
rect 13173 34663 13231 34669
rect 13173 34660 13185 34663
rect 12860 34632 13185 34660
rect 12860 34620 12866 34632
rect 13173 34629 13185 34632
rect 13219 34629 13231 34663
rect 13173 34623 13231 34629
rect 13725 34663 13783 34669
rect 13725 34629 13737 34663
rect 13771 34660 13783 34663
rect 13906 34660 13912 34672
rect 13771 34632 13912 34660
rect 13771 34629 13783 34632
rect 13725 34623 13783 34629
rect 13906 34620 13912 34632
rect 13964 34660 13970 34672
rect 14366 34660 14372 34672
rect 13964 34632 14372 34660
rect 13964 34620 13970 34632
rect 14366 34620 14372 34632
rect 14424 34620 14430 34672
rect 14816 34663 14874 34669
rect 14816 34660 14828 34663
rect 14476 34632 14828 34660
rect 1581 34595 1639 34601
rect 1581 34561 1593 34595
rect 1627 34561 1639 34595
rect 2314 34592 2320 34604
rect 2275 34564 2320 34592
rect 1581 34555 1639 34561
rect 2314 34552 2320 34564
rect 2372 34552 2378 34604
rect 3878 34592 3884 34604
rect 3839 34564 3884 34592
rect 3878 34552 3884 34564
rect 3936 34552 3942 34604
rect 4982 34592 4988 34604
rect 4943 34564 4988 34592
rect 4982 34552 4988 34564
rect 5040 34552 5046 34604
rect 8202 34592 8208 34604
rect 8163 34564 8208 34592
rect 8202 34552 8208 34564
rect 8260 34552 8266 34604
rect 8294 34552 8300 34604
rect 8352 34592 8358 34604
rect 8352 34564 8397 34592
rect 8352 34552 8358 34564
rect 10594 34552 10600 34604
rect 10652 34592 10658 34604
rect 10870 34592 10876 34604
rect 10652 34564 10876 34592
rect 10652 34552 10658 34564
rect 10870 34552 10876 34564
rect 10928 34552 10934 34604
rect 11698 34592 11704 34604
rect 11659 34564 11704 34592
rect 11698 34552 11704 34564
rect 11756 34552 11762 34604
rect 14182 34552 14188 34604
rect 14240 34592 14246 34604
rect 14476 34592 14504 34632
rect 14816 34629 14828 34632
rect 14862 34629 14874 34663
rect 14816 34623 14874 34629
rect 15286 34620 15292 34672
rect 15344 34620 15350 34672
rect 14240 34564 14504 34592
rect 14553 34595 14611 34601
rect 14240 34552 14246 34564
rect 14553 34561 14565 34595
rect 14599 34561 14611 34595
rect 14553 34555 14611 34561
rect 9401 34527 9459 34533
rect 9401 34493 9413 34527
rect 9447 34524 9459 34527
rect 10042 34524 10048 34536
rect 9447 34496 10048 34524
rect 9447 34493 9459 34496
rect 9401 34487 9459 34493
rect 10042 34484 10048 34496
rect 10100 34484 10106 34536
rect 10413 34527 10471 34533
rect 10413 34493 10425 34527
rect 10459 34524 10471 34527
rect 10962 34524 10968 34536
rect 10459 34496 10968 34524
rect 10459 34493 10471 34496
rect 10413 34487 10471 34493
rect 10962 34484 10968 34496
rect 11020 34484 11026 34536
rect 13078 34524 13084 34536
rect 13039 34496 13084 34524
rect 13078 34484 13084 34496
rect 13136 34484 13142 34536
rect 14458 34416 14464 34468
rect 14516 34456 14522 34468
rect 14568 34456 14596 34555
rect 16132 34524 16160 34700
rect 18616 34700 19432 34728
rect 18616 34660 18644 34700
rect 19426 34688 19432 34700
rect 19484 34688 19490 34740
rect 19518 34688 19524 34740
rect 19576 34728 19582 34740
rect 20257 34731 20315 34737
rect 20257 34728 20269 34731
rect 19576 34700 20269 34728
rect 19576 34688 19582 34700
rect 20257 34697 20269 34700
rect 20303 34728 20315 34731
rect 20714 34728 20720 34740
rect 20303 34700 20720 34728
rect 20303 34697 20315 34700
rect 20257 34691 20315 34697
rect 20714 34688 20720 34700
rect 20772 34688 20778 34740
rect 22186 34728 22192 34740
rect 20824 34700 22192 34728
rect 18782 34660 18788 34672
rect 18524 34632 18644 34660
rect 18743 34632 18788 34660
rect 18524 34601 18552 34632
rect 18782 34620 18788 34632
rect 18840 34620 18846 34672
rect 20824 34601 20852 34700
rect 22186 34688 22192 34700
rect 22244 34688 22250 34740
rect 24305 34731 24363 34737
rect 24305 34728 24317 34731
rect 22296 34700 24317 34728
rect 20898 34620 20904 34672
rect 20956 34660 20962 34672
rect 22296 34660 22324 34700
rect 24305 34697 24317 34700
rect 24351 34697 24363 34731
rect 31478 34728 31484 34740
rect 31439 34700 31484 34728
rect 24305 34691 24363 34697
rect 31478 34688 31484 34700
rect 31536 34688 31542 34740
rect 33226 34728 33232 34740
rect 32324 34700 33232 34728
rect 24762 34660 24768 34672
rect 20956 34632 21001 34660
rect 22066 34632 22324 34660
rect 24058 34632 24768 34660
rect 20956 34620 20962 34632
rect 18509 34595 18567 34601
rect 18509 34561 18521 34595
rect 18555 34561 18567 34595
rect 20809 34595 20867 34601
rect 18509 34555 18567 34561
rect 19904 34524 19932 34578
rect 20809 34561 20821 34595
rect 20855 34561 20867 34595
rect 22066 34592 22094 34632
rect 24762 34620 24768 34632
rect 24820 34620 24826 34672
rect 30466 34620 30472 34672
rect 30524 34660 30530 34672
rect 30745 34663 30803 34669
rect 30745 34660 30757 34663
rect 30524 34632 30757 34660
rect 30524 34620 30530 34632
rect 30745 34629 30757 34632
rect 30791 34629 30803 34663
rect 30745 34623 30803 34629
rect 20809 34555 20867 34561
rect 20916 34564 22094 34592
rect 16132 34496 19932 34524
rect 19978 34484 19984 34536
rect 20036 34524 20042 34536
rect 20916 34524 20944 34564
rect 22278 34552 22284 34604
rect 22336 34592 22342 34604
rect 22557 34595 22615 34601
rect 22557 34592 22569 34595
rect 22336 34564 22569 34592
rect 22336 34552 22342 34564
rect 22557 34561 22569 34564
rect 22603 34561 22615 34595
rect 27154 34592 27160 34604
rect 27115 34564 27160 34592
rect 22557 34555 22615 34561
rect 27154 34552 27160 34564
rect 27212 34552 27218 34604
rect 28534 34552 28540 34604
rect 28592 34552 28598 34604
rect 30006 34592 30012 34604
rect 29967 34564 30012 34592
rect 30006 34552 30012 34564
rect 30064 34552 30070 34604
rect 31018 34552 31024 34604
rect 31076 34592 31082 34604
rect 32324 34601 32352 34700
rect 33226 34688 33232 34700
rect 33284 34688 33290 34740
rect 33962 34688 33968 34740
rect 34020 34728 34026 34740
rect 34057 34731 34115 34737
rect 34057 34728 34069 34731
rect 34020 34700 34069 34728
rect 34020 34688 34026 34700
rect 34057 34697 34069 34700
rect 34103 34697 34115 34731
rect 38838 34728 38844 34740
rect 34057 34691 34115 34697
rect 35452 34700 38844 34728
rect 35452 34660 35480 34700
rect 38838 34688 38844 34700
rect 38896 34688 38902 34740
rect 35848 34669 35854 34672
rect 35713 34663 35771 34669
rect 35713 34660 35725 34663
rect 33810 34632 35480 34660
rect 35544 34632 35725 34660
rect 31389 34595 31447 34601
rect 31389 34592 31401 34595
rect 31076 34564 31401 34592
rect 31076 34552 31082 34564
rect 31389 34561 31401 34564
rect 31435 34561 31447 34595
rect 31389 34555 31447 34561
rect 32309 34595 32367 34601
rect 32309 34561 32321 34595
rect 32355 34561 32367 34595
rect 32309 34555 32367 34561
rect 35250 34552 35256 34604
rect 35308 34592 35314 34604
rect 35544 34592 35572 34632
rect 35713 34629 35725 34632
rect 35759 34629 35771 34663
rect 35713 34623 35771 34629
rect 35805 34663 35854 34669
rect 35805 34629 35817 34663
rect 35851 34629 35854 34663
rect 35805 34623 35854 34629
rect 35848 34620 35854 34623
rect 35906 34620 35912 34672
rect 35308 34564 35572 34592
rect 35308 34552 35314 34564
rect 37918 34552 37924 34604
rect 37976 34592 37982 34604
rect 38013 34595 38071 34601
rect 38013 34592 38025 34595
rect 37976 34564 38025 34592
rect 37976 34552 37982 34564
rect 38013 34561 38025 34564
rect 38059 34561 38071 34595
rect 38013 34555 38071 34561
rect 20036 34496 20944 34524
rect 22833 34527 22891 34533
rect 20036 34484 20042 34496
rect 22833 34493 22845 34527
rect 22879 34524 22891 34527
rect 29178 34524 29184 34536
rect 22879 34496 23888 34524
rect 29139 34496 29184 34524
rect 22879 34493 22891 34496
rect 22833 34487 22891 34493
rect 18230 34456 18236 34468
rect 14516 34428 14596 34456
rect 16224 34428 18236 34456
rect 14516 34416 14522 34428
rect 1762 34388 1768 34400
rect 1723 34360 1768 34388
rect 1762 34348 1768 34360
rect 1820 34348 1826 34400
rect 11054 34348 11060 34400
rect 11112 34388 11118 34400
rect 16224 34388 16252 34428
rect 18230 34416 18236 34428
rect 18288 34416 18294 34468
rect 23860 34456 23888 34496
rect 29178 34484 29184 34496
rect 29236 34484 29242 34536
rect 29270 34484 29276 34536
rect 29328 34524 29334 34536
rect 36170 34524 36176 34536
rect 29328 34496 36176 34524
rect 29328 34484 29334 34496
rect 36170 34484 36176 34496
rect 36228 34484 36234 34536
rect 24578 34456 24584 34468
rect 19812 34428 22094 34456
rect 23860 34428 24584 34456
rect 11112 34360 16252 34388
rect 11112 34348 11118 34360
rect 16298 34348 16304 34400
rect 16356 34388 16362 34400
rect 16356 34360 16401 34388
rect 16356 34348 16362 34360
rect 16666 34348 16672 34400
rect 16724 34388 16730 34400
rect 19812 34388 19840 34428
rect 16724 34360 19840 34388
rect 22066 34388 22094 34428
rect 24578 34416 24584 34428
rect 24636 34416 24642 34468
rect 23566 34388 23572 34400
rect 22066 34360 23572 34388
rect 16724 34348 16730 34360
rect 23566 34348 23572 34360
rect 23624 34388 23630 34400
rect 24026 34388 24032 34400
rect 23624 34360 24032 34388
rect 23624 34348 23630 34360
rect 24026 34348 24032 34360
rect 24084 34348 24090 34400
rect 27420 34391 27478 34397
rect 27420 34357 27432 34391
rect 27466 34388 27478 34391
rect 28994 34388 29000 34400
rect 27466 34360 29000 34388
rect 27466 34357 27478 34360
rect 27420 34351 27478 34357
rect 28994 34348 29000 34360
rect 29052 34348 29058 34400
rect 32572 34391 32630 34397
rect 32572 34357 32584 34391
rect 32618 34388 32630 34391
rect 32674 34388 32680 34400
rect 32618 34360 32680 34388
rect 32618 34357 32630 34360
rect 32572 34351 32630 34357
rect 32674 34348 32680 34360
rect 32732 34348 32738 34400
rect 38194 34388 38200 34400
rect 38155 34360 38200 34388
rect 38194 34348 38200 34360
rect 38252 34348 38258 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 9582 34144 9588 34196
rect 9640 34184 9646 34196
rect 9640 34156 13124 34184
rect 9640 34144 9646 34156
rect 11422 34076 11428 34128
rect 11480 34116 11486 34128
rect 12250 34116 12256 34128
rect 11480 34088 12256 34116
rect 11480 34076 11486 34088
rect 12250 34076 12256 34088
rect 12308 34076 12314 34128
rect 13096 34116 13124 34156
rect 13170 34144 13176 34196
rect 13228 34184 13234 34196
rect 13265 34187 13323 34193
rect 13265 34184 13277 34187
rect 13228 34156 13277 34184
rect 13228 34144 13234 34156
rect 13265 34153 13277 34156
rect 13311 34153 13323 34187
rect 13265 34147 13323 34153
rect 13354 34144 13360 34196
rect 13412 34184 13418 34196
rect 14274 34184 14280 34196
rect 13412 34156 14280 34184
rect 13412 34144 13418 34156
rect 14274 34144 14280 34156
rect 14332 34144 14338 34196
rect 14369 34187 14427 34193
rect 14369 34153 14381 34187
rect 14415 34184 14427 34187
rect 15194 34184 15200 34196
rect 14415 34156 15200 34184
rect 14415 34153 14427 34156
rect 14369 34147 14427 34153
rect 15194 34144 15200 34156
rect 15252 34144 15258 34196
rect 15488 34156 18184 34184
rect 15488 34116 15516 34156
rect 13096 34088 15516 34116
rect 18156 34116 18184 34156
rect 18230 34144 18236 34196
rect 18288 34184 18294 34196
rect 19978 34184 19984 34196
rect 18288 34156 19984 34184
rect 18288 34144 18294 34156
rect 19978 34144 19984 34156
rect 20036 34144 20042 34196
rect 25501 34187 25559 34193
rect 25501 34153 25513 34187
rect 25547 34184 25559 34187
rect 27338 34184 27344 34196
rect 25547 34156 27344 34184
rect 25547 34153 25559 34156
rect 25501 34147 25559 34153
rect 27338 34144 27344 34156
rect 27396 34144 27402 34196
rect 30009 34187 30067 34193
rect 30009 34153 30021 34187
rect 30055 34184 30067 34187
rect 30282 34184 30288 34196
rect 30055 34156 30288 34184
rect 30055 34153 30067 34156
rect 30009 34147 30067 34153
rect 30282 34144 30288 34156
rect 30340 34144 30346 34196
rect 34149 34187 34207 34193
rect 34149 34153 34161 34187
rect 34195 34184 34207 34187
rect 35710 34184 35716 34196
rect 34195 34156 35716 34184
rect 34195 34153 34207 34156
rect 34149 34147 34207 34153
rect 35710 34144 35716 34156
rect 35768 34144 35774 34196
rect 18156 34088 19748 34116
rect 15381 34051 15439 34057
rect 15381 34017 15393 34051
rect 15427 34048 15439 34051
rect 16850 34048 16856 34060
rect 15427 34020 16856 34048
rect 15427 34017 15439 34020
rect 15381 34011 15439 34017
rect 2130 33980 2136 33992
rect 2091 33952 2136 33980
rect 2130 33940 2136 33952
rect 2188 33940 2194 33992
rect 2774 33940 2780 33992
rect 2832 33980 2838 33992
rect 2832 33952 2877 33980
rect 2832 33940 2838 33952
rect 6914 33940 6920 33992
rect 6972 33980 6978 33992
rect 9125 33983 9183 33989
rect 9125 33980 9137 33983
rect 6972 33952 9137 33980
rect 6972 33940 6978 33952
rect 9125 33949 9137 33952
rect 9171 33949 9183 33983
rect 9125 33943 9183 33949
rect 11333 33983 11391 33989
rect 11333 33949 11345 33983
rect 11379 33980 11391 33983
rect 11698 33980 11704 33992
rect 11379 33952 11704 33980
rect 11379 33949 11391 33952
rect 11333 33943 11391 33949
rect 11698 33940 11704 33952
rect 11756 33980 11762 33992
rect 11977 33983 12035 33989
rect 11977 33980 11989 33983
rect 11756 33952 11989 33980
rect 11756 33940 11762 33952
rect 11977 33949 11989 33952
rect 12023 33980 12035 33983
rect 12158 33980 12164 33992
rect 12023 33952 12164 33980
rect 12023 33949 12035 33952
rect 11977 33943 12035 33949
rect 12158 33940 12164 33952
rect 12216 33940 12222 33992
rect 12250 33940 12256 33992
rect 12308 33980 12314 33992
rect 13078 33980 13084 33992
rect 12308 33952 13084 33980
rect 12308 33940 12314 33952
rect 13078 33940 13084 33952
rect 13136 33940 13142 33992
rect 13173 33983 13231 33989
rect 13173 33949 13185 33983
rect 13219 33949 13231 33983
rect 14550 33980 14556 33992
rect 14511 33952 14556 33980
rect 13173 33943 13231 33949
rect 11425 33915 11483 33921
rect 11425 33881 11437 33915
rect 11471 33912 11483 33915
rect 13188 33912 13216 33943
rect 14550 33940 14556 33952
rect 14608 33940 14614 33992
rect 11471 33884 12296 33912
rect 13188 33884 14320 33912
rect 11471 33881 11483 33884
rect 11425 33875 11483 33881
rect 1578 33804 1584 33856
rect 1636 33844 1642 33856
rect 1949 33847 2007 33853
rect 1949 33844 1961 33847
rect 1636 33816 1961 33844
rect 1636 33804 1642 33816
rect 1949 33813 1961 33816
rect 1995 33813 2007 33847
rect 2866 33844 2872 33856
rect 2827 33816 2872 33844
rect 1949 33807 2007 33813
rect 2866 33804 2872 33816
rect 2924 33804 2930 33856
rect 9217 33847 9275 33853
rect 9217 33813 9229 33847
rect 9263 33844 9275 33847
rect 11146 33844 11152 33856
rect 9263 33816 11152 33844
rect 9263 33813 9275 33816
rect 9217 33807 9275 33813
rect 11146 33804 11152 33816
rect 11204 33804 11210 33856
rect 12066 33844 12072 33856
rect 12027 33816 12072 33844
rect 12066 33804 12072 33816
rect 12124 33804 12130 33856
rect 12268 33844 12296 33884
rect 13630 33844 13636 33856
rect 12268 33816 13636 33844
rect 13630 33804 13636 33816
rect 13688 33804 13694 33856
rect 14292 33844 14320 33884
rect 14458 33872 14464 33924
rect 14516 33912 14522 33924
rect 15396 33912 15424 34011
rect 16850 34008 16856 34020
rect 16908 34008 16914 34060
rect 19334 34008 19340 34060
rect 19392 34048 19398 34060
rect 19613 34051 19671 34057
rect 19613 34048 19625 34051
rect 19392 34020 19625 34048
rect 19392 34008 19398 34020
rect 19613 34017 19625 34020
rect 19659 34017 19671 34051
rect 19720 34048 19748 34088
rect 32674 34076 32680 34128
rect 32732 34116 32738 34128
rect 32732 34088 35020 34116
rect 32732 34076 32738 34088
rect 19889 34051 19947 34057
rect 19889 34048 19901 34051
rect 19720 34020 19901 34048
rect 19613 34011 19671 34017
rect 19889 34017 19901 34020
rect 19935 34048 19947 34051
rect 22094 34048 22100 34060
rect 19935 34020 22100 34048
rect 19935 34017 19947 34020
rect 19889 34011 19947 34017
rect 22094 34008 22100 34020
rect 22152 34008 22158 34060
rect 22830 34008 22836 34060
rect 22888 34048 22894 34060
rect 22888 34020 28580 34048
rect 22888 34008 22894 34020
rect 17678 33940 17684 33992
rect 17736 33980 17742 33992
rect 18598 33980 18604 33992
rect 17736 33952 18604 33980
rect 17736 33940 17742 33952
rect 18598 33940 18604 33952
rect 18656 33940 18662 33992
rect 22002 33940 22008 33992
rect 22060 33980 22066 33992
rect 22189 33983 22247 33989
rect 22189 33980 22201 33983
rect 22060 33952 22201 33980
rect 22060 33940 22066 33952
rect 22189 33949 22201 33952
rect 22235 33949 22247 33983
rect 25406 33980 25412 33992
rect 25319 33952 25412 33980
rect 22189 33943 22247 33949
rect 25406 33940 25412 33952
rect 25464 33980 25470 33992
rect 26142 33980 26148 33992
rect 25464 33952 26148 33980
rect 25464 33940 25470 33952
rect 26142 33940 26148 33952
rect 26200 33940 26206 33992
rect 14516 33884 15424 33912
rect 15657 33915 15715 33921
rect 14516 33872 14522 33884
rect 15657 33881 15669 33915
rect 15703 33912 15715 33915
rect 15930 33912 15936 33924
rect 15703 33884 15936 33912
rect 15703 33881 15715 33884
rect 15657 33875 15715 33881
rect 15930 33872 15936 33884
rect 15988 33872 15994 33924
rect 16114 33872 16120 33924
rect 16172 33872 16178 33924
rect 19610 33912 19616 33924
rect 16960 33884 19616 33912
rect 15562 33844 15568 33856
rect 14292 33816 15568 33844
rect 15562 33804 15568 33816
rect 15620 33804 15626 33856
rect 15746 33804 15752 33856
rect 15804 33844 15810 33856
rect 16960 33844 16988 33884
rect 19610 33872 19616 33884
rect 19668 33872 19674 33924
rect 19720 33884 20378 33912
rect 17126 33844 17132 33856
rect 15804 33816 16988 33844
rect 17087 33816 17132 33844
rect 15804 33804 15810 33816
rect 17126 33804 17132 33816
rect 17184 33804 17190 33856
rect 17402 33804 17408 33856
rect 17460 33844 17466 33856
rect 19720 33844 19748 33884
rect 21174 33872 21180 33924
rect 21232 33912 21238 33924
rect 22094 33912 22100 33924
rect 21232 33884 22100 33912
rect 21232 33872 21238 33884
rect 22094 33872 22100 33884
rect 22152 33872 22158 33924
rect 22462 33912 22468 33924
rect 22423 33884 22468 33912
rect 22462 33872 22468 33884
rect 22520 33872 22526 33924
rect 24394 33912 24400 33924
rect 23690 33884 24400 33912
rect 24394 33872 24400 33884
rect 24452 33872 24458 33924
rect 27430 33912 27436 33924
rect 27391 33884 27436 33912
rect 27430 33872 27436 33884
rect 27488 33872 27494 33924
rect 27522 33872 27528 33924
rect 27580 33912 27586 33924
rect 28442 33912 28448 33924
rect 27580 33884 27625 33912
rect 28403 33884 28448 33912
rect 27580 33872 27586 33884
rect 28442 33872 28448 33884
rect 28500 33872 28506 33924
rect 28552 33912 28580 34020
rect 30466 34008 30472 34060
rect 30524 34048 30530 34060
rect 31389 34051 31447 34057
rect 31389 34048 31401 34051
rect 30524 34020 31401 34048
rect 30524 34008 30530 34020
rect 31389 34017 31401 34020
rect 31435 34017 31447 34051
rect 31389 34011 31447 34017
rect 34422 34008 34428 34060
rect 34480 34048 34486 34060
rect 34885 34051 34943 34057
rect 34885 34048 34897 34051
rect 34480 34020 34897 34048
rect 34480 34008 34486 34020
rect 34885 34017 34897 34020
rect 34931 34017 34943 34051
rect 34992 34048 35020 34088
rect 36633 34051 36691 34057
rect 36633 34048 36645 34051
rect 34992 34020 36645 34048
rect 34885 34011 34943 34017
rect 36633 34017 36645 34020
rect 36679 34017 36691 34051
rect 36633 34011 36691 34017
rect 29917 33983 29975 33989
rect 29917 33949 29929 33983
rect 29963 33980 29975 33983
rect 31110 33980 31116 33992
rect 29963 33952 31116 33980
rect 29963 33949 29975 33952
rect 29917 33943 29975 33949
rect 31110 33940 31116 33952
rect 31168 33940 31174 33992
rect 34057 33983 34115 33989
rect 34057 33949 34069 33983
rect 34103 33980 34115 33983
rect 34698 33980 34704 33992
rect 34103 33952 34704 33980
rect 34103 33949 34115 33952
rect 34057 33943 34115 33949
rect 34698 33940 34704 33952
rect 34756 33940 34762 33992
rect 31665 33915 31723 33921
rect 31665 33912 31677 33915
rect 28552 33884 31677 33912
rect 31665 33881 31677 33884
rect 31711 33881 31723 33915
rect 31665 33875 31723 33881
rect 32122 33872 32128 33924
rect 32180 33872 32186 33924
rect 34514 33872 34520 33924
rect 34572 33912 34578 33924
rect 35161 33915 35219 33921
rect 35161 33912 35173 33915
rect 34572 33884 35173 33912
rect 34572 33872 34578 33884
rect 35161 33881 35173 33884
rect 35207 33881 35219 33915
rect 35161 33875 35219 33881
rect 35894 33872 35900 33924
rect 35952 33872 35958 33924
rect 17460 33816 19748 33844
rect 17460 33804 17466 33816
rect 19886 33804 19892 33856
rect 19944 33844 19950 33856
rect 21361 33847 21419 33853
rect 21361 33844 21373 33847
rect 19944 33816 21373 33844
rect 19944 33804 19950 33816
rect 21361 33813 21373 33816
rect 21407 33813 21419 33847
rect 21361 33807 21419 33813
rect 23937 33847 23995 33853
rect 23937 33813 23949 33847
rect 23983 33844 23995 33847
rect 24210 33844 24216 33856
rect 23983 33816 24216 33844
rect 23983 33813 23995 33816
rect 23937 33807 23995 33813
rect 24210 33804 24216 33816
rect 24268 33804 24274 33856
rect 31110 33804 31116 33856
rect 31168 33844 31174 33856
rect 33137 33847 33195 33853
rect 33137 33844 33149 33847
rect 31168 33816 33149 33844
rect 31168 33804 31174 33816
rect 33137 33813 33149 33816
rect 33183 33813 33195 33847
rect 33137 33807 33195 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 9030 33600 9036 33652
rect 9088 33640 9094 33652
rect 11793 33643 11851 33649
rect 9088 33612 11744 33640
rect 9088 33600 9094 33612
rect 4525 33575 4583 33581
rect 4525 33541 4537 33575
rect 4571 33572 4583 33575
rect 4614 33572 4620 33584
rect 4571 33544 4620 33572
rect 4571 33541 4583 33544
rect 4525 33535 4583 33541
rect 4614 33532 4620 33544
rect 4672 33532 4678 33584
rect 8018 33572 8024 33584
rect 7979 33544 8024 33572
rect 8018 33532 8024 33544
rect 8076 33532 8082 33584
rect 8113 33575 8171 33581
rect 8113 33541 8125 33575
rect 8159 33572 8171 33575
rect 9214 33572 9220 33584
rect 8159 33544 9220 33572
rect 8159 33541 8171 33544
rect 8113 33535 8171 33541
rect 9214 33532 9220 33544
rect 9272 33532 9278 33584
rect 10410 33572 10416 33584
rect 10371 33544 10416 33572
rect 10410 33532 10416 33544
rect 10468 33532 10474 33584
rect 11716 33572 11744 33612
rect 11793 33609 11805 33643
rect 11839 33640 11851 33643
rect 11974 33640 11980 33652
rect 11839 33612 11980 33640
rect 11839 33609 11851 33612
rect 11793 33603 11851 33609
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 13078 33600 13084 33652
rect 13136 33640 13142 33652
rect 13136 33612 16252 33640
rect 13136 33600 13142 33612
rect 16114 33572 16120 33584
rect 11716 33544 12480 33572
rect 8662 33464 8668 33516
rect 8720 33504 8726 33516
rect 9125 33507 9183 33513
rect 8720 33476 8765 33504
rect 8720 33464 8726 33476
rect 9125 33473 9137 33507
rect 9171 33473 9183 33507
rect 9125 33467 9183 33473
rect 11701 33507 11759 33513
rect 11701 33473 11713 33507
rect 11747 33504 11759 33507
rect 12158 33504 12164 33516
rect 11747 33476 12164 33504
rect 11747 33473 11759 33476
rect 11701 33467 11759 33473
rect 4433 33439 4491 33445
rect 4433 33405 4445 33439
rect 4479 33436 4491 33439
rect 5074 33436 5080 33448
rect 4479 33408 5080 33436
rect 4479 33405 4491 33408
rect 4433 33399 4491 33405
rect 5074 33396 5080 33408
rect 5132 33396 5138 33448
rect 5350 33436 5356 33448
rect 5311 33408 5356 33436
rect 5350 33396 5356 33408
rect 5408 33396 5414 33448
rect 6730 33396 6736 33448
rect 6788 33436 6794 33448
rect 9140 33436 9168 33467
rect 12158 33464 12164 33476
rect 12216 33504 12222 33516
rect 12345 33507 12403 33513
rect 12345 33504 12357 33507
rect 12216 33476 12357 33504
rect 12216 33464 12222 33476
rect 12345 33473 12357 33476
rect 12391 33473 12403 33507
rect 12452 33504 12480 33544
rect 13096 33544 16120 33572
rect 13096 33504 13124 33544
rect 16114 33532 16120 33544
rect 16172 33532 16178 33584
rect 16224 33572 16252 33612
rect 17126 33600 17132 33652
rect 17184 33640 17190 33652
rect 18598 33640 18604 33652
rect 17184 33612 18460 33640
rect 18559 33612 18604 33640
rect 17184 33600 17190 33612
rect 18432 33572 18460 33612
rect 18598 33600 18604 33612
rect 18656 33600 18662 33652
rect 19058 33600 19064 33652
rect 19116 33640 19122 33652
rect 20993 33643 21051 33649
rect 20993 33640 21005 33643
rect 19116 33612 21005 33640
rect 19116 33600 19122 33612
rect 20993 33609 21005 33612
rect 21039 33609 21051 33643
rect 20993 33603 21051 33609
rect 22094 33600 22100 33652
rect 22152 33640 22158 33652
rect 24946 33640 24952 33652
rect 22152 33612 24952 33640
rect 22152 33600 22158 33612
rect 24946 33600 24952 33612
rect 25004 33600 25010 33652
rect 27430 33600 27436 33652
rect 27488 33640 27494 33652
rect 35253 33643 35311 33649
rect 35253 33640 35265 33643
rect 27488 33612 35265 33640
rect 27488 33600 27494 33612
rect 35253 33609 35265 33612
rect 35299 33609 35311 33643
rect 35253 33603 35311 33609
rect 19521 33575 19579 33581
rect 19521 33572 19533 33575
rect 16224 33544 17618 33572
rect 18432 33544 19533 33572
rect 19521 33541 19533 33544
rect 19567 33541 19579 33575
rect 19521 33535 19579 33541
rect 19978 33532 19984 33584
rect 20036 33532 20042 33584
rect 24486 33532 24492 33584
rect 24544 33532 24550 33584
rect 25038 33532 25044 33584
rect 25096 33572 25102 33584
rect 25685 33575 25743 33581
rect 25685 33572 25697 33575
rect 25096 33544 25697 33572
rect 25096 33532 25102 33544
rect 25685 33541 25697 33544
rect 25731 33541 25743 33575
rect 25685 33535 25743 33541
rect 30006 33532 30012 33584
rect 30064 33572 30070 33584
rect 33781 33575 33839 33581
rect 30064 33544 32996 33572
rect 30064 33532 30070 33544
rect 32968 33516 32996 33544
rect 33781 33541 33793 33575
rect 33827 33572 33839 33575
rect 34422 33572 34428 33584
rect 33827 33544 34428 33572
rect 33827 33541 33839 33544
rect 33781 33535 33839 33541
rect 34422 33532 34428 33544
rect 34480 33532 34486 33584
rect 35526 33532 35532 33584
rect 35584 33572 35590 33584
rect 35989 33575 36047 33581
rect 35989 33572 36001 33575
rect 35584 33544 36001 33572
rect 35584 33532 35590 33544
rect 35989 33541 36001 33544
rect 36035 33541 36047 33575
rect 35989 33535 36047 33541
rect 12452 33476 13124 33504
rect 13449 33507 13507 33513
rect 12345 33467 12403 33473
rect 13449 33473 13461 33507
rect 13495 33504 13507 33507
rect 13722 33504 13728 33516
rect 13495 33476 13728 33504
rect 13495 33473 13507 33476
rect 13449 33467 13507 33473
rect 13722 33464 13728 33476
rect 13780 33464 13786 33516
rect 14185 33507 14243 33513
rect 14185 33473 14197 33507
rect 14231 33504 14243 33507
rect 16666 33504 16672 33516
rect 14231 33476 16672 33504
rect 14231 33473 14243 33476
rect 14185 33467 14243 33473
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 16850 33504 16856 33516
rect 16811 33476 16856 33504
rect 16850 33464 16856 33476
rect 16908 33464 16914 33516
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33473 19303 33507
rect 19245 33467 19303 33473
rect 6788 33408 9168 33436
rect 6788 33396 6794 33408
rect 10134 33396 10140 33448
rect 10192 33436 10198 33448
rect 10321 33439 10379 33445
rect 10321 33436 10333 33439
rect 10192 33408 10333 33436
rect 10192 33396 10198 33408
rect 10321 33405 10333 33408
rect 10367 33405 10379 33439
rect 10321 33399 10379 33405
rect 10502 33396 10508 33448
rect 10560 33436 10566 33448
rect 10597 33439 10655 33445
rect 10597 33436 10609 33439
rect 10560 33408 10609 33436
rect 10560 33396 10566 33408
rect 10597 33405 10609 33408
rect 10643 33405 10655 33439
rect 10597 33399 10655 33405
rect 10612 33368 10640 33399
rect 10686 33396 10692 33448
rect 10744 33436 10750 33448
rect 12250 33436 12256 33448
rect 10744 33408 12256 33436
rect 10744 33396 10750 33408
rect 12250 33396 12256 33408
rect 12308 33396 12314 33448
rect 12437 33439 12495 33445
rect 12437 33405 12449 33439
rect 12483 33436 12495 33439
rect 12483 33408 13308 33436
rect 12483 33405 12495 33408
rect 12437 33399 12495 33405
rect 13170 33368 13176 33380
rect 10612 33340 13176 33368
rect 13170 33328 13176 33340
rect 13228 33328 13234 33380
rect 13280 33368 13308 33408
rect 14642 33396 14648 33448
rect 14700 33436 14706 33448
rect 15930 33436 15936 33448
rect 14700 33408 15936 33436
rect 14700 33396 14706 33408
rect 15930 33396 15936 33408
rect 15988 33396 15994 33448
rect 16390 33396 16396 33448
rect 16448 33436 16454 33448
rect 17129 33439 17187 33445
rect 17129 33436 17141 33439
rect 16448 33408 17141 33436
rect 16448 33396 16454 33408
rect 17129 33405 17141 33408
rect 17175 33436 17187 33439
rect 17770 33436 17776 33448
rect 17175 33408 17776 33436
rect 17175 33405 17187 33408
rect 17129 33399 17187 33405
rect 17770 33396 17776 33408
rect 17828 33396 17834 33448
rect 15746 33368 15752 33380
rect 13280 33340 15752 33368
rect 15746 33328 15752 33340
rect 15804 33328 15810 33380
rect 9217 33303 9275 33309
rect 9217 33269 9229 33303
rect 9263 33300 9275 33303
rect 9582 33300 9588 33312
rect 9263 33272 9588 33300
rect 9263 33269 9275 33272
rect 9217 33263 9275 33269
rect 9582 33260 9588 33272
rect 9640 33260 9646 33312
rect 13262 33300 13268 33312
rect 13223 33272 13268 33300
rect 13262 33260 13268 33272
rect 13320 33260 13326 33312
rect 13354 33260 13360 33312
rect 13412 33300 13418 33312
rect 14277 33303 14335 33309
rect 14277 33300 14289 33303
rect 13412 33272 14289 33300
rect 13412 33260 13418 33272
rect 14277 33269 14289 33272
rect 14323 33269 14335 33303
rect 19260 33300 19288 33467
rect 27154 33464 27160 33516
rect 27212 33504 27218 33516
rect 28445 33507 28503 33513
rect 28445 33504 28457 33507
rect 27212 33476 28457 33504
rect 27212 33464 27218 33476
rect 28445 33473 28457 33476
rect 28491 33473 28503 33507
rect 28445 33467 28503 33473
rect 29822 33464 29828 33516
rect 29880 33464 29886 33516
rect 30929 33507 30987 33513
rect 30929 33473 30941 33507
rect 30975 33504 30987 33507
rect 31110 33504 31116 33516
rect 30975 33476 31116 33504
rect 30975 33473 30987 33476
rect 30929 33467 30987 33473
rect 31110 33464 31116 33476
rect 31168 33464 31174 33516
rect 32950 33504 32956 33516
rect 32911 33476 32956 33504
rect 32950 33464 32956 33476
rect 33008 33464 33014 33516
rect 35161 33507 35219 33513
rect 35161 33473 35173 33507
rect 35207 33473 35219 33507
rect 35161 33467 35219 33473
rect 21726 33436 21732 33448
rect 20824 33408 21732 33436
rect 20824 33312 20852 33408
rect 21726 33396 21732 33408
rect 21784 33436 21790 33448
rect 22002 33436 22008 33448
rect 21784 33408 22008 33436
rect 21784 33396 21790 33408
rect 22002 33396 22008 33408
rect 22060 33436 22066 33448
rect 23201 33439 23259 33445
rect 23201 33436 23213 33439
rect 22060 33408 23213 33436
rect 22060 33396 22066 33408
rect 23201 33405 23213 33408
rect 23247 33405 23259 33439
rect 23201 33399 23259 33405
rect 23477 33439 23535 33445
rect 23477 33405 23489 33439
rect 23523 33436 23535 33439
rect 24210 33436 24216 33448
rect 23523 33408 24216 33436
rect 23523 33405 23535 33408
rect 23477 33399 23535 33405
rect 24210 33396 24216 33408
rect 24268 33396 24274 33448
rect 25590 33436 25596 33448
rect 25551 33408 25596 33436
rect 25590 33396 25596 33408
rect 25648 33396 25654 33448
rect 26234 33436 26240 33448
rect 26195 33408 26240 33436
rect 26234 33396 26240 33408
rect 26292 33396 26298 33448
rect 28718 33436 28724 33448
rect 28679 33408 28724 33436
rect 28718 33396 28724 33408
rect 28776 33396 28782 33448
rect 29914 33396 29920 33448
rect 29972 33436 29978 33448
rect 30469 33439 30527 33445
rect 30469 33436 30481 33439
rect 29972 33408 30481 33436
rect 29972 33396 29978 33408
rect 30469 33405 30481 33408
rect 30515 33405 30527 33439
rect 30469 33399 30527 33405
rect 35176 33368 35204 33467
rect 35894 33396 35900 33448
rect 35952 33436 35958 33448
rect 36170 33436 36176 33448
rect 35952 33408 35997 33436
rect 36131 33408 36176 33436
rect 35952 33396 35958 33408
rect 36170 33396 36176 33408
rect 36228 33396 36234 33448
rect 38102 33368 38108 33380
rect 35176 33340 38108 33368
rect 38102 33328 38108 33340
rect 38160 33328 38166 33380
rect 20806 33300 20812 33312
rect 19260 33272 20812 33300
rect 14277 33263 14335 33269
rect 20806 33260 20812 33272
rect 20864 33260 20870 33312
rect 20898 33260 20904 33312
rect 20956 33300 20962 33312
rect 25406 33300 25412 33312
rect 20956 33272 25412 33300
rect 20956 33260 20962 33272
rect 25406 33260 25412 33272
rect 25464 33260 25470 33312
rect 27614 33260 27620 33312
rect 27672 33300 27678 33312
rect 31021 33303 31079 33309
rect 31021 33300 31033 33303
rect 27672 33272 31033 33300
rect 27672 33260 27678 33272
rect 31021 33269 31033 33272
rect 31067 33269 31079 33303
rect 31021 33263 31079 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 3878 33056 3884 33108
rect 3936 33096 3942 33108
rect 8202 33096 8208 33108
rect 3936 33068 8208 33096
rect 3936 33056 3942 33068
rect 8202 33056 8208 33068
rect 8260 33056 8266 33108
rect 9214 33096 9220 33108
rect 9175 33068 9220 33096
rect 9214 33056 9220 33068
rect 9272 33056 9278 33108
rect 10318 33096 10324 33108
rect 10279 33068 10324 33096
rect 10318 33056 10324 33068
rect 10376 33056 10382 33108
rect 11514 33056 11520 33108
rect 11572 33096 11578 33108
rect 34054 33096 34060 33108
rect 11572 33068 34060 33096
rect 11572 33056 11578 33068
rect 34054 33056 34060 33068
rect 34112 33096 34118 33108
rect 34514 33096 34520 33108
rect 34112 33068 34520 33096
rect 34112 33056 34118 33068
rect 34514 33056 34520 33068
rect 34572 33056 34578 33108
rect 13814 33028 13820 33040
rect 13740 33000 13820 33028
rect 5074 32920 5080 32972
rect 5132 32960 5138 32972
rect 11440 32960 11652 32972
rect 13740 32969 13768 33000
rect 13814 32988 13820 33000
rect 13872 33028 13878 33040
rect 14090 33028 14096 33040
rect 13872 33000 14096 33028
rect 13872 32988 13878 33000
rect 14090 32988 14096 33000
rect 14148 32988 14154 33040
rect 14918 32988 14924 33040
rect 14976 33028 14982 33040
rect 20162 33028 20168 33040
rect 14976 33000 20168 33028
rect 14976 32988 14982 33000
rect 20162 32988 20168 33000
rect 20220 32988 20226 33040
rect 22094 32988 22100 33040
rect 22152 33028 22158 33040
rect 22557 33031 22615 33037
rect 22557 33028 22569 33031
rect 22152 33000 22569 33028
rect 22152 32988 22158 33000
rect 22557 32997 22569 33000
rect 22603 32997 22615 33031
rect 25038 33028 25044 33040
rect 24999 33000 25044 33028
rect 22557 32991 22615 32997
rect 25038 32988 25044 33000
rect 25096 32988 25102 33040
rect 13725 32963 13783 32969
rect 5132 32944 13676 32960
rect 5132 32932 11468 32944
rect 11624 32932 13676 32944
rect 5132 32920 5138 32932
rect 1578 32892 1584 32904
rect 1539 32864 1584 32892
rect 1578 32852 1584 32864
rect 1636 32852 1642 32904
rect 7377 32895 7435 32901
rect 7377 32861 7389 32895
rect 7423 32892 7435 32895
rect 8386 32892 8392 32904
rect 7423 32864 8392 32892
rect 7423 32861 7435 32864
rect 7377 32855 7435 32861
rect 8386 32852 8392 32864
rect 8444 32852 8450 32904
rect 9125 32895 9183 32901
rect 9125 32861 9137 32895
rect 9171 32861 9183 32895
rect 10226 32892 10232 32904
rect 10187 32864 10232 32892
rect 9125 32855 9183 32861
rect 1762 32756 1768 32768
rect 1723 32728 1768 32756
rect 1762 32716 1768 32728
rect 1820 32716 1826 32768
rect 7282 32716 7288 32768
rect 7340 32756 7346 32768
rect 7469 32759 7527 32765
rect 7469 32756 7481 32759
rect 7340 32728 7481 32756
rect 7340 32716 7346 32728
rect 7469 32725 7481 32728
rect 7515 32725 7527 32759
rect 9140 32756 9168 32855
rect 10226 32852 10232 32864
rect 10284 32852 10290 32904
rect 10870 32892 10876 32904
rect 10831 32864 10876 32892
rect 10870 32852 10876 32864
rect 10928 32852 10934 32904
rect 11514 32892 11520 32904
rect 11475 32864 11520 32892
rect 11514 32852 11520 32864
rect 11572 32852 11578 32904
rect 11609 32895 11667 32901
rect 11609 32861 11621 32895
rect 11655 32892 11667 32895
rect 12342 32892 12348 32904
rect 11655 32864 12348 32892
rect 11655 32861 11667 32864
rect 11609 32855 11667 32861
rect 12342 32852 12348 32864
rect 12400 32852 12406 32904
rect 10965 32827 11023 32833
rect 10965 32793 10977 32827
rect 11011 32824 11023 32827
rect 11011 32796 12480 32824
rect 11011 32793 11023 32796
rect 10965 32787 11023 32793
rect 11330 32756 11336 32768
rect 9140 32728 11336 32756
rect 7469 32719 7527 32725
rect 11330 32716 11336 32728
rect 11388 32756 11394 32768
rect 12342 32756 12348 32768
rect 11388 32728 12348 32756
rect 11388 32716 11394 32728
rect 12342 32716 12348 32728
rect 12400 32716 12406 32768
rect 12452 32756 12480 32796
rect 12526 32784 12532 32836
rect 12584 32824 12590 32836
rect 12713 32827 12771 32833
rect 12713 32824 12725 32827
rect 12584 32796 12725 32824
rect 12584 32784 12590 32796
rect 12713 32793 12725 32796
rect 12759 32793 12771 32827
rect 12713 32787 12771 32793
rect 12805 32827 12863 32833
rect 12805 32793 12817 32827
rect 12851 32824 12863 32827
rect 13354 32824 13360 32836
rect 12851 32796 13360 32824
rect 12851 32793 12863 32796
rect 12805 32787 12863 32793
rect 13354 32784 13360 32796
rect 13412 32784 13418 32836
rect 13648 32824 13676 32932
rect 13725 32929 13737 32963
rect 13771 32929 13783 32963
rect 13725 32923 13783 32929
rect 17494 32920 17500 32972
rect 17552 32960 17558 32972
rect 20254 32960 20260 32972
rect 17552 32932 20260 32960
rect 17552 32920 17558 32932
rect 20254 32920 20260 32932
rect 20312 32920 20318 32972
rect 20806 32960 20812 32972
rect 20767 32932 20812 32960
rect 20806 32920 20812 32932
rect 20864 32920 20870 32972
rect 25590 32920 25596 32972
rect 25648 32960 25654 32972
rect 25961 32963 26019 32969
rect 25961 32960 25973 32963
rect 25648 32932 25973 32960
rect 25648 32920 25654 32932
rect 25961 32929 25973 32932
rect 26007 32929 26019 32963
rect 25961 32923 26019 32929
rect 27525 32963 27583 32969
rect 27525 32929 27537 32963
rect 27571 32960 27583 32963
rect 27614 32960 27620 32972
rect 27571 32932 27620 32960
rect 27571 32929 27583 32932
rect 27525 32923 27583 32929
rect 27614 32920 27620 32932
rect 27672 32920 27678 32972
rect 28442 32960 28448 32972
rect 28403 32932 28448 32960
rect 28442 32920 28448 32932
rect 28500 32920 28506 32972
rect 14829 32895 14887 32901
rect 14829 32861 14841 32895
rect 14875 32894 14887 32895
rect 14875 32892 15056 32894
rect 16942 32892 16948 32904
rect 14875 32866 16948 32892
rect 14875 32861 14887 32866
rect 15028 32864 16948 32866
rect 14829 32855 14887 32861
rect 16942 32852 16948 32864
rect 17000 32852 17006 32904
rect 24578 32852 24584 32904
rect 24636 32892 24642 32904
rect 24949 32895 25007 32901
rect 24949 32892 24961 32895
rect 24636 32864 24961 32892
rect 24636 32852 24642 32864
rect 24949 32861 24961 32864
rect 24995 32861 25007 32895
rect 24949 32855 25007 32861
rect 27341 32895 27399 32901
rect 27341 32861 27353 32895
rect 27387 32861 27399 32895
rect 37458 32892 37464 32904
rect 37419 32864 37464 32892
rect 27341 32855 27399 32861
rect 13648 32796 15056 32824
rect 13078 32756 13084 32768
rect 12452 32728 13084 32756
rect 13078 32716 13084 32728
rect 13136 32716 13142 32768
rect 13170 32716 13176 32768
rect 13228 32756 13234 32768
rect 14921 32759 14979 32765
rect 14921 32756 14933 32759
rect 13228 32728 14933 32756
rect 13228 32716 13234 32728
rect 14921 32725 14933 32728
rect 14967 32725 14979 32759
rect 15028 32756 15056 32796
rect 17402 32784 17408 32836
rect 17460 32824 17466 32836
rect 21085 32827 21143 32833
rect 21085 32824 21097 32827
rect 17460 32796 21097 32824
rect 17460 32784 17466 32796
rect 21085 32793 21097 32796
rect 21131 32793 21143 32827
rect 21085 32787 21143 32793
rect 21542 32784 21548 32836
rect 21600 32784 21606 32836
rect 27356 32824 27384 32855
rect 37458 32852 37464 32864
rect 37516 32852 37522 32904
rect 37737 32895 37795 32901
rect 37737 32861 37749 32895
rect 37783 32892 37795 32895
rect 38746 32892 38752 32904
rect 37783 32864 38752 32892
rect 37783 32861 37795 32864
rect 37737 32855 37795 32861
rect 38746 32852 38752 32864
rect 38804 32852 38810 32904
rect 28350 32824 28356 32836
rect 27356 32796 28356 32824
rect 27356 32756 27384 32796
rect 28350 32784 28356 32796
rect 28408 32784 28414 32836
rect 28442 32784 28448 32836
rect 28500 32824 28506 32836
rect 37274 32824 37280 32836
rect 28500 32796 37280 32824
rect 28500 32784 28506 32796
rect 37274 32784 37280 32796
rect 37332 32784 37338 32836
rect 15028 32728 27384 32756
rect 14921 32719 14979 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 10321 32555 10379 32561
rect 10321 32521 10333 32555
rect 10367 32552 10379 32555
rect 10410 32552 10416 32564
rect 10367 32524 10416 32552
rect 10367 32521 10379 32524
rect 10321 32515 10379 32521
rect 10410 32512 10416 32524
rect 10468 32512 10474 32564
rect 11793 32555 11851 32561
rect 11793 32521 11805 32555
rect 11839 32552 11851 32555
rect 14918 32552 14924 32564
rect 11839 32524 14924 32552
rect 11839 32521 11851 32524
rect 11793 32515 11851 32521
rect 14918 32512 14924 32524
rect 14976 32512 14982 32564
rect 15194 32512 15200 32564
rect 15252 32552 15258 32564
rect 15252 32524 21312 32552
rect 15252 32512 15258 32524
rect 7282 32484 7288 32496
rect 7243 32456 7288 32484
rect 7282 32444 7288 32456
rect 7340 32444 7346 32496
rect 7837 32487 7895 32493
rect 7837 32453 7849 32487
rect 7883 32484 7895 32487
rect 10134 32484 10140 32496
rect 7883 32456 10140 32484
rect 7883 32453 7895 32456
rect 7837 32447 7895 32453
rect 10134 32444 10140 32456
rect 10192 32444 10198 32496
rect 12986 32484 12992 32496
rect 10244 32456 12992 32484
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32416 1639 32419
rect 2038 32416 2044 32428
rect 1627 32388 2044 32416
rect 1627 32385 1639 32388
rect 1581 32379 1639 32385
rect 2038 32376 2044 32388
rect 2096 32376 2102 32428
rect 10244 32425 10272 32456
rect 12986 32444 12992 32456
rect 13044 32444 13050 32496
rect 13078 32444 13084 32496
rect 13136 32484 13142 32496
rect 15838 32484 15844 32496
rect 13136 32456 15844 32484
rect 13136 32444 13142 32456
rect 15838 32444 15844 32456
rect 15896 32444 15902 32496
rect 17129 32487 17187 32493
rect 17129 32453 17141 32487
rect 17175 32484 17187 32487
rect 17218 32484 17224 32496
rect 17175 32456 17224 32484
rect 17175 32453 17187 32456
rect 17129 32447 17187 32453
rect 17218 32444 17224 32456
rect 17276 32444 17282 32496
rect 18414 32444 18420 32496
rect 18472 32484 18478 32496
rect 19981 32487 20039 32493
rect 19981 32484 19993 32487
rect 18472 32456 19993 32484
rect 18472 32444 18478 32456
rect 19981 32453 19993 32456
rect 20027 32453 20039 32487
rect 19981 32447 20039 32453
rect 10229 32419 10287 32425
rect 10229 32385 10241 32419
rect 10275 32385 10287 32419
rect 10229 32379 10287 32385
rect 10870 32376 10876 32428
rect 10928 32416 10934 32428
rect 11698 32416 11704 32428
rect 10928 32388 11704 32416
rect 10928 32376 10934 32388
rect 11698 32376 11704 32388
rect 11756 32376 11762 32428
rect 12250 32376 12256 32428
rect 12308 32416 12314 32428
rect 12345 32419 12403 32425
rect 12345 32416 12357 32419
rect 12308 32388 12357 32416
rect 12308 32376 12314 32388
rect 12345 32385 12357 32388
rect 12391 32385 12403 32419
rect 12345 32379 12403 32385
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32416 13691 32419
rect 14918 32416 14924 32428
rect 13679 32388 14924 32416
rect 13679 32385 13691 32388
rect 13633 32379 13691 32385
rect 14918 32376 14924 32388
rect 14976 32376 14982 32428
rect 16850 32416 16856 32428
rect 16684 32388 16856 32416
rect 7190 32348 7196 32360
rect 7151 32320 7196 32348
rect 7190 32308 7196 32320
rect 7248 32308 7254 32360
rect 14550 32348 14556 32360
rect 12636 32320 14556 32348
rect 10226 32240 10232 32292
rect 10284 32280 10290 32292
rect 12437 32283 12495 32289
rect 10284 32252 10732 32280
rect 10284 32240 10290 32252
rect 1762 32212 1768 32224
rect 1723 32184 1768 32212
rect 1762 32172 1768 32184
rect 1820 32172 1826 32224
rect 10134 32172 10140 32224
rect 10192 32212 10198 32224
rect 10594 32212 10600 32224
rect 10192 32184 10600 32212
rect 10192 32172 10198 32184
rect 10594 32172 10600 32184
rect 10652 32172 10658 32224
rect 10704 32212 10732 32252
rect 12437 32249 12449 32283
rect 12483 32280 12495 32283
rect 12636 32280 12664 32320
rect 14550 32308 14556 32320
rect 14608 32308 14614 32360
rect 15102 32308 15108 32360
rect 15160 32348 15166 32360
rect 16684 32348 16712 32388
rect 16850 32376 16856 32388
rect 16908 32376 16914 32428
rect 18230 32376 18236 32428
rect 18288 32376 18294 32428
rect 21082 32376 21088 32428
rect 21140 32376 21146 32428
rect 15160 32320 16712 32348
rect 16776 32320 18184 32348
rect 15160 32308 15166 32320
rect 12483 32252 12664 32280
rect 12483 32249 12495 32252
rect 12437 32243 12495 32249
rect 15378 32240 15384 32292
rect 15436 32280 15442 32292
rect 16776 32280 16804 32320
rect 15436 32252 16804 32280
rect 18156 32280 18184 32320
rect 19242 32308 19248 32360
rect 19300 32348 19306 32360
rect 19705 32351 19763 32357
rect 19705 32348 19717 32351
rect 19300 32320 19717 32348
rect 19300 32308 19306 32320
rect 19705 32317 19717 32320
rect 19751 32317 19763 32351
rect 19705 32311 19763 32317
rect 21284 32280 21312 32524
rect 21450 32512 21456 32564
rect 21508 32552 21514 32564
rect 28718 32552 28724 32564
rect 21508 32524 28724 32552
rect 21508 32512 21514 32524
rect 28718 32512 28724 32524
rect 28776 32512 28782 32564
rect 38102 32552 38108 32564
rect 38063 32524 38108 32552
rect 38102 32512 38108 32524
rect 38160 32512 38166 32564
rect 23106 32416 23112 32428
rect 23067 32388 23112 32416
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 26142 32376 26148 32428
rect 26200 32376 26206 32428
rect 38286 32416 38292 32428
rect 38247 32388 38292 32416
rect 38286 32376 38292 32388
rect 38344 32376 38350 32428
rect 21726 32308 21732 32360
rect 21784 32348 21790 32360
rect 22002 32348 22008 32360
rect 21784 32320 22008 32348
rect 21784 32308 21790 32320
rect 22002 32308 22008 32320
rect 22060 32348 22066 32360
rect 23845 32351 23903 32357
rect 23845 32348 23857 32351
rect 22060 32320 23857 32348
rect 22060 32308 22066 32320
rect 23845 32317 23857 32320
rect 23891 32348 23903 32351
rect 24765 32351 24823 32357
rect 24765 32348 24777 32351
rect 23891 32320 24777 32348
rect 23891 32317 23903 32320
rect 23845 32311 23903 32317
rect 24765 32317 24777 32320
rect 24811 32317 24823 32351
rect 24765 32311 24823 32317
rect 25041 32351 25099 32357
rect 25041 32317 25053 32351
rect 25087 32348 25099 32351
rect 26234 32348 26240 32360
rect 25087 32320 26240 32348
rect 25087 32317 25099 32320
rect 25041 32311 25099 32317
rect 26234 32308 26240 32320
rect 26292 32308 26298 32360
rect 22646 32280 22652 32292
rect 18156 32252 19334 32280
rect 21284 32252 22652 32280
rect 15436 32240 15442 32252
rect 13725 32215 13783 32221
rect 13725 32212 13737 32215
rect 10704 32184 13737 32212
rect 13725 32181 13737 32184
rect 13771 32181 13783 32215
rect 13725 32175 13783 32181
rect 15010 32172 15016 32224
rect 15068 32212 15074 32224
rect 16758 32212 16764 32224
rect 15068 32184 16764 32212
rect 15068 32172 15074 32184
rect 16758 32172 16764 32184
rect 16816 32172 16822 32224
rect 16850 32172 16856 32224
rect 16908 32212 16914 32224
rect 18506 32212 18512 32224
rect 16908 32184 18512 32212
rect 16908 32172 16914 32184
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 18598 32172 18604 32224
rect 18656 32212 18662 32224
rect 19306 32212 19334 32252
rect 22646 32240 22652 32252
rect 22704 32240 22710 32292
rect 21450 32212 21456 32224
rect 18656 32184 18701 32212
rect 19306 32184 21456 32212
rect 18656 32172 18662 32184
rect 21450 32172 21456 32184
rect 21508 32172 21514 32224
rect 26326 32172 26332 32224
rect 26384 32212 26390 32224
rect 26513 32215 26571 32221
rect 26513 32212 26525 32215
rect 26384 32184 26525 32212
rect 26384 32172 26390 32184
rect 26513 32181 26525 32184
rect 26559 32181 26571 32215
rect 26513 32175 26571 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 9217 32011 9275 32017
rect 9217 31977 9229 32011
rect 9263 32008 9275 32011
rect 12066 32008 12072 32020
rect 9263 31980 12072 32008
rect 9263 31977 9275 31980
rect 9217 31971 9275 31977
rect 12066 31968 12072 31980
rect 12124 32008 12130 32020
rect 12124 31980 12756 32008
rect 12124 31968 12130 31980
rect 11146 31872 11152 31884
rect 11107 31844 11152 31872
rect 11146 31832 11152 31844
rect 11204 31832 11210 31884
rect 12161 31875 12219 31881
rect 12161 31841 12173 31875
rect 12207 31872 12219 31875
rect 12526 31872 12532 31884
rect 12207 31844 12532 31872
rect 12207 31841 12219 31844
rect 12161 31835 12219 31841
rect 12526 31832 12532 31844
rect 12584 31832 12590 31884
rect 12728 31881 12756 31980
rect 21082 31968 21088 32020
rect 21140 32008 21146 32020
rect 24673 32011 24731 32017
rect 24673 32008 24685 32011
rect 21140 31980 24685 32008
rect 21140 31968 21146 31980
rect 24673 31977 24685 31980
rect 24719 31977 24731 32011
rect 24673 31971 24731 31977
rect 26973 32011 27031 32017
rect 26973 31977 26985 32011
rect 27019 32008 27031 32011
rect 27522 32008 27528 32020
rect 27019 31980 27528 32008
rect 27019 31977 27031 31980
rect 26973 31971 27031 31977
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 35894 31968 35900 32020
rect 35952 32008 35958 32020
rect 36173 32011 36231 32017
rect 36173 32008 36185 32011
rect 35952 31980 36185 32008
rect 35952 31968 35958 31980
rect 36173 31977 36185 31980
rect 36219 31977 36231 32011
rect 36173 31971 36231 31977
rect 12802 31900 12808 31952
rect 12860 31940 12866 31952
rect 15010 31940 15016 31952
rect 12860 31912 15016 31940
rect 12860 31900 12866 31912
rect 15010 31900 15016 31912
rect 15068 31900 15074 31952
rect 16666 31900 16672 31952
rect 16724 31940 16730 31952
rect 16853 31943 16911 31949
rect 16853 31940 16865 31943
rect 16724 31912 16865 31940
rect 16724 31900 16730 31912
rect 16853 31909 16865 31912
rect 16899 31940 16911 31943
rect 24026 31940 24032 31952
rect 16899 31912 19564 31940
rect 23987 31912 24032 31940
rect 16899 31909 16911 31912
rect 16853 31903 16911 31909
rect 12713 31875 12771 31881
rect 12713 31841 12725 31875
rect 12759 31841 12771 31875
rect 13354 31872 13360 31884
rect 13315 31844 13360 31872
rect 12713 31835 12771 31841
rect 13354 31832 13360 31844
rect 13412 31832 13418 31884
rect 15378 31872 15384 31884
rect 15291 31844 15384 31872
rect 15378 31832 15384 31844
rect 15436 31872 15442 31884
rect 17862 31872 17868 31884
rect 15436 31844 17868 31872
rect 15436 31832 15442 31844
rect 17862 31832 17868 31844
rect 17920 31832 17926 31884
rect 18506 31832 18512 31884
rect 18564 31872 18570 31884
rect 19242 31872 19248 31884
rect 18564 31844 19248 31872
rect 18564 31832 18570 31844
rect 19242 31832 19248 31844
rect 19300 31872 19306 31884
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 19300 31844 19441 31872
rect 19300 31832 19306 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 19536 31872 19564 31912
rect 24026 31900 24032 31912
rect 24084 31900 24090 31952
rect 33502 31900 33508 31952
rect 33560 31940 33566 31952
rect 34054 31940 34060 31952
rect 33560 31912 34060 31940
rect 33560 31900 33566 31912
rect 34054 31900 34060 31912
rect 34112 31900 34118 31952
rect 19705 31875 19763 31881
rect 19705 31872 19717 31875
rect 19536 31844 19717 31872
rect 19429 31835 19487 31841
rect 19705 31841 19717 31844
rect 19751 31841 19763 31875
rect 19705 31835 19763 31841
rect 20070 31832 20076 31884
rect 20128 31872 20134 31884
rect 21177 31875 21235 31881
rect 21177 31872 21189 31875
rect 20128 31844 21189 31872
rect 20128 31832 20134 31844
rect 21177 31841 21189 31844
rect 21223 31841 21235 31875
rect 21177 31835 21235 31841
rect 21634 31832 21640 31884
rect 21692 31872 21698 31884
rect 22557 31875 22615 31881
rect 22557 31872 22569 31875
rect 21692 31844 22569 31872
rect 21692 31832 21698 31844
rect 22557 31841 22569 31844
rect 22603 31841 22615 31875
rect 22557 31835 22615 31841
rect 22646 31832 22652 31884
rect 22704 31872 22710 31884
rect 28074 31872 28080 31884
rect 22704 31844 23796 31872
rect 22704 31832 22710 31844
rect 9122 31804 9128 31816
rect 9083 31776 9128 31804
rect 9122 31764 9128 31776
rect 9180 31764 9186 31816
rect 9766 31804 9772 31816
rect 9727 31776 9772 31804
rect 9766 31764 9772 31776
rect 9824 31764 9830 31816
rect 9858 31764 9864 31816
rect 9916 31804 9922 31816
rect 15102 31804 15108 31816
rect 9916 31776 9961 31804
rect 15063 31776 15108 31804
rect 9916 31764 9922 31776
rect 15102 31764 15108 31776
rect 15160 31764 15166 31816
rect 16758 31764 16764 31816
rect 16816 31804 16822 31816
rect 17402 31804 17408 31816
rect 16816 31776 17408 31804
rect 16816 31764 16822 31776
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 21082 31764 21088 31816
rect 21140 31804 21146 31816
rect 21140 31776 21772 31804
rect 21140 31764 21146 31776
rect 11238 31736 11244 31748
rect 11199 31708 11244 31736
rect 11238 31696 11244 31708
rect 11296 31696 11302 31748
rect 12802 31736 12808 31748
rect 12763 31708 12808 31736
rect 12802 31696 12808 31708
rect 12860 31696 12866 31748
rect 15838 31696 15844 31748
rect 15896 31696 15902 31748
rect 20162 31696 20168 31748
rect 20220 31696 20226 31748
rect 21744 31736 21772 31776
rect 22002 31764 22008 31816
rect 22060 31804 22066 31816
rect 22281 31807 22339 31813
rect 22281 31804 22293 31807
rect 22060 31776 22293 31804
rect 22060 31764 22066 31776
rect 22281 31773 22293 31776
rect 22327 31773 22339 31807
rect 23768 31804 23796 31844
rect 27540 31844 28080 31872
rect 24581 31807 24639 31813
rect 24581 31804 24593 31807
rect 23768 31776 24593 31804
rect 22281 31767 22339 31773
rect 24581 31773 24593 31776
rect 24627 31773 24639 31807
rect 24581 31767 24639 31773
rect 24946 31764 24952 31816
rect 25004 31804 25010 31816
rect 27540 31813 27568 31844
rect 28074 31832 28080 31844
rect 28132 31832 28138 31884
rect 32306 31872 32312 31884
rect 32267 31844 32312 31872
rect 32306 31832 32312 31844
rect 32364 31872 32370 31884
rect 35526 31872 35532 31884
rect 32364 31844 35532 31872
rect 32364 31832 32370 31844
rect 35526 31832 35532 31844
rect 35584 31832 35590 31884
rect 26881 31807 26939 31813
rect 26881 31804 26893 31807
rect 25004 31776 26893 31804
rect 25004 31764 25010 31776
rect 26881 31773 26893 31776
rect 26927 31773 26939 31807
rect 26881 31767 26939 31773
rect 27525 31807 27583 31813
rect 27525 31773 27537 31807
rect 27571 31773 27583 31807
rect 27525 31767 27583 31773
rect 27617 31807 27675 31813
rect 27617 31773 27629 31807
rect 27663 31804 27675 31807
rect 27706 31804 27712 31816
rect 27663 31776 27712 31804
rect 27663 31773 27675 31776
rect 27617 31767 27675 31773
rect 27706 31764 27712 31776
rect 27764 31764 27770 31816
rect 30374 31764 30380 31816
rect 30432 31804 30438 31816
rect 32033 31807 32091 31813
rect 32033 31804 32045 31807
rect 30432 31776 32045 31804
rect 30432 31764 30438 31776
rect 32033 31773 32045 31776
rect 32079 31773 32091 31807
rect 33594 31804 33600 31816
rect 33442 31776 33600 31804
rect 32033 31767 32091 31773
rect 33594 31764 33600 31776
rect 33652 31764 33658 31816
rect 34054 31804 34060 31816
rect 34015 31776 34060 31804
rect 34054 31764 34060 31776
rect 34112 31764 34118 31816
rect 36078 31804 36084 31816
rect 36039 31776 36084 31804
rect 36078 31764 36084 31776
rect 36136 31764 36142 31816
rect 21744 31708 23046 31736
rect 9398 31628 9404 31680
rect 9456 31668 9462 31680
rect 22462 31668 22468 31680
rect 9456 31640 22468 31668
rect 9456 31628 9462 31640
rect 22462 31628 22468 31640
rect 22520 31668 22526 31680
rect 23842 31668 23848 31680
rect 22520 31640 23848 31668
rect 22520 31628 22526 31640
rect 23842 31628 23848 31640
rect 23900 31628 23906 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 4249 31467 4307 31473
rect 4249 31433 4261 31467
rect 4295 31464 4307 31467
rect 4614 31464 4620 31476
rect 4295 31436 4620 31464
rect 4295 31433 4307 31436
rect 4249 31427 4307 31433
rect 4614 31424 4620 31436
rect 4672 31424 4678 31476
rect 6641 31467 6699 31473
rect 6641 31433 6653 31467
rect 6687 31464 6699 31467
rect 7190 31464 7196 31476
rect 6687 31436 7196 31464
rect 6687 31433 6699 31436
rect 6641 31427 6699 31433
rect 7190 31424 7196 31436
rect 7248 31464 7254 31476
rect 11793 31467 11851 31473
rect 7248 31436 8156 31464
rect 7248 31424 7254 31436
rect 8128 31405 8156 31436
rect 11793 31433 11805 31467
rect 11839 31464 11851 31467
rect 12802 31464 12808 31476
rect 11839 31436 12808 31464
rect 11839 31433 11851 31436
rect 11793 31427 11851 31433
rect 12802 31424 12808 31436
rect 12860 31424 12866 31476
rect 23934 31464 23940 31476
rect 15028 31436 23940 31464
rect 8113 31399 8171 31405
rect 8113 31365 8125 31399
rect 8159 31365 8171 31399
rect 8113 31359 8171 31365
rect 8205 31399 8263 31405
rect 8205 31365 8217 31399
rect 8251 31396 8263 31399
rect 9953 31399 10011 31405
rect 9953 31396 9965 31399
rect 8251 31368 9965 31396
rect 8251 31365 8263 31368
rect 8205 31359 8263 31365
rect 9953 31365 9965 31368
rect 9999 31365 10011 31399
rect 11054 31396 11060 31408
rect 9953 31359 10011 31365
rect 10428 31368 11060 31396
rect 4157 31331 4215 31337
rect 4157 31297 4169 31331
rect 4203 31328 4215 31331
rect 5258 31328 5264 31340
rect 4203 31300 5264 31328
rect 4203 31297 4215 31300
rect 4157 31291 4215 31297
rect 5258 31288 5264 31300
rect 5316 31288 5322 31340
rect 6549 31331 6607 31337
rect 6549 31297 6561 31331
rect 6595 31328 6607 31331
rect 6638 31328 6644 31340
rect 6595 31300 6644 31328
rect 6595 31297 6607 31300
rect 6549 31291 6607 31297
rect 6638 31288 6644 31300
rect 6696 31288 6702 31340
rect 9217 31331 9275 31337
rect 9217 31297 9229 31331
rect 9263 31297 9275 31331
rect 9217 31291 9275 31297
rect 9861 31331 9919 31337
rect 9861 31297 9873 31331
rect 9907 31328 9919 31331
rect 10428 31328 10456 31368
rect 11054 31356 11060 31368
rect 11112 31356 11118 31408
rect 13357 31399 13415 31405
rect 13357 31365 13369 31399
rect 13403 31396 13415 31399
rect 13403 31368 14412 31396
rect 13403 31365 13415 31368
rect 13357 31359 13415 31365
rect 9907 31300 10456 31328
rect 10505 31331 10563 31337
rect 9907 31297 9919 31300
rect 9861 31291 9919 31297
rect 10505 31297 10517 31331
rect 10551 31297 10563 31331
rect 11698 31328 11704 31340
rect 11659 31300 11704 31328
rect 10505 31291 10563 31297
rect 6362 31220 6368 31272
rect 6420 31260 6426 31272
rect 9232 31260 9260 31291
rect 6420 31232 9260 31260
rect 6420 31220 6426 31232
rect 8665 31195 8723 31201
rect 8665 31161 8677 31195
rect 8711 31192 8723 31195
rect 10410 31192 10416 31204
rect 8711 31164 10416 31192
rect 8711 31161 8723 31164
rect 8665 31155 8723 31161
rect 10410 31152 10416 31164
rect 10468 31152 10474 31204
rect 10520 31192 10548 31291
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 12434 31220 12440 31272
rect 12492 31260 12498 31272
rect 13265 31263 13323 31269
rect 13265 31260 13277 31263
rect 12492 31232 13277 31260
rect 12492 31220 12498 31232
rect 13265 31229 13277 31232
rect 13311 31229 13323 31263
rect 14090 31260 14096 31272
rect 14051 31232 14096 31260
rect 13265 31223 13323 31229
rect 14090 31220 14096 31232
rect 14148 31220 14154 31272
rect 14384 31260 14412 31368
rect 15028 31337 15056 31436
rect 23934 31424 23940 31436
rect 23992 31424 23998 31476
rect 32582 31424 32588 31476
rect 32640 31464 32646 31476
rect 35802 31464 35808 31476
rect 32640 31436 35808 31464
rect 32640 31424 32646 31436
rect 35802 31424 35808 31436
rect 35860 31424 35866 31476
rect 20530 31396 20536 31408
rect 20102 31368 20536 31396
rect 20530 31356 20536 31368
rect 20588 31356 20594 31408
rect 25406 31356 25412 31408
rect 25464 31396 25470 31408
rect 33410 31396 33416 31408
rect 25464 31368 33416 31396
rect 25464 31356 25470 31368
rect 33410 31356 33416 31368
rect 33468 31356 33474 31408
rect 37366 31396 37372 31408
rect 35006 31368 37372 31396
rect 37366 31356 37372 31368
rect 37424 31356 37430 31408
rect 15013 31331 15071 31337
rect 15013 31297 15025 31331
rect 15059 31297 15071 31331
rect 15013 31291 15071 31297
rect 18506 31288 18512 31340
rect 18564 31328 18570 31340
rect 18601 31331 18659 31337
rect 18601 31328 18613 31331
rect 18564 31300 18613 31328
rect 18564 31288 18570 31300
rect 18601 31297 18613 31300
rect 18647 31297 18659 31331
rect 18601 31291 18659 31297
rect 35713 31331 35771 31337
rect 35713 31297 35725 31331
rect 35759 31328 35771 31331
rect 35802 31328 35808 31340
rect 35759 31300 35808 31328
rect 35759 31297 35771 31300
rect 35713 31291 35771 31297
rect 35802 31288 35808 31300
rect 35860 31288 35866 31340
rect 15105 31263 15163 31269
rect 15105 31260 15117 31263
rect 14384 31232 15117 31260
rect 15105 31229 15117 31232
rect 15151 31229 15163 31263
rect 15105 31223 15163 31229
rect 18877 31263 18935 31269
rect 18877 31229 18889 31263
rect 18923 31260 18935 31263
rect 19242 31260 19248 31272
rect 18923 31232 19248 31260
rect 18923 31229 18935 31232
rect 18877 31223 18935 31229
rect 19242 31220 19248 31232
rect 19300 31220 19306 31272
rect 32214 31220 32220 31272
rect 32272 31260 32278 31272
rect 33505 31263 33563 31269
rect 33505 31260 33517 31263
rect 32272 31232 33517 31260
rect 32272 31220 32278 31232
rect 33505 31229 33517 31232
rect 33551 31229 33563 31263
rect 33505 31223 33563 31229
rect 33781 31263 33839 31269
rect 33781 31229 33793 31263
rect 33827 31260 33839 31263
rect 36630 31260 36636 31272
rect 33827 31232 36636 31260
rect 33827 31229 33839 31232
rect 33781 31223 33839 31229
rect 36630 31220 36636 31232
rect 36688 31220 36694 31272
rect 10520 31164 12434 31192
rect 9309 31127 9367 31133
rect 9309 31093 9321 31127
rect 9355 31124 9367 31127
rect 9674 31124 9680 31136
rect 9355 31096 9680 31124
rect 9355 31093 9367 31096
rect 9309 31087 9367 31093
rect 9674 31084 9680 31096
rect 9732 31084 9738 31136
rect 10597 31127 10655 31133
rect 10597 31093 10609 31127
rect 10643 31124 10655 31127
rect 10778 31124 10784 31136
rect 10643 31096 10784 31124
rect 10643 31093 10655 31096
rect 10597 31087 10655 31093
rect 10778 31084 10784 31096
rect 10836 31084 10842 31136
rect 12406 31124 12434 31164
rect 14550 31152 14556 31204
rect 14608 31192 14614 31204
rect 16114 31192 16120 31204
rect 14608 31164 16120 31192
rect 14608 31152 14614 31164
rect 16114 31152 16120 31164
rect 16172 31152 16178 31204
rect 20162 31124 20168 31136
rect 12406 31096 20168 31124
rect 20162 31084 20168 31096
rect 20220 31084 20226 31136
rect 20349 31127 20407 31133
rect 20349 31093 20361 31127
rect 20395 31124 20407 31127
rect 27430 31124 27436 31136
rect 20395 31096 27436 31124
rect 20395 31093 20407 31096
rect 20349 31087 20407 31093
rect 27430 31084 27436 31096
rect 27488 31084 27494 31136
rect 35253 31127 35311 31133
rect 35253 31093 35265 31127
rect 35299 31124 35311 31127
rect 35526 31124 35532 31136
rect 35299 31096 35532 31124
rect 35299 31093 35311 31096
rect 35253 31087 35311 31093
rect 35526 31084 35532 31096
rect 35584 31084 35590 31136
rect 35805 31127 35863 31133
rect 35805 31093 35817 31127
rect 35851 31124 35863 31127
rect 36446 31124 36452 31136
rect 35851 31096 36452 31124
rect 35851 31093 35863 31096
rect 35805 31087 35863 31093
rect 36446 31084 36452 31096
rect 36504 31084 36510 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 8386 30880 8392 30932
rect 8444 30920 8450 30932
rect 8444 30892 10640 30920
rect 8444 30880 8450 30892
rect 10226 30852 10232 30864
rect 9508 30824 10232 30852
rect 9508 30793 9536 30824
rect 10226 30812 10232 30824
rect 10284 30812 10290 30864
rect 10612 30852 10640 30892
rect 11698 30880 11704 30932
rect 11756 30920 11762 30932
rect 24670 30920 24676 30932
rect 11756 30892 24676 30920
rect 11756 30880 11762 30892
rect 24670 30880 24676 30892
rect 24728 30880 24734 30932
rect 24844 30923 24902 30929
rect 24844 30889 24856 30923
rect 24890 30920 24902 30923
rect 26694 30920 26700 30932
rect 24890 30892 26700 30920
rect 24890 30889 24902 30892
rect 24844 30883 24902 30889
rect 26694 30880 26700 30892
rect 26752 30880 26758 30932
rect 31008 30923 31066 30929
rect 31008 30889 31020 30923
rect 31054 30920 31066 30923
rect 34238 30920 34244 30932
rect 31054 30892 34244 30920
rect 31054 30889 31066 30892
rect 31008 30883 31066 30889
rect 34238 30880 34244 30892
rect 34296 30880 34302 30932
rect 14277 30855 14335 30861
rect 10612 30824 14228 30852
rect 9493 30787 9551 30793
rect 9493 30753 9505 30787
rect 9539 30753 9551 30787
rect 9493 30747 9551 30753
rect 9582 30744 9588 30796
rect 9640 30784 9646 30796
rect 10689 30787 10747 30793
rect 10689 30784 10701 30787
rect 9640 30756 10701 30784
rect 9640 30744 9646 30756
rect 10689 30753 10701 30756
rect 10735 30753 10747 30787
rect 10689 30747 10747 30753
rect 11701 30787 11759 30793
rect 11701 30753 11713 30787
rect 11747 30784 11759 30787
rect 13262 30784 13268 30796
rect 11747 30756 13268 30784
rect 11747 30753 11759 30756
rect 11701 30747 11759 30753
rect 13262 30744 13268 30756
rect 13320 30744 13326 30796
rect 13446 30784 13452 30796
rect 13407 30756 13452 30784
rect 13446 30744 13452 30756
rect 13504 30744 13510 30796
rect 14200 30784 14228 30824
rect 14277 30821 14289 30855
rect 14323 30852 14335 30855
rect 14323 30824 15332 30852
rect 14323 30821 14335 30824
rect 14277 30815 14335 30821
rect 14200 30756 15056 30784
rect 1581 30719 1639 30725
rect 1581 30685 1593 30719
rect 1627 30716 1639 30719
rect 4706 30716 4712 30728
rect 1627 30688 4712 30716
rect 1627 30685 1639 30688
rect 1581 30679 1639 30685
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 12158 30716 12164 30728
rect 12119 30688 12164 30716
rect 12158 30676 12164 30688
rect 12216 30676 12222 30728
rect 14458 30716 14464 30728
rect 14419 30688 14464 30716
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 9582 30608 9588 30660
rect 9640 30648 9646 30660
rect 10137 30651 10195 30657
rect 9640 30620 9685 30648
rect 9640 30608 9646 30620
rect 10137 30617 10149 30651
rect 10183 30617 10195 30651
rect 10137 30611 10195 30617
rect 1762 30580 1768 30592
rect 1723 30552 1768 30580
rect 1762 30540 1768 30552
rect 1820 30540 1826 30592
rect 10152 30580 10180 30611
rect 10778 30608 10784 30660
rect 10836 30648 10842 30660
rect 13081 30651 13139 30657
rect 10836 30620 10881 30648
rect 10836 30608 10842 30620
rect 13081 30617 13093 30651
rect 13127 30617 13139 30651
rect 13081 30611 13139 30617
rect 13173 30651 13231 30657
rect 13173 30617 13185 30651
rect 13219 30648 13231 30651
rect 14826 30648 14832 30660
rect 13219 30620 14832 30648
rect 13219 30617 13231 30620
rect 13173 30611 13231 30617
rect 10594 30580 10600 30592
rect 10152 30552 10600 30580
rect 10594 30540 10600 30552
rect 10652 30540 10658 30592
rect 12253 30583 12311 30589
rect 12253 30549 12265 30583
rect 12299 30580 12311 30583
rect 12802 30580 12808 30592
rect 12299 30552 12808 30580
rect 12299 30549 12311 30552
rect 12253 30543 12311 30549
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 12986 30540 12992 30592
rect 13044 30580 13050 30592
rect 13096 30580 13124 30611
rect 14826 30608 14832 30620
rect 14884 30608 14890 30660
rect 15028 30648 15056 30756
rect 15102 30744 15108 30796
rect 15160 30784 15166 30796
rect 15197 30787 15255 30793
rect 15197 30784 15209 30787
rect 15160 30756 15209 30784
rect 15160 30744 15166 30756
rect 15197 30753 15209 30756
rect 15243 30753 15255 30787
rect 15304 30784 15332 30824
rect 15562 30784 15568 30796
rect 15304 30756 15568 30784
rect 15197 30747 15255 30753
rect 15562 30744 15568 30756
rect 15620 30744 15626 30796
rect 16758 30744 16764 30796
rect 16816 30784 16822 30796
rect 17221 30787 17279 30793
rect 17221 30784 17233 30787
rect 16816 30756 17233 30784
rect 16816 30744 16822 30756
rect 17221 30753 17233 30756
rect 17267 30753 17279 30787
rect 17221 30747 17279 30753
rect 18506 30744 18512 30796
rect 18564 30784 18570 30796
rect 18693 30787 18751 30793
rect 18693 30784 18705 30787
rect 18564 30756 18705 30784
rect 18564 30744 18570 30756
rect 18693 30753 18705 30756
rect 18739 30753 18751 30787
rect 18693 30747 18751 30753
rect 19613 30787 19671 30793
rect 19613 30753 19625 30787
rect 19659 30784 19671 30787
rect 21818 30784 21824 30796
rect 19659 30756 21824 30784
rect 19659 30753 19671 30756
rect 19613 30747 19671 30753
rect 21818 30744 21824 30756
rect 21876 30744 21882 30796
rect 23842 30784 23848 30796
rect 23803 30756 23848 30784
rect 23842 30744 23848 30756
rect 23900 30744 23906 30796
rect 24581 30787 24639 30793
rect 24581 30753 24593 30787
rect 24627 30784 24639 30787
rect 26142 30784 26148 30796
rect 24627 30756 26148 30784
rect 24627 30753 24639 30756
rect 24581 30747 24639 30753
rect 26142 30744 26148 30756
rect 26200 30744 26206 30796
rect 30745 30787 30803 30793
rect 30745 30753 30757 30787
rect 30791 30784 30803 30787
rect 32214 30784 32220 30796
rect 30791 30756 32220 30784
rect 30791 30753 30803 30756
rect 30745 30747 30803 30753
rect 32214 30744 32220 30756
rect 32272 30784 32278 30796
rect 34149 30787 34207 30793
rect 34149 30784 34161 30787
rect 32272 30756 34161 30784
rect 32272 30744 32278 30756
rect 34149 30753 34161 30756
rect 34195 30753 34207 30787
rect 34149 30747 34207 30753
rect 35894 30744 35900 30796
rect 35952 30784 35958 30796
rect 36265 30787 36323 30793
rect 36265 30784 36277 30787
rect 35952 30756 36277 30784
rect 35952 30744 35958 30756
rect 36265 30753 36277 30756
rect 36311 30753 36323 30787
rect 36446 30784 36452 30796
rect 36407 30756 36452 30784
rect 36265 30747 36323 30753
rect 36446 30744 36452 30756
rect 36504 30744 36510 30796
rect 37274 30784 37280 30796
rect 37235 30756 37280 30784
rect 37274 30744 37280 30756
rect 37332 30744 37338 30796
rect 16850 30676 16856 30728
rect 16908 30716 16914 30728
rect 17957 30719 18015 30725
rect 17957 30716 17969 30719
rect 16908 30688 17969 30716
rect 16908 30676 16914 30688
rect 17957 30685 17969 30688
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 32950 30676 32956 30728
rect 33008 30716 33014 30728
rect 33413 30719 33471 30725
rect 33413 30716 33425 30719
rect 33008 30688 33425 30716
rect 33008 30676 33014 30688
rect 33413 30685 33425 30688
rect 33459 30685 33471 30719
rect 33413 30679 33471 30685
rect 15473 30651 15531 30657
rect 15473 30648 15485 30651
rect 15028 30620 15485 30648
rect 15473 30617 15485 30620
rect 15519 30617 15531 30651
rect 15473 30611 15531 30617
rect 13044 30552 13124 30580
rect 15488 30580 15516 30611
rect 15746 30608 15752 30660
rect 15804 30648 15810 30660
rect 19889 30651 19947 30657
rect 15804 30620 15962 30648
rect 15804 30608 15810 30620
rect 19889 30617 19901 30651
rect 19935 30648 19947 30651
rect 19978 30648 19984 30660
rect 19935 30620 19984 30648
rect 19935 30617 19947 30620
rect 19889 30611 19947 30617
rect 19978 30608 19984 30620
rect 20036 30608 20042 30660
rect 20088 30620 20378 30648
rect 17402 30580 17408 30592
rect 15488 30552 17408 30580
rect 13044 30540 13050 30552
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 17862 30540 17868 30592
rect 17920 30580 17926 30592
rect 20088 30580 20116 30620
rect 21450 30608 21456 30660
rect 21508 30648 21514 30660
rect 22097 30651 22155 30657
rect 22097 30648 22109 30651
rect 21508 30620 22109 30648
rect 21508 30608 21514 30620
rect 22097 30617 22109 30620
rect 22143 30617 22155 30651
rect 26605 30651 26663 30657
rect 22097 30611 22155 30617
rect 22296 30620 22586 30648
rect 25240 30620 25346 30648
rect 17920 30552 20116 30580
rect 17920 30540 17926 30552
rect 20898 30540 20904 30592
rect 20956 30580 20962 30592
rect 21266 30580 21272 30592
rect 20956 30552 21272 30580
rect 20956 30540 20962 30552
rect 21266 30540 21272 30552
rect 21324 30580 21330 30592
rect 21361 30583 21419 30589
rect 21361 30580 21373 30583
rect 21324 30552 21373 30580
rect 21324 30540 21330 30552
rect 21361 30549 21373 30552
rect 21407 30549 21419 30583
rect 21361 30543 21419 30549
rect 21910 30540 21916 30592
rect 21968 30580 21974 30592
rect 22296 30580 22324 30620
rect 25240 30592 25268 30620
rect 26605 30617 26617 30651
rect 26651 30617 26663 30651
rect 26605 30611 26663 30617
rect 21968 30552 22324 30580
rect 21968 30540 21974 30552
rect 25222 30540 25228 30592
rect 25280 30540 25286 30592
rect 25866 30540 25872 30592
rect 25924 30580 25930 30592
rect 26234 30580 26240 30592
rect 25924 30552 26240 30580
rect 25924 30540 25930 30552
rect 26234 30540 26240 30552
rect 26292 30580 26298 30592
rect 26620 30580 26648 30611
rect 28626 30608 28632 30660
rect 28684 30648 28690 30660
rect 32766 30648 32772 30660
rect 28684 30620 31510 30648
rect 32727 30620 32772 30648
rect 28684 30608 28690 30620
rect 32766 30608 32772 30620
rect 32824 30608 32830 30660
rect 26292 30552 26648 30580
rect 26292 30540 26298 30552
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 8386 30336 8392 30388
rect 8444 30376 8450 30388
rect 8662 30376 8668 30388
rect 8444 30348 8668 30376
rect 8444 30336 8450 30348
rect 8662 30336 8668 30348
rect 8720 30336 8726 30388
rect 9217 30379 9275 30385
rect 9217 30345 9229 30379
rect 9263 30376 9275 30379
rect 9582 30376 9588 30388
rect 9263 30348 9588 30376
rect 9263 30345 9275 30348
rect 9217 30339 9275 30345
rect 9582 30336 9588 30348
rect 9640 30336 9646 30388
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 16574 30376 16580 30388
rect 12860 30348 16580 30376
rect 12860 30336 12866 30348
rect 16574 30336 16580 30348
rect 16632 30336 16638 30388
rect 24670 30336 24676 30388
rect 24728 30376 24734 30388
rect 29638 30376 29644 30388
rect 24728 30348 29644 30376
rect 24728 30336 24734 30348
rect 29638 30336 29644 30348
rect 29696 30336 29702 30388
rect 10226 30268 10232 30320
rect 10284 30308 10290 30320
rect 10494 30311 10552 30317
rect 10494 30308 10506 30311
rect 10284 30280 10506 30308
rect 10284 30268 10290 30280
rect 10494 30277 10506 30280
rect 10540 30277 10552 30311
rect 10494 30271 10552 30277
rect 10597 30311 10655 30317
rect 10597 30277 10609 30311
rect 10643 30308 10655 30311
rect 11514 30308 11520 30320
rect 10643 30280 11520 30308
rect 10643 30277 10655 30280
rect 10597 30271 10655 30277
rect 11514 30268 11520 30280
rect 11572 30268 11578 30320
rect 11885 30311 11943 30317
rect 11885 30277 11897 30311
rect 11931 30308 11943 30311
rect 13449 30311 13507 30317
rect 13449 30308 13461 30311
rect 11931 30280 13461 30308
rect 11931 30277 11943 30280
rect 11885 30271 11943 30277
rect 13449 30277 13461 30280
rect 13495 30277 13507 30311
rect 15102 30308 15108 30320
rect 13449 30271 13507 30277
rect 14568 30280 15108 30308
rect 8202 30200 8208 30252
rect 8260 30240 8266 30252
rect 9122 30240 9128 30252
rect 8260 30212 9128 30240
rect 8260 30200 8266 30212
rect 9122 30200 9128 30212
rect 9180 30200 9186 30252
rect 9766 30240 9772 30252
rect 9727 30212 9772 30240
rect 9766 30200 9772 30212
rect 9824 30200 9830 30252
rect 13357 30243 13415 30249
rect 13357 30209 13369 30243
rect 13403 30240 13415 30243
rect 14366 30240 14372 30252
rect 13403 30212 14372 30240
rect 13403 30209 13415 30212
rect 13357 30203 13415 30209
rect 14366 30200 14372 30212
rect 14424 30200 14430 30252
rect 14568 30249 14596 30280
rect 15102 30268 15108 30280
rect 15160 30268 15166 30320
rect 15286 30268 15292 30320
rect 15344 30268 15350 30320
rect 16114 30268 16120 30320
rect 16172 30308 16178 30320
rect 16172 30280 19458 30308
rect 16172 30268 16178 30280
rect 36262 30268 36268 30320
rect 36320 30268 36326 30320
rect 14553 30243 14611 30249
rect 14553 30209 14565 30243
rect 14599 30209 14611 30243
rect 14553 30203 14611 30209
rect 18506 30200 18512 30252
rect 18564 30240 18570 30252
rect 18693 30243 18751 30249
rect 18693 30240 18705 30243
rect 18564 30212 18705 30240
rect 18564 30200 18570 30212
rect 18693 30209 18705 30212
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 23106 30200 23112 30252
rect 23164 30240 23170 30252
rect 27614 30240 27620 30252
rect 23164 30212 27620 30240
rect 23164 30200 23170 30212
rect 27614 30200 27620 30212
rect 27672 30240 27678 30252
rect 29089 30243 29147 30249
rect 29089 30240 29101 30243
rect 27672 30212 29101 30240
rect 27672 30200 27678 30212
rect 29089 30209 29101 30212
rect 29135 30240 29147 30243
rect 30006 30240 30012 30252
rect 29135 30212 30012 30240
rect 29135 30209 29147 30212
rect 29089 30203 29147 30209
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 38286 30240 38292 30252
rect 38247 30212 38292 30240
rect 38286 30200 38292 30212
rect 38344 30200 38350 30252
rect 9861 30175 9919 30181
rect 9861 30141 9873 30175
rect 9907 30172 9919 30175
rect 11790 30172 11796 30184
rect 9907 30144 11376 30172
rect 11751 30144 11796 30172
rect 9907 30141 9919 30144
rect 9861 30135 9919 30141
rect 10410 30064 10416 30116
rect 10468 30104 10474 30116
rect 11057 30107 11115 30113
rect 11057 30104 11069 30107
rect 10468 30076 11069 30104
rect 10468 30064 10474 30076
rect 11057 30073 11069 30076
rect 11103 30073 11115 30107
rect 11348 30104 11376 30144
rect 11790 30132 11796 30144
rect 11848 30132 11854 30184
rect 12437 30175 12495 30181
rect 12437 30141 12449 30175
rect 12483 30172 12495 30175
rect 13906 30172 13912 30184
rect 12483 30144 13912 30172
rect 12483 30141 12495 30144
rect 12437 30135 12495 30141
rect 13906 30132 13912 30144
rect 13964 30132 13970 30184
rect 14829 30175 14887 30181
rect 14829 30172 14841 30175
rect 14660 30144 14841 30172
rect 12250 30104 12256 30116
rect 11348 30076 12256 30104
rect 11057 30067 11115 30073
rect 12250 30064 12256 30076
rect 12308 30064 12314 30116
rect 14274 30064 14280 30116
rect 14332 30104 14338 30116
rect 14660 30104 14688 30144
rect 14829 30141 14841 30144
rect 14875 30172 14887 30175
rect 18598 30172 18604 30184
rect 14875 30144 18604 30172
rect 14875 30141 14887 30144
rect 14829 30135 14887 30141
rect 18598 30132 18604 30144
rect 18656 30132 18662 30184
rect 18969 30175 19027 30181
rect 18969 30172 18981 30175
rect 18708 30144 18981 30172
rect 14332 30076 14688 30104
rect 14332 30064 14338 30076
rect 16022 30064 16028 30116
rect 16080 30104 16086 30116
rect 16758 30104 16764 30116
rect 16080 30076 16764 30104
rect 16080 30064 16086 30076
rect 16758 30064 16764 30076
rect 16816 30064 16822 30116
rect 18322 30064 18328 30116
rect 18380 30104 18386 30116
rect 18708 30104 18736 30144
rect 18969 30141 18981 30144
rect 19015 30172 19027 30175
rect 19058 30172 19064 30184
rect 19015 30144 19064 30172
rect 19015 30141 19027 30144
rect 18969 30135 19027 30141
rect 19058 30132 19064 30144
rect 19116 30132 19122 30184
rect 29730 30132 29736 30184
rect 29788 30172 29794 30184
rect 29825 30175 29883 30181
rect 29825 30172 29837 30175
rect 29788 30144 29837 30172
rect 29788 30132 29794 30144
rect 29825 30141 29837 30144
rect 29871 30172 29883 30175
rect 30374 30172 30380 30184
rect 29871 30144 30380 30172
rect 29871 30141 29883 30144
rect 29825 30135 29883 30141
rect 30374 30132 30380 30144
rect 30432 30132 30438 30184
rect 34790 30132 34796 30184
rect 34848 30172 34854 30184
rect 34977 30175 35035 30181
rect 34977 30172 34989 30175
rect 34848 30144 34989 30172
rect 34848 30132 34854 30144
rect 34977 30141 34989 30144
rect 35023 30141 35035 30175
rect 35250 30172 35256 30184
rect 35211 30144 35256 30172
rect 34977 30135 35035 30141
rect 35250 30132 35256 30144
rect 35308 30132 35314 30184
rect 37550 30104 37556 30116
rect 18380 30076 18736 30104
rect 36280 30076 37556 30104
rect 18380 30064 18386 30076
rect 10870 29996 10876 30048
rect 10928 30036 10934 30048
rect 12158 30036 12164 30048
rect 10928 30008 12164 30036
rect 10928 29996 10934 30008
rect 12158 29996 12164 30008
rect 12216 30036 12222 30048
rect 16114 30036 16120 30048
rect 12216 30008 16120 30036
rect 12216 29996 12222 30008
rect 16114 29996 16120 30008
rect 16172 29996 16178 30048
rect 16298 29996 16304 30048
rect 16356 30036 16362 30048
rect 16356 30008 16401 30036
rect 16356 29996 16362 30008
rect 19150 29996 19156 30048
rect 19208 30036 19214 30048
rect 20441 30039 20499 30045
rect 20441 30036 20453 30039
rect 19208 30008 20453 30036
rect 19208 29996 19214 30008
rect 20441 30005 20453 30008
rect 20487 30005 20499 30039
rect 20441 29999 20499 30005
rect 26878 29996 26884 30048
rect 26936 30036 26942 30048
rect 36280 30036 36308 30076
rect 37550 30064 37556 30076
rect 37608 30064 37614 30116
rect 26936 30008 36308 30036
rect 26936 29996 26942 30008
rect 36630 29996 36636 30048
rect 36688 30036 36694 30048
rect 36725 30039 36783 30045
rect 36725 30036 36737 30039
rect 36688 30008 36737 30036
rect 36688 29996 36694 30008
rect 36725 30005 36737 30008
rect 36771 30005 36783 30039
rect 36725 29999 36783 30005
rect 38105 30039 38163 30045
rect 38105 30005 38117 30039
rect 38151 30036 38163 30039
rect 38470 30036 38476 30048
rect 38151 30008 38476 30036
rect 38151 30005 38163 30008
rect 38105 29999 38163 30005
rect 38470 29996 38476 30008
rect 38528 29996 38534 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 11514 29832 11520 29844
rect 11475 29804 11520 29832
rect 11514 29792 11520 29804
rect 11572 29792 11578 29844
rect 14826 29832 14832 29844
rect 14787 29804 14832 29832
rect 14826 29792 14832 29804
rect 14884 29792 14890 29844
rect 19334 29832 19340 29844
rect 14936 29804 19340 29832
rect 2130 29724 2136 29776
rect 2188 29764 2194 29776
rect 9766 29764 9772 29776
rect 2188 29736 9772 29764
rect 2188 29724 2194 29736
rect 9766 29724 9772 29736
rect 9824 29724 9830 29776
rect 10873 29767 10931 29773
rect 10873 29733 10885 29767
rect 10919 29764 10931 29767
rect 14936 29764 14964 29804
rect 19334 29792 19340 29804
rect 19392 29792 19398 29844
rect 29178 29832 29184 29844
rect 19444 29804 29184 29832
rect 15378 29764 15384 29776
rect 10919 29736 14964 29764
rect 15028 29736 15384 29764
rect 10919 29733 10931 29736
rect 10873 29727 10931 29733
rect 9950 29656 9956 29708
rect 10008 29696 10014 29708
rect 11790 29696 11796 29708
rect 10008 29668 11796 29696
rect 10008 29656 10014 29668
rect 11790 29656 11796 29668
rect 11848 29656 11854 29708
rect 12250 29696 12256 29708
rect 12211 29668 12256 29696
rect 12250 29656 12256 29668
rect 12308 29656 12314 29708
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 1854 29628 1860 29640
rect 1627 29600 1860 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 1854 29588 1860 29600
rect 1912 29588 1918 29640
rect 10781 29631 10839 29637
rect 10781 29597 10793 29631
rect 10827 29628 10839 29631
rect 10870 29628 10876 29640
rect 10827 29600 10876 29628
rect 10827 29597 10839 29600
rect 10781 29591 10839 29597
rect 10870 29588 10876 29600
rect 10928 29588 10934 29640
rect 11422 29628 11428 29640
rect 11383 29600 11428 29628
rect 11422 29588 11428 29600
rect 11480 29588 11486 29640
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29628 14795 29631
rect 15028 29628 15056 29736
rect 15378 29724 15384 29736
rect 15436 29724 15442 29776
rect 16758 29724 16764 29776
rect 16816 29764 16822 29776
rect 19444 29764 19472 29804
rect 29178 29792 29184 29804
rect 29236 29792 29242 29844
rect 29840 29804 31064 29832
rect 16816 29736 19472 29764
rect 16816 29724 16822 29736
rect 26326 29724 26332 29776
rect 26384 29764 26390 29776
rect 29840 29764 29868 29804
rect 26384 29736 29868 29764
rect 31036 29764 31064 29804
rect 31202 29792 31208 29844
rect 31260 29832 31266 29844
rect 33965 29835 34023 29841
rect 33965 29832 33977 29835
rect 31260 29804 33977 29832
rect 31260 29792 31266 29804
rect 33965 29801 33977 29804
rect 34011 29801 34023 29835
rect 33965 29795 34023 29801
rect 31036 29736 32076 29764
rect 26384 29724 26390 29736
rect 15654 29656 15660 29708
rect 15712 29696 15718 29708
rect 16022 29696 16028 29708
rect 15712 29668 16028 29696
rect 15712 29656 15718 29668
rect 16022 29656 16028 29668
rect 16080 29656 16086 29708
rect 16114 29656 16120 29708
rect 16172 29696 16178 29708
rect 23014 29696 23020 29708
rect 16172 29668 23020 29696
rect 16172 29656 16178 29668
rect 23014 29656 23020 29668
rect 23072 29656 23078 29708
rect 26142 29656 26148 29708
rect 26200 29696 26206 29708
rect 29730 29696 29736 29708
rect 26200 29668 29736 29696
rect 26200 29656 26206 29668
rect 29730 29656 29736 29668
rect 29788 29656 29794 29708
rect 30466 29656 30472 29708
rect 30524 29696 30530 29708
rect 31757 29699 31815 29705
rect 31757 29696 31769 29699
rect 30524 29668 31769 29696
rect 30524 29656 30530 29668
rect 31757 29665 31769 29668
rect 31803 29665 31815 29699
rect 31757 29659 31815 29665
rect 14783 29600 15056 29628
rect 14783 29597 14795 29600
rect 14737 29591 14795 29597
rect 15102 29588 15108 29640
rect 15160 29628 15166 29640
rect 15381 29631 15439 29637
rect 15381 29628 15393 29631
rect 15160 29600 15393 29628
rect 15160 29588 15166 29600
rect 15381 29597 15393 29600
rect 15427 29597 15439 29631
rect 17402 29628 17408 29640
rect 17363 29600 17408 29628
rect 15381 29591 15439 29597
rect 17402 29588 17408 29600
rect 17460 29588 17466 29640
rect 20622 29628 20628 29640
rect 20583 29600 20628 29628
rect 20622 29588 20628 29600
rect 20680 29588 20686 29640
rect 27433 29631 27491 29637
rect 27433 29597 27445 29631
rect 27479 29628 27491 29631
rect 27614 29628 27620 29640
rect 27479 29600 27620 29628
rect 27479 29597 27491 29600
rect 27433 29591 27491 29597
rect 27614 29588 27620 29600
rect 27672 29588 27678 29640
rect 4065 29563 4123 29569
rect 4065 29529 4077 29563
rect 4111 29560 4123 29563
rect 7742 29560 7748 29572
rect 4111 29532 7748 29560
rect 4111 29529 4123 29532
rect 4065 29523 4123 29529
rect 7742 29520 7748 29532
rect 7800 29520 7806 29572
rect 9122 29520 9128 29572
rect 9180 29560 9186 29572
rect 12342 29560 12348 29572
rect 9180 29532 9996 29560
rect 12303 29532 12348 29560
rect 9180 29520 9186 29532
rect 1762 29492 1768 29504
rect 1723 29464 1768 29492
rect 1762 29452 1768 29464
rect 1820 29452 1826 29504
rect 4157 29495 4215 29501
rect 4157 29461 4169 29495
rect 4203 29492 4215 29495
rect 9858 29492 9864 29504
rect 4203 29464 9864 29492
rect 4203 29461 4215 29464
rect 4157 29455 4215 29461
rect 9858 29452 9864 29464
rect 9916 29452 9922 29504
rect 9968 29492 9996 29532
rect 12342 29520 12348 29532
rect 12400 29520 12406 29572
rect 13265 29563 13323 29569
rect 13265 29529 13277 29563
rect 13311 29560 13323 29563
rect 13446 29560 13452 29572
rect 13311 29532 13452 29560
rect 13311 29529 13323 29532
rect 13265 29523 13323 29529
rect 13446 29520 13452 29532
rect 13504 29520 13510 29572
rect 15654 29560 15660 29572
rect 13556 29532 15660 29560
rect 13556 29492 13584 29532
rect 15654 29520 15660 29532
rect 15712 29520 15718 29572
rect 15764 29532 16146 29560
rect 9968 29464 13584 29492
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 15764 29492 15792 29532
rect 16942 29520 16948 29572
rect 17000 29560 17006 29572
rect 20901 29563 20959 29569
rect 20901 29560 20913 29563
rect 17000 29532 20913 29560
rect 17000 29520 17006 29532
rect 20901 29529 20913 29532
rect 20947 29529 20959 29563
rect 20901 29523 20959 29529
rect 21174 29520 21180 29572
rect 21232 29560 21238 29572
rect 22649 29563 22707 29569
rect 21232 29532 21390 29560
rect 21232 29520 21238 29532
rect 22649 29529 22661 29563
rect 22695 29560 22707 29563
rect 23934 29560 23940 29572
rect 22695 29532 23940 29560
rect 22695 29529 22707 29532
rect 22649 29523 22707 29529
rect 23934 29520 23940 29532
rect 23992 29520 23998 29572
rect 25685 29563 25743 29569
rect 25685 29529 25697 29563
rect 25731 29560 25743 29563
rect 25731 29532 29224 29560
rect 25731 29529 25743 29532
rect 25685 29523 25743 29529
rect 13688 29464 15792 29492
rect 13688 29452 13694 29464
rect 16666 29452 16672 29504
rect 16724 29492 16730 29504
rect 26878 29492 26884 29504
rect 16724 29464 26884 29492
rect 16724 29452 16730 29464
rect 26878 29452 26884 29464
rect 26936 29452 26942 29504
rect 29196 29492 29224 29532
rect 29638 29520 29644 29572
rect 29696 29560 29702 29572
rect 30009 29563 30067 29569
rect 30009 29560 30021 29563
rect 29696 29532 30021 29560
rect 29696 29520 29702 29532
rect 30009 29529 30021 29532
rect 30055 29529 30067 29563
rect 31386 29560 31392 29572
rect 31234 29532 31392 29560
rect 30009 29523 30067 29529
rect 31386 29520 31392 29532
rect 31444 29520 31450 29572
rect 32048 29560 32076 29736
rect 32214 29696 32220 29708
rect 32175 29668 32220 29696
rect 32214 29656 32220 29668
rect 32272 29696 32278 29708
rect 34790 29696 34796 29708
rect 32272 29668 34796 29696
rect 32272 29656 32278 29668
rect 34790 29656 34796 29668
rect 34848 29696 34854 29708
rect 34885 29699 34943 29705
rect 34885 29696 34897 29699
rect 34848 29668 34897 29696
rect 34848 29656 34854 29668
rect 34885 29665 34897 29668
rect 34931 29665 34943 29699
rect 34885 29659 34943 29665
rect 32493 29563 32551 29569
rect 32493 29560 32505 29563
rect 32048 29532 32505 29560
rect 32493 29529 32505 29532
rect 32539 29529 32551 29563
rect 32493 29523 32551 29529
rect 32950 29520 32956 29572
rect 33008 29520 33014 29572
rect 35158 29560 35164 29572
rect 33796 29532 34100 29560
rect 35119 29532 35164 29560
rect 33796 29492 33824 29532
rect 29196 29464 33824 29492
rect 34072 29492 34100 29532
rect 35158 29520 35164 29532
rect 35216 29520 35222 29572
rect 36906 29560 36912 29572
rect 36386 29532 36492 29560
rect 36867 29532 36912 29560
rect 35434 29492 35440 29504
rect 34072 29464 35440 29492
rect 35434 29452 35440 29464
rect 35492 29452 35498 29504
rect 36464 29492 36492 29532
rect 36906 29520 36912 29532
rect 36964 29520 36970 29572
rect 38102 29560 38108 29572
rect 38063 29532 38108 29560
rect 38102 29520 38108 29532
rect 38160 29520 38166 29572
rect 36998 29492 37004 29504
rect 36464 29464 37004 29492
rect 36998 29452 37004 29464
rect 37056 29452 37062 29504
rect 38194 29492 38200 29504
rect 38155 29464 38200 29492
rect 38194 29452 38200 29464
rect 38252 29452 38258 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 4706 29288 4712 29300
rect 4667 29260 4712 29288
rect 4706 29248 4712 29260
rect 4764 29248 4770 29300
rect 11698 29288 11704 29300
rect 9784 29260 11704 29288
rect 8018 29180 8024 29232
rect 8076 29220 8082 29232
rect 9784 29229 9812 29260
rect 11698 29248 11704 29260
rect 11756 29248 11762 29300
rect 11793 29291 11851 29297
rect 11793 29257 11805 29291
rect 11839 29288 11851 29291
rect 12342 29288 12348 29300
rect 11839 29260 12348 29288
rect 11839 29257 11851 29260
rect 11793 29251 11851 29257
rect 12342 29248 12348 29260
rect 12400 29248 12406 29300
rect 16666 29288 16672 29300
rect 13004 29260 16672 29288
rect 9677 29223 9735 29229
rect 9677 29220 9689 29223
rect 8076 29192 9689 29220
rect 8076 29180 8082 29192
rect 9677 29189 9689 29192
rect 9723 29189 9735 29223
rect 9677 29183 9735 29189
rect 9769 29223 9827 29229
rect 9769 29189 9781 29223
rect 9815 29189 9827 29223
rect 9769 29183 9827 29189
rect 9858 29180 9864 29232
rect 9916 29220 9922 29232
rect 13004 29220 13032 29260
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 16850 29248 16856 29300
rect 16908 29288 16914 29300
rect 23106 29288 23112 29300
rect 16908 29260 23112 29288
rect 16908 29248 16914 29260
rect 13170 29220 13176 29232
rect 9916 29192 13032 29220
rect 13131 29192 13176 29220
rect 9916 29180 9922 29192
rect 13170 29180 13176 29192
rect 13228 29180 13234 29232
rect 14090 29220 14096 29232
rect 14051 29192 14096 29220
rect 14090 29180 14096 29192
rect 14148 29180 14154 29232
rect 16574 29180 16580 29232
rect 16632 29220 16638 29232
rect 20548 29229 20576 29260
rect 23106 29248 23112 29260
rect 23164 29248 23170 29300
rect 31294 29248 31300 29300
rect 31352 29288 31358 29300
rect 35158 29288 35164 29300
rect 31352 29260 35164 29288
rect 31352 29248 31358 29260
rect 35158 29248 35164 29260
rect 35216 29248 35222 29300
rect 20533 29223 20591 29229
rect 16632 29192 19090 29220
rect 16632 29180 16638 29192
rect 20533 29189 20545 29223
rect 20579 29189 20591 29223
rect 20533 29183 20591 29189
rect 28258 29180 28264 29232
rect 28316 29180 28322 29232
rect 34054 29180 34060 29232
rect 34112 29180 34118 29232
rect 4893 29155 4951 29161
rect 4893 29121 4905 29155
rect 4939 29152 4951 29155
rect 6822 29152 6828 29164
rect 4939 29124 6828 29152
rect 4939 29121 4951 29124
rect 4893 29115 4951 29121
rect 6822 29112 6828 29124
rect 6880 29112 6886 29164
rect 11054 29112 11060 29164
rect 11112 29152 11118 29164
rect 11701 29155 11759 29161
rect 11701 29152 11713 29155
rect 11112 29124 11713 29152
rect 11112 29112 11118 29124
rect 11701 29121 11713 29124
rect 11747 29152 11759 29155
rect 12250 29152 12256 29164
rect 11747 29124 12256 29152
rect 11747 29121 11759 29124
rect 11701 29115 11759 29121
rect 12250 29112 12256 29124
rect 12308 29112 12314 29164
rect 14553 29155 14611 29161
rect 14553 29121 14565 29155
rect 14599 29152 14611 29155
rect 14642 29152 14648 29164
rect 14599 29124 14648 29152
rect 14599 29121 14611 29124
rect 14553 29115 14611 29121
rect 14642 29112 14648 29124
rect 14700 29112 14706 29164
rect 16850 29152 16856 29164
rect 16811 29124 16856 29152
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 22002 29152 22008 29164
rect 21963 29124 22008 29152
rect 22002 29112 22008 29124
rect 22060 29112 22066 29164
rect 26142 29112 26148 29164
rect 26200 29152 26206 29164
rect 27249 29155 27307 29161
rect 27249 29152 27261 29155
rect 26200 29124 27261 29152
rect 26200 29112 26206 29124
rect 27249 29121 27261 29124
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 32214 29112 32220 29164
rect 32272 29152 32278 29164
rect 32769 29155 32827 29161
rect 32769 29152 32781 29155
rect 32272 29124 32781 29152
rect 32272 29112 32278 29124
rect 32769 29121 32781 29124
rect 32815 29121 32827 29155
rect 38286 29152 38292 29164
rect 38247 29124 38292 29152
rect 32769 29115 32827 29121
rect 38286 29112 38292 29124
rect 38344 29112 38350 29164
rect 1578 29084 1584 29096
rect 1539 29056 1584 29084
rect 1578 29044 1584 29056
rect 1636 29044 1642 29096
rect 1857 29087 1915 29093
rect 1857 29053 1869 29087
rect 1903 29084 1915 29087
rect 1946 29084 1952 29096
rect 1903 29056 1952 29084
rect 1903 29053 1915 29056
rect 1857 29047 1915 29053
rect 1946 29044 1952 29056
rect 2004 29044 2010 29096
rect 10689 29087 10747 29093
rect 10689 29053 10701 29087
rect 10735 29084 10747 29087
rect 10735 29056 12434 29084
rect 10735 29053 10747 29056
rect 10689 29047 10747 29053
rect 12406 29016 12434 29056
rect 12710 29044 12716 29096
rect 12768 29084 12774 29096
rect 13081 29087 13139 29093
rect 13081 29084 13093 29087
rect 12768 29056 13093 29084
rect 12768 29044 12774 29056
rect 13081 29053 13093 29056
rect 13127 29053 13139 29087
rect 13081 29047 13139 29053
rect 16390 29044 16396 29096
rect 16448 29084 16454 29096
rect 16942 29084 16948 29096
rect 16448 29056 16948 29084
rect 16448 29044 16454 29056
rect 16942 29044 16948 29056
rect 17000 29044 17006 29096
rect 17681 29087 17739 29093
rect 17681 29053 17693 29087
rect 17727 29084 17739 29087
rect 17770 29084 17776 29096
rect 17727 29056 17776 29084
rect 17727 29053 17739 29056
rect 17681 29047 17739 29053
rect 17770 29044 17776 29056
rect 17828 29044 17834 29096
rect 18138 29044 18144 29096
rect 18196 29084 18202 29096
rect 18325 29087 18383 29093
rect 18325 29084 18337 29087
rect 18196 29056 18337 29084
rect 18196 29044 18202 29056
rect 18325 29053 18337 29056
rect 18371 29053 18383 29087
rect 18325 29047 18383 29053
rect 18432 29056 19656 29084
rect 13446 29016 13452 29028
rect 12406 28988 13452 29016
rect 13446 28976 13452 28988
rect 13504 28976 13510 29028
rect 14642 29016 14648 29028
rect 14603 28988 14648 29016
rect 14642 28976 14648 28988
rect 14700 28976 14706 29028
rect 16114 28976 16120 29028
rect 16172 29016 16178 29028
rect 16172 28988 16620 29016
rect 16172 28976 16178 28988
rect 11422 28908 11428 28960
rect 11480 28948 11486 28960
rect 16482 28948 16488 28960
rect 11480 28920 16488 28948
rect 11480 28908 11486 28920
rect 16482 28908 16488 28920
rect 16540 28908 16546 28960
rect 16592 28948 16620 28988
rect 17494 28976 17500 29028
rect 17552 29016 17558 29028
rect 18432 29016 18460 29056
rect 17552 28988 18460 29016
rect 19628 29016 19656 29056
rect 20714 29044 20720 29096
rect 20772 29084 20778 29096
rect 21269 29087 21327 29093
rect 21269 29084 21281 29087
rect 20772 29056 21281 29084
rect 20772 29044 20778 29056
rect 21269 29053 21281 29056
rect 21315 29053 21327 29087
rect 21269 29047 21327 29053
rect 33134 29044 33140 29096
rect 33192 29084 33198 29096
rect 34517 29087 34575 29093
rect 34517 29084 34529 29087
rect 33192 29056 34529 29084
rect 33192 29044 33198 29056
rect 34517 29053 34529 29056
rect 34563 29053 34575 29087
rect 34517 29047 34575 29053
rect 36538 29044 36544 29096
rect 36596 29084 36602 29096
rect 39206 29084 39212 29096
rect 36596 29056 39212 29084
rect 36596 29044 36602 29056
rect 39206 29044 39212 29056
rect 39264 29044 39270 29096
rect 22097 29019 22155 29025
rect 22097 29016 22109 29019
rect 19628 28988 22109 29016
rect 17552 28976 17558 28988
rect 22097 28985 22109 28988
rect 22143 28985 22155 29019
rect 28994 29016 29000 29028
rect 28907 28988 29000 29016
rect 22097 28979 22155 28985
rect 28994 28976 29000 28988
rect 29052 29016 29058 29028
rect 29270 29016 29276 29028
rect 29052 28988 29276 29016
rect 29052 28976 29058 28988
rect 29270 28976 29276 28988
rect 29328 28976 29334 29028
rect 38102 29016 38108 29028
rect 38063 28988 38108 29016
rect 38102 28976 38108 28988
rect 38160 28976 38166 29028
rect 16758 28948 16764 28960
rect 16592 28920 16764 28948
rect 16758 28908 16764 28920
rect 16816 28908 16822 28960
rect 17954 28908 17960 28960
rect 18012 28948 18018 28960
rect 18582 28951 18640 28957
rect 18582 28948 18594 28951
rect 18012 28920 18594 28948
rect 18012 28908 18018 28920
rect 18582 28917 18594 28920
rect 18628 28948 18640 28951
rect 19150 28948 19156 28960
rect 18628 28920 19156 28948
rect 18628 28917 18640 28920
rect 18582 28911 18640 28917
rect 19150 28908 19156 28920
rect 19208 28908 19214 28960
rect 20070 28948 20076 28960
rect 20031 28920 20076 28948
rect 20070 28908 20076 28920
rect 20128 28908 20134 28960
rect 27338 28908 27344 28960
rect 27396 28948 27402 28960
rect 27506 28951 27564 28957
rect 27506 28948 27518 28951
rect 27396 28920 27518 28948
rect 27396 28908 27402 28920
rect 27506 28917 27518 28920
rect 27552 28917 27564 28951
rect 27506 28911 27564 28917
rect 33032 28951 33090 28957
rect 33032 28917 33044 28951
rect 33078 28948 33090 28951
rect 35434 28948 35440 28960
rect 33078 28920 35440 28948
rect 33078 28917 33090 28920
rect 33032 28911 33090 28917
rect 35434 28908 35440 28920
rect 35492 28908 35498 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 6822 28704 6828 28756
rect 6880 28744 6886 28756
rect 6917 28747 6975 28753
rect 6917 28744 6929 28747
rect 6880 28716 6929 28744
rect 6880 28704 6886 28716
rect 6917 28713 6929 28716
rect 6963 28713 6975 28747
rect 11238 28744 11244 28756
rect 11199 28716 11244 28744
rect 6917 28707 6975 28713
rect 11238 28704 11244 28716
rect 11296 28704 11302 28756
rect 32858 28744 32864 28756
rect 12406 28716 32864 28744
rect 8481 28679 8539 28685
rect 8481 28645 8493 28679
rect 8527 28676 8539 28679
rect 12406 28676 12434 28716
rect 32858 28704 32864 28716
rect 32916 28704 32922 28756
rect 8527 28648 12434 28676
rect 8527 28645 8539 28648
rect 8481 28639 8539 28645
rect 12526 28636 12532 28688
rect 12584 28676 12590 28688
rect 16114 28676 16120 28688
rect 12584 28648 16120 28676
rect 12584 28636 12590 28648
rect 16114 28636 16120 28648
rect 16172 28636 16178 28688
rect 7653 28611 7711 28617
rect 7653 28577 7665 28611
rect 7699 28608 7711 28611
rect 10045 28611 10103 28617
rect 10045 28608 10057 28611
rect 7699 28580 10057 28608
rect 7699 28577 7711 28580
rect 7653 28571 7711 28577
rect 10045 28577 10057 28580
rect 10091 28577 10103 28611
rect 10045 28571 10103 28577
rect 11882 28568 11888 28620
rect 11940 28608 11946 28620
rect 12069 28611 12127 28617
rect 12069 28608 12081 28611
rect 11940 28580 12081 28608
rect 11940 28568 11946 28580
rect 12069 28577 12081 28580
rect 12115 28577 12127 28611
rect 12069 28571 12127 28577
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 12492 28580 12537 28608
rect 12492 28568 12498 28580
rect 15102 28568 15108 28620
rect 15160 28608 15166 28620
rect 16209 28611 16267 28617
rect 16209 28608 16221 28611
rect 15160 28580 16221 28608
rect 15160 28568 15166 28580
rect 16209 28577 16221 28580
rect 16255 28608 16267 28611
rect 17770 28608 17776 28620
rect 16255 28580 17776 28608
rect 16255 28577 16267 28580
rect 16209 28571 16267 28577
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 20714 28608 20720 28620
rect 20364 28580 20720 28608
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28540 4583 28543
rect 4614 28540 4620 28552
rect 4571 28512 4620 28540
rect 4571 28509 4583 28512
rect 4525 28503 4583 28509
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 5169 28543 5227 28549
rect 5169 28509 5181 28543
rect 5215 28509 5227 28543
rect 5169 28503 5227 28509
rect 6825 28543 6883 28549
rect 6825 28509 6837 28543
rect 6871 28540 6883 28543
rect 7190 28540 7196 28552
rect 6871 28512 7196 28540
rect 6871 28509 6883 28512
rect 6825 28503 6883 28509
rect 5184 28472 5212 28503
rect 7190 28500 7196 28512
rect 7248 28500 7254 28552
rect 7558 28540 7564 28552
rect 7519 28512 7564 28540
rect 7558 28500 7564 28512
rect 7616 28500 7622 28552
rect 11149 28543 11207 28549
rect 11149 28509 11161 28543
rect 11195 28540 11207 28543
rect 11790 28540 11796 28552
rect 11195 28512 11796 28540
rect 11195 28509 11207 28512
rect 11149 28503 11207 28509
rect 11790 28500 11796 28512
rect 11848 28500 11854 28552
rect 13538 28540 13544 28552
rect 13499 28512 13544 28540
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 18138 28500 18144 28552
rect 18196 28540 18202 28552
rect 20364 28549 20392 28580
rect 20714 28568 20720 28580
rect 20772 28568 20778 28620
rect 32214 28568 32220 28620
rect 32272 28608 32278 28620
rect 32493 28611 32551 28617
rect 32493 28608 32505 28611
rect 32272 28580 32505 28608
rect 32272 28568 32278 28580
rect 32493 28577 32505 28580
rect 32539 28577 32551 28611
rect 32493 28571 32551 28577
rect 20349 28543 20407 28549
rect 20349 28540 20361 28543
rect 18196 28512 20361 28540
rect 18196 28500 18202 28512
rect 20349 28509 20361 28512
rect 20395 28509 20407 28543
rect 20349 28503 20407 28509
rect 4356 28444 5212 28472
rect 8297 28475 8355 28481
rect 4356 28413 4384 28444
rect 8297 28441 8309 28475
rect 8343 28472 8355 28475
rect 8386 28472 8392 28484
rect 8343 28444 8392 28472
rect 8343 28441 8355 28444
rect 8297 28435 8355 28441
rect 8386 28432 8392 28444
rect 8444 28432 8450 28484
rect 10042 28432 10048 28484
rect 10100 28472 10106 28484
rect 10137 28475 10195 28481
rect 10137 28472 10149 28475
rect 10100 28444 10149 28472
rect 10100 28432 10106 28444
rect 10137 28441 10149 28444
rect 10183 28441 10195 28475
rect 10137 28435 10195 28441
rect 10689 28475 10747 28481
rect 10689 28441 10701 28475
rect 10735 28472 10747 28475
rect 10778 28472 10784 28484
rect 10735 28444 10784 28472
rect 10735 28441 10747 28444
rect 10689 28435 10747 28441
rect 10778 28432 10784 28444
rect 10836 28432 10842 28484
rect 12161 28475 12219 28481
rect 12161 28441 12173 28475
rect 12207 28441 12219 28475
rect 12161 28435 12219 28441
rect 4341 28407 4399 28413
rect 4341 28373 4353 28407
rect 4387 28373 4399 28407
rect 4982 28404 4988 28416
rect 4943 28376 4988 28404
rect 4341 28367 4399 28373
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 12176 28404 12204 28435
rect 12250 28432 12256 28484
rect 12308 28472 12314 28484
rect 16482 28472 16488 28484
rect 12308 28444 16344 28472
rect 16443 28444 16488 28472
rect 12308 28432 12314 28444
rect 13633 28407 13691 28413
rect 13633 28404 13645 28407
rect 12176 28376 13645 28404
rect 13633 28373 13645 28376
rect 13679 28373 13691 28407
rect 16316 28404 16344 28444
rect 16482 28432 16488 28444
rect 16540 28432 16546 28484
rect 18506 28472 18512 28484
rect 17710 28444 18512 28472
rect 18506 28432 18512 28444
rect 18564 28432 18570 28484
rect 19426 28472 19432 28484
rect 19260 28444 19432 28472
rect 17957 28407 18015 28413
rect 17957 28404 17969 28407
rect 16316 28376 17969 28404
rect 13633 28367 13691 28373
rect 17957 28373 17969 28376
rect 18003 28404 18015 28407
rect 19260 28404 19288 28444
rect 19426 28432 19432 28444
rect 19484 28432 19490 28484
rect 20070 28432 20076 28484
rect 20128 28472 20134 28484
rect 20625 28475 20683 28481
rect 20625 28472 20637 28475
rect 20128 28444 20637 28472
rect 20128 28432 20134 28444
rect 20625 28441 20637 28444
rect 20671 28441 20683 28475
rect 32766 28472 32772 28484
rect 20625 28435 20683 28441
rect 20732 28444 21114 28472
rect 32727 28444 32772 28472
rect 18003 28376 19288 28404
rect 18003 28373 18015 28376
rect 17957 28367 18015 28373
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 20732 28404 20760 28444
rect 32766 28432 32772 28444
rect 32824 28472 32830 28484
rect 33042 28472 33048 28484
rect 32824 28444 33048 28472
rect 32824 28432 32830 28444
rect 33042 28432 33048 28444
rect 33100 28432 33106 28484
rect 33778 28432 33784 28484
rect 33836 28432 33842 28484
rect 19392 28376 20760 28404
rect 19392 28364 19398 28376
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 22097 28407 22155 28413
rect 22097 28404 22109 28407
rect 20864 28376 22109 28404
rect 20864 28364 20870 28376
rect 22097 28373 22109 28376
rect 22143 28373 22155 28407
rect 34238 28404 34244 28416
rect 34199 28376 34244 28404
rect 22097 28367 22155 28373
rect 34238 28364 34244 28376
rect 34296 28364 34302 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 11882 28200 11888 28212
rect 7760 28172 11888 28200
rect 7466 28024 7472 28076
rect 7524 28064 7530 28076
rect 7760 28073 7788 28172
rect 11882 28160 11888 28172
rect 11940 28160 11946 28212
rect 12526 28200 12532 28212
rect 12406 28172 12532 28200
rect 9306 28092 9312 28144
rect 9364 28092 9370 28144
rect 7745 28067 7803 28073
rect 7745 28064 7757 28067
rect 7524 28036 7757 28064
rect 7524 28024 7530 28036
rect 7745 28033 7757 28036
rect 7791 28033 7803 28067
rect 7745 28027 7803 28033
rect 9125 28067 9183 28073
rect 9125 28033 9137 28067
rect 9171 28064 9183 28067
rect 9324 28064 9352 28092
rect 9171 28036 9352 28064
rect 10229 28067 10287 28073
rect 9171 28033 9183 28036
rect 9125 28027 9183 28033
rect 10229 28033 10241 28067
rect 10275 28033 10287 28067
rect 10229 28027 10287 28033
rect 11701 28067 11759 28073
rect 11701 28033 11713 28067
rect 11747 28064 11759 28067
rect 12406 28064 12434 28172
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 16298 28200 16304 28212
rect 12636 28172 16304 28200
rect 11747 28036 12434 28064
rect 11747 28033 11759 28036
rect 11701 28027 11759 28033
rect 4982 27956 4988 28008
rect 5040 27996 5046 28008
rect 9309 27999 9367 28005
rect 9309 27996 9321 27999
rect 5040 27968 9321 27996
rect 5040 27956 5046 27968
rect 9309 27965 9321 27968
rect 9355 27965 9367 27999
rect 9309 27959 9367 27965
rect 10244 27928 10272 28027
rect 12636 27928 12664 28172
rect 16298 28160 16304 28172
rect 16356 28160 16362 28212
rect 16482 28160 16488 28212
rect 16540 28200 16546 28212
rect 23290 28200 23296 28212
rect 16540 28172 23296 28200
rect 16540 28160 16546 28172
rect 23290 28160 23296 28172
rect 23348 28160 23354 28212
rect 12989 28135 13047 28141
rect 12989 28101 13001 28135
rect 13035 28132 13047 28135
rect 14366 28132 14372 28144
rect 13035 28104 14372 28132
rect 13035 28101 13047 28104
rect 12989 28095 13047 28101
rect 14366 28092 14372 28104
rect 14424 28092 14430 28144
rect 15102 28132 15108 28144
rect 14568 28104 15108 28132
rect 14568 28076 14596 28104
rect 15102 28092 15108 28104
rect 15160 28092 15166 28144
rect 17494 28132 17500 28144
rect 16054 28104 17500 28132
rect 17494 28092 17500 28104
rect 17552 28092 17558 28144
rect 20530 28132 20536 28144
rect 19274 28104 20536 28132
rect 20530 28092 20536 28104
rect 20588 28092 20594 28144
rect 21358 28092 21364 28144
rect 21416 28132 21422 28144
rect 21416 28104 22770 28132
rect 21416 28092 21422 28104
rect 26878 28092 26884 28144
rect 26936 28132 26942 28144
rect 27430 28132 27436 28144
rect 26936 28104 27436 28132
rect 26936 28092 26942 28104
rect 27430 28092 27436 28104
rect 27488 28092 27494 28144
rect 28718 28132 28724 28144
rect 28658 28104 28724 28132
rect 28718 28092 28724 28104
rect 28776 28092 28782 28144
rect 29178 28132 29184 28144
rect 29091 28104 29184 28132
rect 29178 28092 29184 28104
rect 29236 28132 29242 28144
rect 29638 28132 29644 28144
rect 29236 28104 29644 28132
rect 29236 28092 29242 28104
rect 29638 28092 29644 28104
rect 29696 28092 29702 28144
rect 32490 28092 32496 28144
rect 32548 28132 32554 28144
rect 33413 28135 33471 28141
rect 33413 28132 33425 28135
rect 32548 28104 33425 28132
rect 32548 28092 32554 28104
rect 33413 28101 33425 28104
rect 33459 28101 33471 28135
rect 34790 28132 34796 28144
rect 34638 28104 34796 28132
rect 33413 28095 33471 28101
rect 34790 28092 34796 28104
rect 34848 28092 34854 28144
rect 14550 28064 14556 28076
rect 14463 28036 14556 28064
rect 14550 28024 14556 28036
rect 14608 28024 14614 28076
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 22005 28067 22063 28073
rect 22005 28064 22017 28067
rect 20772 28036 22017 28064
rect 20772 28024 20778 28036
rect 22005 28033 22017 28036
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 12897 27999 12955 28005
rect 12897 27965 12909 27999
rect 12943 27996 12955 27999
rect 13078 27996 13084 28008
rect 12943 27968 13084 27996
rect 12943 27965 12955 27968
rect 12897 27959 12955 27965
rect 13078 27956 13084 27968
rect 13136 27956 13142 28008
rect 13354 27996 13360 28008
rect 13315 27968 13360 27996
rect 13354 27956 13360 27968
rect 13412 27956 13418 28008
rect 14826 27956 14832 28008
rect 14884 27996 14890 28008
rect 14884 27968 14929 27996
rect 14884 27956 14890 27968
rect 15562 27956 15568 28008
rect 15620 27996 15626 28008
rect 17218 27996 17224 28008
rect 15620 27968 17224 27996
rect 15620 27956 15626 27968
rect 17218 27956 17224 27968
rect 17276 27956 17282 28008
rect 17770 27996 17776 28008
rect 17731 27968 17776 27996
rect 17770 27956 17776 27968
rect 17828 27956 17834 28008
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 17880 27968 18061 27996
rect 10244 27900 12664 27928
rect 7834 27860 7840 27872
rect 7795 27832 7840 27860
rect 7834 27820 7840 27832
rect 7892 27820 7898 27872
rect 7926 27820 7932 27872
rect 7984 27860 7990 27872
rect 9493 27863 9551 27869
rect 9493 27860 9505 27863
rect 7984 27832 9505 27860
rect 7984 27820 7990 27832
rect 9493 27829 9505 27832
rect 9539 27829 9551 27863
rect 10318 27860 10324 27872
rect 10279 27832 10324 27860
rect 9493 27823 9551 27829
rect 10318 27820 10324 27832
rect 10376 27820 10382 27872
rect 11514 27820 11520 27872
rect 11572 27860 11578 27872
rect 11793 27863 11851 27869
rect 11793 27860 11805 27863
rect 11572 27832 11805 27860
rect 11572 27820 11578 27832
rect 11793 27829 11805 27832
rect 11839 27829 11851 27863
rect 11793 27823 11851 27829
rect 11882 27820 11888 27872
rect 11940 27860 11946 27872
rect 16301 27863 16359 27869
rect 16301 27860 16313 27863
rect 11940 27832 16313 27860
rect 11940 27820 11946 27832
rect 16301 27829 16313 27832
rect 16347 27860 16359 27863
rect 17880 27860 17908 27968
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 18414 27956 18420 28008
rect 18472 27996 18478 28008
rect 19797 27999 19855 28005
rect 19797 27996 19809 27999
rect 18472 27968 19809 27996
rect 18472 27956 18478 27968
rect 19797 27965 19809 27968
rect 19843 27965 19855 27999
rect 19797 27959 19855 27965
rect 20162 27956 20168 28008
rect 20220 27996 20226 28008
rect 24029 27999 24087 28005
rect 24029 27996 24041 27999
rect 20220 27968 24041 27996
rect 20220 27956 20226 27968
rect 24029 27965 24041 27968
rect 24075 27996 24087 27999
rect 26326 27996 26332 28008
rect 24075 27968 26332 27996
rect 24075 27965 24087 27968
rect 24029 27959 24087 27965
rect 26326 27956 26332 27968
rect 26384 27956 26390 28008
rect 26418 27956 26424 28008
rect 26476 27996 26482 28008
rect 27157 27999 27215 28005
rect 27157 27996 27169 27999
rect 26476 27968 27169 27996
rect 26476 27956 26482 27968
rect 27157 27965 27169 27968
rect 27203 27965 27215 27999
rect 33134 27996 33140 28008
rect 33095 27968 33140 27996
rect 27157 27959 27215 27965
rect 33134 27956 33140 27968
rect 33192 27956 33198 28008
rect 19242 27888 19248 27940
rect 19300 27928 19306 27940
rect 20806 27928 20812 27940
rect 19300 27900 20812 27928
rect 19300 27888 19306 27900
rect 20806 27888 20812 27900
rect 20864 27888 20870 27940
rect 16347 27832 17908 27860
rect 22268 27863 22326 27869
rect 16347 27829 16359 27832
rect 16301 27823 16359 27829
rect 22268 27829 22280 27863
rect 22314 27860 22326 27863
rect 30466 27860 30472 27872
rect 22314 27832 30472 27860
rect 22314 27829 22326 27832
rect 22268 27823 22326 27829
rect 30466 27820 30472 27832
rect 30524 27860 30530 27872
rect 30926 27860 30932 27872
rect 30524 27832 30932 27860
rect 30524 27820 30530 27832
rect 30926 27820 30932 27832
rect 30984 27820 30990 27872
rect 33870 27820 33876 27872
rect 33928 27860 33934 27872
rect 34885 27863 34943 27869
rect 34885 27860 34897 27863
rect 33928 27832 34897 27860
rect 33928 27820 33934 27832
rect 34885 27829 34897 27832
rect 34931 27829 34943 27863
rect 34885 27823 34943 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 4614 27616 4620 27668
rect 4672 27656 4678 27668
rect 7098 27656 7104 27668
rect 4672 27628 7104 27656
rect 4672 27616 4678 27628
rect 7098 27616 7104 27628
rect 7156 27616 7162 27668
rect 7190 27616 7196 27668
rect 7248 27656 7254 27668
rect 7248 27628 7696 27656
rect 7248 27616 7254 27628
rect 7285 27591 7343 27597
rect 7285 27557 7297 27591
rect 7331 27557 7343 27591
rect 7668 27588 7696 27628
rect 13538 27616 13544 27668
rect 13596 27656 13602 27668
rect 15920 27659 15978 27665
rect 15920 27656 15932 27659
rect 13596 27628 15932 27656
rect 13596 27616 13602 27628
rect 15920 27625 15932 27628
rect 15966 27656 15978 27659
rect 25958 27656 25964 27668
rect 15966 27628 25964 27656
rect 15966 27625 15978 27628
rect 15920 27619 15978 27625
rect 25958 27616 25964 27628
rect 26016 27616 26022 27668
rect 27154 27616 27160 27668
rect 27212 27656 27218 27668
rect 32842 27659 32900 27665
rect 32842 27656 32854 27659
rect 27212 27628 32854 27656
rect 27212 27616 27218 27628
rect 32842 27625 32854 27628
rect 32888 27625 32900 27659
rect 32842 27619 32900 27625
rect 34606 27616 34612 27668
rect 34664 27656 34670 27668
rect 35148 27659 35206 27665
rect 35148 27656 35160 27659
rect 34664 27628 35160 27656
rect 34664 27616 34670 27628
rect 35148 27625 35160 27628
rect 35194 27656 35206 27659
rect 36906 27656 36912 27668
rect 35194 27628 36912 27656
rect 35194 27625 35206 27628
rect 35148 27619 35206 27625
rect 36906 27616 36912 27628
rect 36964 27616 36970 27668
rect 8297 27591 8355 27597
rect 8297 27588 8309 27591
rect 7668 27560 8309 27588
rect 7285 27551 7343 27557
rect 8297 27557 8309 27560
rect 8343 27557 8355 27591
rect 8297 27551 8355 27557
rect 6825 27455 6883 27461
rect 6825 27421 6837 27455
rect 6871 27452 6883 27455
rect 7300 27452 7328 27551
rect 12894 27548 12900 27600
rect 12952 27548 12958 27600
rect 14366 27588 14372 27600
rect 14327 27560 14372 27588
rect 14366 27548 14372 27560
rect 14424 27548 14430 27600
rect 14826 27548 14832 27600
rect 14884 27588 14890 27600
rect 15378 27588 15384 27600
rect 14884 27560 15384 27588
rect 14884 27548 14890 27560
rect 15378 27548 15384 27560
rect 15436 27548 15442 27600
rect 7834 27480 7840 27532
rect 7892 27520 7898 27532
rect 8113 27523 8171 27529
rect 8113 27520 8125 27523
rect 7892 27492 8125 27520
rect 7892 27480 7898 27492
rect 8113 27489 8125 27492
rect 8159 27489 8171 27523
rect 12912 27520 12940 27548
rect 12989 27523 13047 27529
rect 12989 27520 13001 27523
rect 12912 27492 13001 27520
rect 8113 27483 8171 27489
rect 12989 27489 13001 27492
rect 13035 27489 13047 27523
rect 12989 27483 13047 27489
rect 13170 27480 13176 27532
rect 13228 27520 13234 27532
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 13228 27492 13277 27520
rect 13228 27480 13234 27492
rect 13265 27489 13277 27492
rect 13311 27489 13323 27523
rect 13265 27483 13323 27489
rect 14090 27480 14096 27532
rect 14148 27520 14154 27532
rect 14844 27520 14872 27548
rect 14148 27492 14872 27520
rect 15657 27523 15715 27529
rect 14148 27480 14154 27492
rect 15657 27489 15669 27523
rect 15703 27520 15715 27523
rect 17770 27520 17776 27532
rect 15703 27492 17776 27520
rect 15703 27489 15715 27492
rect 15657 27483 15715 27489
rect 17770 27480 17776 27492
rect 17828 27520 17834 27532
rect 19429 27523 19487 27529
rect 19429 27520 19441 27523
rect 17828 27492 19441 27520
rect 17828 27480 17834 27492
rect 19429 27489 19441 27492
rect 19475 27489 19487 27523
rect 19429 27483 19487 27489
rect 21177 27523 21235 27529
rect 21177 27489 21189 27523
rect 21223 27520 21235 27523
rect 23198 27520 23204 27532
rect 21223 27492 23204 27520
rect 21223 27489 21235 27492
rect 21177 27483 21235 27489
rect 23198 27480 23204 27492
rect 23256 27480 23262 27532
rect 23290 27480 23296 27532
rect 23348 27520 23354 27532
rect 28445 27523 28503 27529
rect 28445 27520 28457 27523
rect 23348 27492 28457 27520
rect 23348 27480 23354 27492
rect 28445 27489 28457 27492
rect 28491 27489 28503 27523
rect 28445 27483 28503 27489
rect 30101 27523 30159 27529
rect 30101 27489 30113 27523
rect 30147 27520 30159 27523
rect 31110 27520 31116 27532
rect 30147 27492 31116 27520
rect 30147 27489 30159 27492
rect 30101 27483 30159 27489
rect 31110 27480 31116 27492
rect 31168 27480 31174 27532
rect 32585 27523 32643 27529
rect 32585 27489 32597 27523
rect 32631 27520 32643 27523
rect 33226 27520 33232 27532
rect 32631 27492 33232 27520
rect 32631 27489 32643 27492
rect 32585 27483 32643 27489
rect 33226 27480 33232 27492
rect 33284 27480 33290 27532
rect 37274 27520 37280 27532
rect 33980 27492 37280 27520
rect 7466 27452 7472 27464
rect 6871 27424 7328 27452
rect 7427 27424 7472 27452
rect 6871 27421 6883 27424
rect 6825 27415 6883 27421
rect 7466 27412 7472 27424
rect 7524 27412 7530 27464
rect 7926 27452 7932 27464
rect 7887 27424 7932 27452
rect 7926 27412 7932 27424
rect 7984 27412 7990 27464
rect 12069 27455 12127 27461
rect 12069 27421 12081 27455
rect 12115 27452 12127 27455
rect 12342 27452 12348 27464
rect 12115 27424 12348 27452
rect 12115 27421 12127 27424
rect 12069 27415 12127 27421
rect 12342 27412 12348 27424
rect 12400 27452 12406 27464
rect 12802 27452 12808 27464
rect 12400 27424 12808 27452
rect 12400 27412 12406 27424
rect 12802 27412 12808 27424
rect 12860 27412 12866 27464
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27452 14335 27455
rect 15562 27452 15568 27464
rect 14323 27424 15568 27452
rect 14323 27421 14335 27424
rect 14277 27415 14335 27421
rect 15562 27412 15568 27424
rect 15620 27412 15626 27464
rect 26418 27412 26424 27464
rect 26476 27452 26482 27464
rect 26697 27455 26755 27461
rect 26697 27452 26709 27455
rect 26476 27424 26709 27452
rect 26476 27412 26482 27424
rect 26697 27421 26709 27424
rect 26743 27421 26755 27455
rect 32398 27452 32404 27464
rect 31510 27424 32404 27452
rect 26697 27415 26755 27421
rect 32398 27412 32404 27424
rect 32456 27412 32462 27464
rect 33980 27438 34008 27492
rect 37274 27480 37280 27492
rect 37332 27480 37338 27532
rect 34422 27412 34428 27464
rect 34480 27452 34486 27464
rect 34885 27455 34943 27461
rect 34885 27452 34897 27455
rect 34480 27424 34897 27452
rect 34480 27412 34486 27424
rect 34885 27421 34897 27424
rect 34931 27421 34943 27455
rect 38286 27452 38292 27464
rect 38247 27424 38292 27452
rect 34885 27415 34943 27421
rect 38286 27412 38292 27424
rect 38344 27412 38350 27464
rect 1670 27384 1676 27396
rect 1631 27356 1676 27384
rect 1670 27344 1676 27356
rect 1728 27344 1734 27396
rect 1857 27387 1915 27393
rect 1857 27353 1869 27387
rect 1903 27384 1915 27387
rect 5442 27384 5448 27396
rect 1903 27356 5448 27384
rect 1903 27353 1915 27356
rect 1857 27347 1915 27353
rect 5442 27344 5448 27356
rect 5500 27344 5506 27396
rect 10226 27344 10232 27396
rect 10284 27384 10290 27396
rect 11425 27387 11483 27393
rect 11425 27384 11437 27387
rect 10284 27356 11437 27384
rect 10284 27344 10290 27356
rect 11425 27353 11437 27356
rect 11471 27353 11483 27387
rect 11425 27347 11483 27353
rect 11514 27344 11520 27396
rect 11572 27384 11578 27396
rect 13078 27384 13084 27396
rect 11572 27356 11617 27384
rect 13039 27356 13084 27384
rect 11572 27344 11578 27356
rect 13078 27344 13084 27356
rect 13136 27344 13142 27396
rect 19705 27387 19763 27393
rect 15856 27356 16422 27384
rect 6641 27319 6699 27325
rect 6641 27285 6653 27319
rect 6687 27316 6699 27319
rect 7006 27316 7012 27328
rect 6687 27288 7012 27316
rect 6687 27285 6699 27288
rect 6641 27279 6699 27285
rect 7006 27276 7012 27288
rect 7064 27276 7070 27328
rect 12066 27276 12072 27328
rect 12124 27316 12130 27328
rect 15856 27316 15884 27356
rect 19705 27353 19717 27387
rect 19751 27353 19763 27387
rect 22462 27384 22468 27396
rect 20930 27356 22468 27384
rect 19705 27347 19763 27353
rect 17402 27316 17408 27328
rect 12124 27288 15884 27316
rect 17363 27288 17408 27316
rect 12124 27276 12130 27288
rect 17402 27276 17408 27288
rect 17460 27276 17466 27328
rect 19720 27316 19748 27347
rect 22462 27344 22468 27356
rect 22520 27344 22526 27396
rect 26970 27384 26976 27396
rect 26931 27356 26976 27384
rect 26970 27344 26976 27356
rect 27028 27344 27034 27396
rect 29086 27384 29092 27396
rect 28198 27356 29092 27384
rect 29086 27344 29092 27356
rect 29144 27344 29150 27396
rect 30377 27387 30435 27393
rect 30377 27353 30389 27387
rect 30423 27384 30435 27387
rect 30466 27384 30472 27396
rect 30423 27356 30472 27384
rect 30423 27353 30435 27356
rect 30377 27347 30435 27353
rect 30466 27344 30472 27356
rect 30524 27344 30530 27396
rect 31662 27344 31668 27396
rect 31720 27384 31726 27396
rect 32125 27387 32183 27393
rect 32125 27384 32137 27387
rect 31720 27356 32137 27384
rect 31720 27344 31726 27356
rect 32125 27353 32137 27356
rect 32171 27353 32183 27387
rect 39574 27384 39580 27396
rect 36386 27356 39580 27384
rect 32125 27347 32183 27353
rect 39574 27344 39580 27356
rect 39632 27344 39638 27396
rect 21542 27316 21548 27328
rect 19720 27288 21548 27316
rect 21542 27276 21548 27288
rect 21600 27276 21606 27328
rect 31754 27276 31760 27328
rect 31812 27316 31818 27328
rect 32306 27316 32312 27328
rect 31812 27288 32312 27316
rect 31812 27276 31818 27288
rect 32306 27276 32312 27288
rect 32364 27316 32370 27328
rect 34333 27319 34391 27325
rect 34333 27316 34345 27319
rect 32364 27288 34345 27316
rect 32364 27276 32370 27288
rect 34333 27285 34345 27288
rect 34379 27285 34391 27319
rect 34333 27279 34391 27285
rect 35526 27276 35532 27328
rect 35584 27316 35590 27328
rect 36633 27319 36691 27325
rect 36633 27316 36645 27319
rect 35584 27288 36645 27316
rect 35584 27276 35590 27288
rect 36633 27285 36645 27288
rect 36679 27285 36691 27319
rect 36633 27279 36691 27285
rect 38105 27319 38163 27325
rect 38105 27285 38117 27319
rect 38151 27316 38163 27319
rect 39298 27316 39304 27328
rect 38151 27288 39304 27316
rect 38151 27285 38163 27288
rect 38105 27279 38163 27285
rect 39298 27276 39304 27288
rect 39356 27276 39362 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 12066 27112 12072 27124
rect 12027 27084 12072 27112
rect 12066 27072 12072 27084
rect 12124 27072 12130 27124
rect 13078 27072 13084 27124
rect 13136 27112 13142 27124
rect 16945 27115 17003 27121
rect 16945 27112 16957 27115
rect 13136 27084 16957 27112
rect 13136 27072 13142 27084
rect 16945 27081 16957 27084
rect 16991 27081 17003 27115
rect 16945 27075 17003 27081
rect 20530 27072 20536 27124
rect 20588 27112 20594 27124
rect 21361 27115 21419 27121
rect 21361 27112 21373 27115
rect 20588 27084 21373 27112
rect 20588 27072 20594 27084
rect 21361 27081 21373 27084
rect 21407 27081 21419 27115
rect 21361 27075 21419 27081
rect 21542 27072 21548 27124
rect 21600 27112 21606 27124
rect 31662 27112 31668 27124
rect 21600 27084 31668 27112
rect 21600 27072 21606 27084
rect 31662 27072 31668 27084
rect 31720 27072 31726 27124
rect 34606 27112 34612 27124
rect 32968 27084 34612 27112
rect 6822 27004 6828 27056
rect 6880 27044 6886 27056
rect 8481 27047 8539 27053
rect 8481 27044 8493 27047
rect 6880 27016 8493 27044
rect 6880 27004 6886 27016
rect 8481 27013 8493 27016
rect 8527 27013 8539 27047
rect 8481 27007 8539 27013
rect 8573 27047 8631 27053
rect 8573 27013 8585 27047
rect 8619 27044 8631 27047
rect 10318 27044 10324 27056
rect 8619 27016 10324 27044
rect 8619 27013 8631 27016
rect 8573 27007 8631 27013
rect 10318 27004 10324 27016
rect 10376 27004 10382 27056
rect 11514 27004 11520 27056
rect 11572 27044 11578 27056
rect 12710 27044 12716 27056
rect 11572 27016 12716 27044
rect 11572 27004 11578 27016
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 14182 27004 14188 27056
rect 14240 27044 14246 27056
rect 14240 27016 15318 27044
rect 14240 27004 14246 27016
rect 18874 27004 18880 27056
rect 18932 27004 18938 27056
rect 7006 26976 7012 26988
rect 6967 26948 7012 26976
rect 7006 26936 7012 26948
rect 7064 26936 7070 26988
rect 11977 26979 12035 26985
rect 11977 26945 11989 26979
rect 12023 26976 12035 26979
rect 12802 26976 12808 26988
rect 12023 26948 12808 26976
rect 12023 26945 12035 26948
rect 11977 26939 12035 26945
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 14550 26976 14556 26988
rect 14511 26948 14556 26976
rect 14550 26936 14556 26948
rect 14608 26936 14614 26988
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26976 16911 26979
rect 17954 26976 17960 26988
rect 16899 26948 17960 26976
rect 16899 26945 16911 26948
rect 16853 26939 16911 26945
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18138 26976 18144 26988
rect 18099 26948 18144 26976
rect 18138 26936 18144 26948
rect 18196 26936 18202 26988
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26976 21327 26979
rect 22002 26976 22008 26988
rect 21315 26948 22008 26976
rect 21315 26945 21327 26948
rect 21269 26939 21327 26945
rect 22002 26936 22008 26948
rect 22060 26936 22066 26988
rect 27614 26976 27620 26988
rect 27575 26948 27620 26976
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 5994 26868 6000 26920
rect 6052 26908 6058 26920
rect 6825 26911 6883 26917
rect 6825 26908 6837 26911
rect 6052 26880 6837 26908
rect 6052 26868 6058 26880
rect 6825 26877 6837 26880
rect 6871 26877 6883 26911
rect 6825 26871 6883 26877
rect 9493 26911 9551 26917
rect 9493 26877 9505 26911
rect 9539 26908 9551 26911
rect 10042 26908 10048 26920
rect 9539 26880 10048 26908
rect 9539 26877 9551 26880
rect 9493 26871 9551 26877
rect 10042 26868 10048 26880
rect 10100 26908 10106 26920
rect 10686 26908 10692 26920
rect 10100 26880 10692 26908
rect 10100 26868 10106 26880
rect 10686 26868 10692 26880
rect 10744 26868 10750 26920
rect 14090 26908 14096 26920
rect 10888 26880 14096 26908
rect 7190 26840 7196 26852
rect 7151 26812 7196 26840
rect 7190 26800 7196 26812
rect 7248 26800 7254 26852
rect 10888 26784 10916 26880
rect 14090 26868 14096 26880
rect 14148 26868 14154 26920
rect 14829 26911 14887 26917
rect 14829 26877 14841 26911
rect 14875 26908 14887 26911
rect 16298 26908 16304 26920
rect 14875 26880 16304 26908
rect 14875 26877 14887 26880
rect 14829 26871 14887 26877
rect 16298 26868 16304 26880
rect 16356 26868 16362 26920
rect 18046 26868 18052 26920
rect 18104 26908 18110 26920
rect 18414 26908 18420 26920
rect 18104 26880 18420 26908
rect 18104 26868 18110 26880
rect 18414 26868 18420 26880
rect 18472 26868 18478 26920
rect 26418 26868 26424 26920
rect 26476 26908 26482 26920
rect 28353 26911 28411 26917
rect 28353 26908 28365 26911
rect 26476 26880 28365 26908
rect 26476 26868 26482 26880
rect 28353 26877 28365 26880
rect 28399 26908 28411 26911
rect 29362 26908 29368 26920
rect 28399 26880 29368 26908
rect 28399 26877 28411 26880
rect 28353 26871 28411 26877
rect 29362 26868 29368 26880
rect 29420 26908 29426 26920
rect 29549 26911 29607 26917
rect 29549 26908 29561 26911
rect 29420 26880 29561 26908
rect 29420 26868 29426 26880
rect 29549 26877 29561 26880
rect 29595 26877 29607 26911
rect 29825 26911 29883 26917
rect 29825 26908 29837 26911
rect 29549 26871 29607 26877
rect 29656 26880 29837 26908
rect 15838 26800 15844 26852
rect 15896 26840 15902 26852
rect 17310 26840 17316 26852
rect 15896 26812 17316 26840
rect 15896 26800 15902 26812
rect 17310 26800 17316 26812
rect 17368 26800 17374 26852
rect 21450 26840 21456 26852
rect 19904 26812 21456 26840
rect 7098 26732 7104 26784
rect 7156 26772 7162 26784
rect 10870 26772 10876 26784
rect 7156 26744 10876 26772
rect 7156 26732 7162 26744
rect 10870 26732 10876 26744
rect 10928 26732 10934 26784
rect 11790 26732 11796 26784
rect 11848 26772 11854 26784
rect 15930 26772 15936 26784
rect 11848 26744 15936 26772
rect 11848 26732 11854 26744
rect 15930 26732 15936 26744
rect 15988 26732 15994 26784
rect 16301 26775 16359 26781
rect 16301 26741 16313 26775
rect 16347 26772 16359 26775
rect 16390 26772 16396 26784
rect 16347 26744 16396 26772
rect 16347 26741 16359 26744
rect 16301 26735 16359 26741
rect 16390 26732 16396 26744
rect 16448 26732 16454 26784
rect 18782 26732 18788 26784
rect 18840 26772 18846 26784
rect 19904 26781 19932 26812
rect 21450 26800 21456 26812
rect 21508 26800 21514 26852
rect 29656 26840 29684 26880
rect 29825 26877 29837 26880
rect 29871 26908 29883 26911
rect 30374 26908 30380 26920
rect 29871 26880 30380 26908
rect 29871 26877 29883 26880
rect 29825 26871 29883 26877
rect 30374 26868 30380 26880
rect 30432 26868 30438 26920
rect 30944 26908 30972 26962
rect 31018 26908 31024 26920
rect 30944 26880 31024 26908
rect 31018 26868 31024 26880
rect 31076 26868 31082 26920
rect 22066 26812 29684 26840
rect 19889 26775 19947 26781
rect 19889 26772 19901 26775
rect 18840 26744 19901 26772
rect 18840 26732 18846 26744
rect 19889 26741 19901 26744
rect 19935 26741 19947 26775
rect 19889 26735 19947 26741
rect 20530 26732 20536 26784
rect 20588 26772 20594 26784
rect 22066 26772 22094 26812
rect 30834 26800 30840 26852
rect 30892 26840 30898 26852
rect 32968 26840 32996 27084
rect 34606 27072 34612 27084
rect 34664 27072 34670 27124
rect 33042 27004 33048 27056
rect 33100 27044 33106 27056
rect 33781 27047 33839 27053
rect 33781 27044 33793 27047
rect 33100 27016 33793 27044
rect 33100 27004 33106 27016
rect 33781 27013 33793 27016
rect 33827 27013 33839 27047
rect 38562 27044 38568 27056
rect 35006 27016 38568 27044
rect 33781 27007 33839 27013
rect 38562 27004 38568 27016
rect 38620 27004 38626 27056
rect 33134 26868 33140 26920
rect 33192 26908 33198 26920
rect 33505 26911 33563 26917
rect 33505 26908 33517 26911
rect 33192 26880 33517 26908
rect 33192 26868 33198 26880
rect 33505 26877 33517 26880
rect 33551 26877 33563 26911
rect 33505 26871 33563 26877
rect 35529 26911 35587 26917
rect 35529 26877 35541 26911
rect 35575 26908 35587 26911
rect 35618 26908 35624 26920
rect 35575 26880 35624 26908
rect 35575 26877 35587 26880
rect 35529 26871 35587 26877
rect 30892 26812 32996 26840
rect 30892 26800 30898 26812
rect 20588 26744 22094 26772
rect 20588 26732 20594 26744
rect 30190 26732 30196 26784
rect 30248 26772 30254 26784
rect 31294 26772 31300 26784
rect 30248 26744 31300 26772
rect 30248 26732 30254 26744
rect 31294 26732 31300 26744
rect 31352 26732 31358 26784
rect 33520 26772 33548 26871
rect 35618 26868 35624 26880
rect 35676 26868 35682 26920
rect 33594 26772 33600 26784
rect 33507 26744 33600 26772
rect 33594 26732 33600 26744
rect 33652 26772 33658 26784
rect 34422 26772 34428 26784
rect 33652 26744 34428 26772
rect 33652 26732 33658 26744
rect 34422 26732 34428 26744
rect 34480 26732 34486 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1581 26571 1639 26577
rect 1581 26537 1593 26571
rect 1627 26568 1639 26571
rect 7558 26568 7564 26580
rect 1627 26540 7564 26568
rect 1627 26537 1639 26540
rect 1581 26531 1639 26537
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 22738 26568 22744 26580
rect 10336 26540 22744 26568
rect 7837 26503 7895 26509
rect 7837 26469 7849 26503
rect 7883 26500 7895 26503
rect 10226 26500 10232 26512
rect 7883 26472 10232 26500
rect 7883 26469 7895 26472
rect 7837 26463 7895 26469
rect 10226 26460 10232 26472
rect 10284 26460 10290 26512
rect 6822 26392 6828 26444
rect 6880 26432 6886 26444
rect 9217 26435 9275 26441
rect 9217 26432 9229 26435
rect 6880 26404 9229 26432
rect 6880 26392 6886 26404
rect 9217 26401 9229 26404
rect 9263 26401 9275 26435
rect 9217 26395 9275 26401
rect 1762 26364 1768 26376
rect 1723 26336 1768 26364
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 4706 26324 4712 26376
rect 4764 26364 4770 26376
rect 5442 26364 5448 26376
rect 4764 26336 5448 26364
rect 4764 26324 4770 26336
rect 5442 26324 5448 26336
rect 5500 26364 5506 26376
rect 7745 26367 7803 26373
rect 7745 26364 7757 26367
rect 5500 26336 7757 26364
rect 5500 26324 5506 26336
rect 7745 26333 7757 26336
rect 7791 26333 7803 26367
rect 7745 26327 7803 26333
rect 8846 26324 8852 26376
rect 8904 26364 8910 26376
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8904 26336 9137 26364
rect 8904 26324 8910 26336
rect 9125 26333 9137 26336
rect 9171 26364 9183 26367
rect 10336 26364 10364 26540
rect 22738 26528 22744 26540
rect 22796 26528 22802 26580
rect 27801 26571 27859 26577
rect 27801 26537 27813 26571
rect 27847 26568 27859 26571
rect 34698 26568 34704 26580
rect 27847 26540 34704 26568
rect 27847 26537 27859 26540
rect 27801 26531 27859 26537
rect 34698 26528 34704 26540
rect 34756 26528 34762 26580
rect 12710 26460 12716 26512
rect 12768 26500 12774 26512
rect 15562 26500 15568 26512
rect 12768 26472 15568 26500
rect 12768 26460 12774 26472
rect 15562 26460 15568 26472
rect 15620 26460 15626 26512
rect 27430 26460 27436 26512
rect 27488 26500 27494 26512
rect 30834 26500 30840 26512
rect 27488 26472 30840 26500
rect 27488 26460 27494 26472
rect 30834 26460 30840 26472
rect 30892 26460 30898 26512
rect 33042 26460 33048 26512
rect 33100 26500 33106 26512
rect 33229 26503 33287 26509
rect 33229 26500 33241 26503
rect 33100 26472 33241 26500
rect 33100 26460 33106 26472
rect 33229 26469 33241 26472
rect 33275 26469 33287 26503
rect 33229 26463 33287 26469
rect 38105 26503 38163 26509
rect 38105 26469 38117 26503
rect 38151 26500 38163 26503
rect 39390 26500 39396 26512
rect 38151 26472 39396 26500
rect 38151 26469 38163 26472
rect 38105 26463 38163 26469
rect 39390 26460 39396 26472
rect 39448 26460 39454 26512
rect 10686 26392 10692 26444
rect 10744 26432 10750 26444
rect 13354 26432 13360 26444
rect 10744 26404 13360 26432
rect 10744 26392 10750 26404
rect 13354 26392 13360 26404
rect 13412 26392 13418 26444
rect 14550 26392 14556 26444
rect 14608 26432 14614 26444
rect 15657 26435 15715 26441
rect 15657 26432 15669 26435
rect 14608 26404 15669 26432
rect 14608 26392 14614 26404
rect 15657 26401 15669 26404
rect 15703 26401 15715 26435
rect 15930 26432 15936 26444
rect 15843 26404 15936 26432
rect 15657 26395 15715 26401
rect 15930 26392 15936 26404
rect 15988 26432 15994 26444
rect 17402 26432 17408 26444
rect 15988 26404 17408 26432
rect 15988 26392 15994 26404
rect 17402 26392 17408 26404
rect 17460 26392 17466 26444
rect 20714 26432 20720 26444
rect 20675 26404 20720 26432
rect 20714 26392 20720 26404
rect 20772 26392 20778 26444
rect 22741 26435 22799 26441
rect 22741 26401 22753 26435
rect 22787 26432 22799 26435
rect 22830 26432 22836 26444
rect 22787 26404 22836 26432
rect 22787 26401 22799 26404
rect 22741 26395 22799 26401
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 26053 26435 26111 26441
rect 26053 26401 26065 26435
rect 26099 26432 26111 26435
rect 26418 26432 26424 26444
rect 26099 26404 26424 26432
rect 26099 26401 26111 26404
rect 26053 26395 26111 26401
rect 26418 26392 26424 26404
rect 26476 26392 26482 26444
rect 30558 26392 30564 26444
rect 30616 26432 30622 26444
rect 31110 26432 31116 26444
rect 30616 26404 31116 26432
rect 30616 26392 30622 26404
rect 31110 26392 31116 26404
rect 31168 26432 31174 26444
rect 31481 26435 31539 26441
rect 31481 26432 31493 26435
rect 31168 26404 31493 26432
rect 31168 26392 31174 26404
rect 31481 26401 31493 26404
rect 31527 26432 31539 26435
rect 33594 26432 33600 26444
rect 31527 26404 33600 26432
rect 31527 26401 31539 26404
rect 31481 26395 31539 26401
rect 33594 26392 33600 26404
rect 33652 26392 33658 26444
rect 34422 26392 34428 26444
rect 34480 26432 34486 26444
rect 35621 26435 35679 26441
rect 35621 26432 35633 26435
rect 34480 26404 35633 26432
rect 34480 26392 34486 26404
rect 35621 26401 35633 26404
rect 35667 26401 35679 26435
rect 35621 26395 35679 26401
rect 10870 26364 10876 26376
rect 9171 26336 10364 26364
rect 10831 26336 10876 26364
rect 9171 26333 9183 26336
rect 9125 26327 9183 26333
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 37642 26364 37648 26376
rect 32890 26336 37648 26364
rect 37642 26324 37648 26336
rect 37700 26324 37706 26376
rect 38286 26364 38292 26376
rect 38247 26336 38292 26364
rect 38286 26324 38292 26336
rect 38344 26324 38350 26376
rect 8294 26256 8300 26308
rect 8352 26296 8358 26308
rect 10965 26299 11023 26305
rect 10965 26296 10977 26299
rect 8352 26268 10977 26296
rect 8352 26256 8358 26268
rect 10965 26265 10977 26268
rect 11011 26265 11023 26299
rect 12710 26296 12716 26308
rect 12671 26268 12716 26296
rect 10965 26259 11023 26265
rect 12710 26256 12716 26268
rect 12768 26256 12774 26308
rect 12805 26299 12863 26305
rect 12805 26265 12817 26299
rect 12851 26296 12863 26299
rect 12851 26268 13676 26296
rect 12851 26265 12863 26268
rect 12805 26259 12863 26265
rect 5442 26228 5448 26240
rect 5403 26200 5448 26228
rect 5442 26188 5448 26200
rect 5500 26188 5506 26240
rect 13648 26228 13676 26268
rect 14826 26256 14832 26308
rect 14884 26296 14890 26308
rect 14884 26268 16422 26296
rect 14884 26256 14890 26268
rect 20346 26256 20352 26308
rect 20404 26296 20410 26308
rect 20993 26299 21051 26305
rect 20993 26296 21005 26299
rect 20404 26268 21005 26296
rect 20404 26256 20410 26268
rect 20993 26265 21005 26268
rect 21039 26265 21051 26299
rect 22554 26296 22560 26308
rect 22218 26268 22560 26296
rect 20993 26259 21051 26265
rect 22554 26256 22560 26268
rect 22612 26256 22618 26308
rect 26326 26296 26332 26308
rect 26287 26268 26332 26296
rect 26326 26256 26332 26268
rect 26384 26256 26390 26308
rect 29546 26296 29552 26308
rect 27554 26268 29552 26296
rect 29546 26256 29552 26268
rect 29604 26256 29610 26308
rect 31754 26256 31760 26308
rect 31812 26296 31818 26308
rect 31812 26268 31857 26296
rect 31812 26256 31818 26268
rect 34514 26256 34520 26308
rect 34572 26296 34578 26308
rect 34885 26299 34943 26305
rect 34885 26296 34897 26299
rect 34572 26268 34897 26296
rect 34572 26256 34578 26268
rect 34885 26265 34897 26268
rect 34931 26265 34943 26299
rect 34885 26259 34943 26265
rect 13814 26228 13820 26240
rect 13648 26200 13820 26228
rect 13814 26188 13820 26200
rect 13872 26188 13878 26240
rect 16758 26188 16764 26240
rect 16816 26228 16822 26240
rect 17405 26231 17463 26237
rect 17405 26228 17417 26231
rect 16816 26200 17417 26228
rect 16816 26188 16822 26200
rect 17405 26197 17417 26200
rect 17451 26197 17463 26231
rect 17405 26191 17463 26197
rect 25038 26188 25044 26240
rect 25096 26228 25102 26240
rect 25866 26228 25872 26240
rect 25096 26200 25872 26228
rect 25096 26188 25102 26200
rect 25866 26188 25872 26200
rect 25924 26188 25930 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 5258 25984 5264 26036
rect 5316 26024 5322 26036
rect 10962 26024 10968 26036
rect 5316 25996 10968 26024
rect 5316 25984 5322 25996
rect 10962 25984 10968 25996
rect 11020 25984 11026 26036
rect 11698 25984 11704 26036
rect 11756 26024 11762 26036
rect 11793 26027 11851 26033
rect 11793 26024 11805 26027
rect 11756 25996 11805 26024
rect 11756 25984 11762 25996
rect 11793 25993 11805 25996
rect 11839 25993 11851 26027
rect 13814 26024 13820 26036
rect 13775 25996 13820 26024
rect 11793 25987 11851 25993
rect 13814 25984 13820 25996
rect 13872 25984 13878 26036
rect 15930 25984 15936 26036
rect 15988 26024 15994 26036
rect 20162 26024 20168 26036
rect 15988 25996 20168 26024
rect 15988 25984 15994 25996
rect 20162 25984 20168 25996
rect 20220 25984 20226 26036
rect 26602 26024 26608 26036
rect 24780 25996 26608 26024
rect 9493 25959 9551 25965
rect 9493 25925 9505 25959
rect 9539 25956 9551 25959
rect 10229 25959 10287 25965
rect 10229 25956 10241 25959
rect 9539 25928 10241 25956
rect 9539 25925 9551 25928
rect 9493 25919 9551 25925
rect 10229 25925 10241 25928
rect 10275 25925 10287 25959
rect 10229 25919 10287 25925
rect 19058 25916 19064 25968
rect 19116 25956 19122 25968
rect 24670 25956 24676 25968
rect 19116 25928 20378 25956
rect 24426 25928 24676 25956
rect 19116 25916 19122 25928
rect 24670 25916 24676 25928
rect 24728 25916 24734 25968
rect 5353 25891 5411 25897
rect 5353 25857 5365 25891
rect 5399 25888 5411 25891
rect 5442 25888 5448 25900
rect 5399 25860 5448 25888
rect 5399 25857 5411 25860
rect 5353 25851 5411 25857
rect 5442 25848 5448 25860
rect 5500 25848 5506 25900
rect 7098 25848 7104 25900
rect 7156 25888 7162 25900
rect 7469 25891 7527 25897
rect 7469 25888 7481 25891
rect 7156 25860 7481 25888
rect 7156 25848 7162 25860
rect 7469 25857 7481 25860
rect 7515 25857 7527 25891
rect 9398 25888 9404 25900
rect 9359 25860 9404 25888
rect 7469 25851 7527 25857
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25888 11759 25891
rect 13725 25891 13783 25897
rect 11747 25860 13676 25888
rect 11747 25857 11759 25860
rect 11701 25851 11759 25857
rect 5534 25820 5540 25832
rect 5495 25792 5540 25820
rect 5534 25780 5540 25792
rect 5592 25780 5598 25832
rect 8757 25823 8815 25829
rect 8757 25789 8769 25823
rect 8803 25820 8815 25823
rect 9214 25820 9220 25832
rect 8803 25792 9220 25820
rect 8803 25789 8815 25792
rect 8757 25783 8815 25789
rect 9214 25780 9220 25792
rect 9272 25780 9278 25832
rect 9674 25780 9680 25832
rect 9732 25820 9738 25832
rect 10137 25823 10195 25829
rect 10137 25820 10149 25823
rect 9732 25792 10149 25820
rect 9732 25780 9738 25792
rect 10137 25789 10149 25792
rect 10183 25789 10195 25823
rect 10137 25783 10195 25789
rect 10781 25823 10839 25829
rect 10781 25789 10793 25823
rect 10827 25820 10839 25823
rect 10827 25792 10916 25820
rect 10827 25789 10839 25792
rect 10781 25783 10839 25789
rect 10888 25764 10916 25792
rect 10870 25712 10876 25764
rect 10928 25712 10934 25764
rect 5994 25684 6000 25696
rect 5955 25656 6000 25684
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 7558 25684 7564 25696
rect 7519 25656 7564 25684
rect 7558 25644 7564 25656
rect 7616 25644 7622 25696
rect 7834 25644 7840 25696
rect 7892 25684 7898 25696
rect 11716 25684 11744 25851
rect 13648 25820 13676 25860
rect 13725 25857 13737 25891
rect 13771 25888 13783 25891
rect 14274 25888 14280 25900
rect 13771 25860 14280 25888
rect 13771 25857 13783 25860
rect 13725 25851 13783 25857
rect 14274 25848 14280 25860
rect 14332 25848 14338 25900
rect 15286 25820 15292 25832
rect 13648 25792 15292 25820
rect 15286 25780 15292 25792
rect 15344 25780 15350 25832
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 19484 25792 19625 25820
rect 19484 25780 19490 25792
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19889 25823 19947 25829
rect 19889 25820 19901 25823
rect 19613 25783 19671 25789
rect 19720 25792 19901 25820
rect 19518 25712 19524 25764
rect 19576 25752 19582 25764
rect 19720 25752 19748 25792
rect 19889 25789 19901 25792
rect 19935 25789 19947 25823
rect 22922 25820 22928 25832
rect 22883 25792 22928 25820
rect 19889 25783 19947 25789
rect 22922 25780 22928 25792
rect 22980 25780 22986 25832
rect 23198 25820 23204 25832
rect 23159 25792 23204 25820
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 24673 25823 24731 25829
rect 24673 25789 24685 25823
rect 24719 25820 24731 25823
rect 24780 25820 24808 25996
rect 26602 25984 26608 25996
rect 26660 26024 26666 26036
rect 37734 26024 37740 26036
rect 26660 25996 29684 26024
rect 37695 25996 37740 26024
rect 26660 25984 26666 25996
rect 28074 25916 28080 25968
rect 28132 25916 28138 25968
rect 29656 25965 29684 25996
rect 37734 25984 37740 25996
rect 37792 25984 37798 26036
rect 29641 25959 29699 25965
rect 29641 25925 29653 25959
rect 29687 25925 29699 25959
rect 29641 25919 29699 25925
rect 33870 25916 33876 25968
rect 33928 25956 33934 25968
rect 33965 25959 34023 25965
rect 33965 25956 33977 25959
rect 33928 25928 33977 25956
rect 33928 25916 33934 25928
rect 33965 25925 33977 25928
rect 34011 25925 34023 25959
rect 35710 25956 35716 25968
rect 35190 25928 35716 25956
rect 33965 25919 34023 25925
rect 35710 25916 35716 25928
rect 35768 25916 35774 25968
rect 26418 25848 26424 25900
rect 26476 25888 26482 25900
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 26476 25860 27169 25888
rect 26476 25848 26482 25860
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 29362 25888 29368 25900
rect 29323 25860 29368 25888
rect 27157 25851 27215 25857
rect 29362 25848 29368 25860
rect 29420 25848 29426 25900
rect 30742 25848 30748 25900
rect 30800 25848 30806 25900
rect 33594 25848 33600 25900
rect 33652 25888 33658 25900
rect 33689 25891 33747 25897
rect 33689 25888 33701 25891
rect 33652 25860 33701 25888
rect 33652 25848 33658 25860
rect 33689 25857 33701 25860
rect 33735 25857 33747 25891
rect 33689 25851 33747 25857
rect 37921 25891 37979 25897
rect 37921 25857 37933 25891
rect 37967 25888 37979 25891
rect 38654 25888 38660 25900
rect 37967 25860 38660 25888
rect 37967 25857 37979 25860
rect 37921 25851 37979 25857
rect 38654 25848 38660 25860
rect 38712 25848 38718 25900
rect 24719 25792 24808 25820
rect 24719 25789 24731 25792
rect 24673 25783 24731 25789
rect 24854 25780 24860 25832
rect 24912 25820 24918 25832
rect 27433 25823 27491 25829
rect 27433 25820 27445 25823
rect 24912 25792 27445 25820
rect 24912 25780 24918 25792
rect 27433 25789 27445 25792
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 35713 25823 35771 25829
rect 35713 25789 35725 25823
rect 35759 25789 35771 25823
rect 35713 25783 35771 25789
rect 19576 25724 19748 25752
rect 19576 25712 19582 25724
rect 28534 25712 28540 25764
rect 28592 25752 28598 25764
rect 28592 25724 29040 25752
rect 28592 25712 28598 25724
rect 7892 25656 11744 25684
rect 7892 25644 7898 25656
rect 14366 25644 14372 25696
rect 14424 25684 14430 25696
rect 19242 25684 19248 25696
rect 14424 25656 19248 25684
rect 14424 25644 14430 25656
rect 19242 25644 19248 25656
rect 19300 25644 19306 25696
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 21361 25687 21419 25693
rect 21361 25684 21373 25687
rect 21048 25656 21373 25684
rect 21048 25644 21054 25656
rect 21361 25653 21373 25656
rect 21407 25653 21419 25687
rect 21361 25647 21419 25653
rect 27430 25644 27436 25696
rect 27488 25684 27494 25696
rect 28905 25687 28963 25693
rect 28905 25684 28917 25687
rect 27488 25656 28917 25684
rect 27488 25644 27494 25656
rect 28905 25653 28917 25656
rect 28951 25653 28963 25687
rect 29012 25684 29040 25724
rect 30668 25724 31754 25752
rect 30668 25684 30696 25724
rect 29012 25656 30696 25684
rect 28905 25647 28963 25653
rect 30834 25644 30840 25696
rect 30892 25684 30898 25696
rect 31113 25687 31171 25693
rect 31113 25684 31125 25687
rect 30892 25656 31125 25684
rect 30892 25644 30898 25656
rect 31113 25653 31125 25656
rect 31159 25653 31171 25687
rect 31726 25684 31754 25724
rect 35728 25684 35756 25783
rect 31726 25656 35756 25684
rect 31113 25647 31171 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 7926 25480 7932 25492
rect 7887 25452 7932 25480
rect 7926 25440 7932 25452
rect 7984 25440 7990 25492
rect 9398 25440 9404 25492
rect 9456 25480 9462 25492
rect 17037 25483 17095 25489
rect 9456 25452 16988 25480
rect 9456 25440 9462 25452
rect 16960 25412 16988 25452
rect 17037 25449 17049 25483
rect 17083 25480 17095 25483
rect 21634 25480 21640 25492
rect 17083 25452 21640 25480
rect 17083 25449 17095 25452
rect 17037 25443 17095 25449
rect 21634 25440 21640 25452
rect 21692 25440 21698 25492
rect 22360 25483 22418 25489
rect 22360 25449 22372 25483
rect 22406 25480 22418 25483
rect 22830 25480 22836 25492
rect 22406 25452 22836 25480
rect 22406 25449 22418 25452
rect 22360 25443 22418 25449
rect 22830 25440 22836 25452
rect 22888 25480 22894 25492
rect 26881 25483 26939 25489
rect 26881 25480 26893 25483
rect 22888 25452 26893 25480
rect 22888 25440 22894 25452
rect 26881 25449 26893 25452
rect 26927 25449 26939 25483
rect 26881 25443 26939 25449
rect 30374 25440 30380 25492
rect 30432 25480 30438 25492
rect 32309 25483 32367 25489
rect 32309 25480 32321 25483
rect 30432 25452 32321 25480
rect 30432 25440 30438 25452
rect 32309 25449 32321 25452
rect 32355 25449 32367 25483
rect 32309 25443 32367 25449
rect 35342 25440 35348 25492
rect 35400 25480 35406 25492
rect 37185 25483 37243 25489
rect 37185 25480 37197 25483
rect 35400 25452 37197 25480
rect 35400 25440 35406 25452
rect 37185 25449 37197 25452
rect 37231 25449 37243 25483
rect 37185 25443 37243 25449
rect 20254 25412 20260 25424
rect 16960 25384 20260 25412
rect 20254 25372 20260 25384
rect 20312 25372 20318 25424
rect 22112 25384 22232 25412
rect 2866 25304 2872 25356
rect 2924 25344 2930 25356
rect 4893 25347 4951 25353
rect 4893 25344 4905 25347
rect 2924 25316 4905 25344
rect 2924 25304 2930 25316
rect 4893 25313 4905 25316
rect 4939 25313 4951 25347
rect 4893 25307 4951 25313
rect 7285 25347 7343 25353
rect 7285 25313 7297 25347
rect 7331 25344 7343 25347
rect 8018 25344 8024 25356
rect 7331 25316 8024 25344
rect 7331 25313 7343 25316
rect 7285 25307 7343 25313
rect 8018 25304 8024 25316
rect 8076 25304 8082 25356
rect 9214 25344 9220 25356
rect 9175 25316 9220 25344
rect 9214 25304 9220 25316
rect 9272 25304 9278 25356
rect 10962 25304 10968 25356
rect 11020 25344 11026 25356
rect 22112 25344 22140 25384
rect 11020 25316 22140 25344
rect 22204 25344 22232 25384
rect 25038 25344 25044 25356
rect 22204 25316 25044 25344
rect 11020 25304 11026 25316
rect 5074 25276 5080 25288
rect 5035 25248 5080 25276
rect 5074 25236 5080 25248
rect 5132 25236 5138 25288
rect 7469 25279 7527 25285
rect 7469 25245 7481 25279
rect 7515 25276 7527 25279
rect 8294 25276 8300 25288
rect 7515 25248 8300 25276
rect 7515 25245 7527 25248
rect 7469 25239 7527 25245
rect 8294 25236 8300 25248
rect 8352 25236 8358 25288
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 14366 25276 14372 25288
rect 10459 25248 14372 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 14366 25236 14372 25248
rect 14424 25236 14430 25288
rect 14660 25285 14688 25316
rect 25038 25304 25044 25316
rect 25096 25304 25102 25356
rect 25133 25347 25191 25353
rect 25133 25313 25145 25347
rect 25179 25344 25191 25347
rect 26418 25344 26424 25356
rect 25179 25316 26424 25344
rect 25179 25313 25191 25316
rect 25133 25307 25191 25313
rect 26418 25304 26424 25316
rect 26476 25304 26482 25356
rect 30558 25344 30564 25356
rect 30519 25316 30564 25344
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 34698 25304 34704 25356
rect 34756 25344 34762 25356
rect 35161 25347 35219 25353
rect 35161 25344 35173 25347
rect 34756 25316 35173 25344
rect 34756 25304 34762 25316
rect 35161 25313 35173 25316
rect 35207 25313 35219 25347
rect 35161 25307 35219 25313
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25245 14703 25279
rect 14645 25239 14703 25245
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25245 15347 25279
rect 15289 25239 15347 25245
rect 9309 25211 9367 25217
rect 9309 25177 9321 25211
rect 9355 25177 9367 25211
rect 9858 25208 9864 25220
rect 9819 25180 9864 25208
rect 9309 25171 9367 25177
rect 5537 25143 5595 25149
rect 5537 25109 5549 25143
rect 5583 25140 5595 25143
rect 5626 25140 5632 25152
rect 5583 25112 5632 25140
rect 5583 25109 5595 25112
rect 5537 25103 5595 25109
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 9324 25140 9352 25171
rect 9858 25168 9864 25180
rect 9916 25168 9922 25220
rect 10505 25143 10563 25149
rect 10505 25140 10517 25143
rect 9324 25112 10517 25140
rect 10505 25109 10517 25112
rect 10551 25109 10563 25143
rect 14734 25140 14740 25152
rect 14695 25112 14740 25140
rect 10505 25103 10563 25109
rect 14734 25100 14740 25112
rect 14792 25100 14798 25152
rect 15304 25140 15332 25239
rect 16850 25236 16856 25288
rect 16908 25276 16914 25288
rect 17681 25279 17739 25285
rect 17681 25276 17693 25279
rect 16908 25248 17693 25276
rect 16908 25236 16914 25248
rect 17681 25245 17693 25248
rect 17727 25245 17739 25279
rect 22086 25279 22144 25285
rect 22086 25276 22098 25279
rect 17681 25239 17739 25245
rect 22066 25245 22098 25276
rect 22132 25245 22144 25279
rect 22066 25239 22144 25245
rect 15565 25211 15623 25217
rect 15565 25177 15577 25211
rect 15611 25208 15623 25211
rect 16942 25208 16948 25220
rect 15611 25180 15976 25208
rect 16790 25180 16948 25208
rect 15611 25177 15623 25180
rect 15565 25171 15623 25177
rect 15746 25140 15752 25152
rect 15304 25112 15752 25140
rect 15746 25100 15752 25112
rect 15804 25100 15810 25152
rect 15948 25140 15976 25180
rect 16942 25168 16948 25180
rect 17000 25168 17006 25220
rect 18138 25168 18144 25220
rect 18196 25208 18202 25220
rect 18417 25211 18475 25217
rect 18417 25208 18429 25211
rect 18196 25180 18429 25208
rect 18196 25168 18202 25180
rect 18417 25177 18429 25180
rect 18463 25177 18475 25211
rect 22066 25208 22094 25239
rect 34606 25236 34612 25288
rect 34664 25276 34670 25288
rect 34885 25279 34943 25285
rect 34885 25276 34897 25279
rect 34664 25248 34897 25276
rect 34664 25236 34670 25248
rect 34885 25245 34897 25248
rect 34931 25245 34943 25279
rect 37090 25276 37096 25288
rect 37051 25248 37096 25276
rect 34885 25239 34943 25245
rect 37090 25236 37096 25248
rect 37148 25236 37154 25288
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 22278 25208 22284 25220
rect 22066 25180 22284 25208
rect 18417 25171 18475 25177
rect 22278 25168 22284 25180
rect 22336 25168 22342 25220
rect 24946 25208 24952 25220
rect 23598 25180 24952 25208
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 25038 25168 25044 25220
rect 25096 25208 25102 25220
rect 25406 25208 25412 25220
rect 25096 25180 25412 25208
rect 25096 25168 25102 25180
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 27522 25208 27528 25220
rect 26634 25180 27528 25208
rect 27522 25168 27528 25180
rect 27580 25168 27586 25220
rect 30834 25208 30840 25220
rect 30795 25180 30840 25208
rect 30834 25168 30840 25180
rect 30892 25168 30898 25220
rect 31846 25168 31852 25220
rect 31904 25168 31910 25220
rect 36170 25168 36176 25220
rect 36228 25168 36234 25220
rect 16850 25140 16856 25152
rect 15948 25112 16856 25140
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 21174 25100 21180 25152
rect 21232 25140 21238 25152
rect 21358 25140 21364 25152
rect 21232 25112 21364 25140
rect 21232 25100 21238 25112
rect 21358 25100 21364 25112
rect 21416 25100 21422 25152
rect 23845 25143 23903 25149
rect 23845 25109 23857 25143
rect 23891 25140 23903 25143
rect 25590 25140 25596 25152
rect 23891 25112 25596 25140
rect 23891 25109 23903 25112
rect 23845 25103 23903 25109
rect 25590 25100 25596 25112
rect 25648 25100 25654 25152
rect 35342 25100 35348 25152
rect 35400 25140 35406 25152
rect 36633 25143 36691 25149
rect 36633 25140 36645 25143
rect 35400 25112 36645 25140
rect 35400 25100 35406 25112
rect 36633 25109 36645 25112
rect 36679 25109 36691 25143
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 36633 25103 36691 25109
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 5074 24896 5080 24948
rect 5132 24936 5138 24948
rect 5261 24939 5319 24945
rect 5261 24936 5273 24939
rect 5132 24908 5273 24936
rect 5132 24896 5138 24908
rect 5261 24905 5273 24908
rect 5307 24905 5319 24939
rect 5261 24899 5319 24905
rect 16298 24896 16304 24948
rect 16356 24936 16362 24948
rect 18690 24936 18696 24948
rect 16356 24908 18696 24936
rect 16356 24896 16362 24908
rect 18690 24896 18696 24908
rect 18748 24896 18754 24948
rect 23842 24896 23848 24948
rect 23900 24936 23906 24948
rect 38010 24936 38016 24948
rect 23900 24908 38016 24936
rect 23900 24896 23906 24908
rect 38010 24896 38016 24908
rect 38068 24896 38074 24948
rect 10229 24871 10287 24877
rect 10229 24868 10241 24871
rect 9968 24840 10241 24868
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 3970 24800 3976 24812
rect 1627 24772 3976 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 3970 24760 3976 24772
rect 4028 24760 4034 24812
rect 4065 24803 4123 24809
rect 4065 24769 4077 24803
rect 4111 24800 4123 24803
rect 4614 24800 4620 24812
rect 4111 24772 4620 24800
rect 4111 24769 4123 24772
rect 4065 24763 4123 24769
rect 4614 24760 4620 24772
rect 4672 24760 4678 24812
rect 4709 24803 4767 24809
rect 4709 24769 4721 24803
rect 4755 24769 4767 24803
rect 4709 24763 4767 24769
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24769 5227 24803
rect 5810 24800 5816 24812
rect 5771 24772 5816 24800
rect 5169 24763 5227 24769
rect 4724 24732 4752 24763
rect 3896 24704 4752 24732
rect 5184 24732 5212 24763
rect 5810 24760 5816 24772
rect 5868 24760 5874 24812
rect 6822 24800 6828 24812
rect 6783 24772 6828 24800
rect 6822 24760 6828 24772
rect 6880 24760 6886 24812
rect 7009 24803 7067 24809
rect 7009 24769 7021 24803
rect 7055 24800 7067 24803
rect 7558 24800 7564 24812
rect 7055 24772 7564 24800
rect 7055 24769 7067 24772
rect 7009 24763 7067 24769
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 7926 24800 7932 24812
rect 7800 24772 7932 24800
rect 7800 24760 7806 24772
rect 7926 24760 7932 24772
rect 7984 24760 7990 24812
rect 9122 24760 9128 24812
rect 9180 24800 9186 24812
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 9180 24772 9413 24800
rect 9180 24760 9186 24772
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 9401 24763 9459 24769
rect 9493 24803 9551 24809
rect 9493 24769 9505 24803
rect 9539 24800 9551 24803
rect 9968 24800 9996 24840
rect 10229 24837 10241 24840
rect 10275 24837 10287 24871
rect 10229 24831 10287 24837
rect 12161 24871 12219 24877
rect 12161 24837 12173 24871
rect 12207 24868 12219 24871
rect 18322 24868 18328 24880
rect 12207 24840 12756 24868
rect 12207 24837 12219 24840
rect 12161 24831 12219 24837
rect 9539 24772 9996 24800
rect 9539 24769 9551 24772
rect 9493 24763 9551 24769
rect 8570 24732 8576 24744
rect 5184 24704 8576 24732
rect 3896 24673 3924 24704
rect 8570 24692 8576 24704
rect 8628 24692 8634 24744
rect 10137 24735 10195 24741
rect 10137 24701 10149 24735
rect 10183 24732 10195 24735
rect 10226 24732 10232 24744
rect 10183 24704 10232 24732
rect 10183 24701 10195 24704
rect 10137 24695 10195 24701
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 11146 24732 11152 24744
rect 11107 24704 11152 24732
rect 11146 24692 11152 24704
rect 11204 24732 11210 24744
rect 12069 24735 12127 24741
rect 12069 24732 12081 24735
rect 11204 24704 12081 24732
rect 11204 24692 11210 24704
rect 12069 24701 12081 24704
rect 12115 24701 12127 24735
rect 12728 24732 12756 24840
rect 17972 24840 18328 24868
rect 13173 24803 13231 24809
rect 13173 24769 13185 24803
rect 13219 24800 13231 24803
rect 17972 24800 18000 24840
rect 18322 24828 18328 24840
rect 18380 24828 18386 24880
rect 22833 24871 22891 24877
rect 22833 24837 22845 24871
rect 22879 24868 22891 24871
rect 22922 24868 22928 24880
rect 22879 24840 22928 24868
rect 22879 24837 22891 24840
rect 22833 24831 22891 24837
rect 22922 24828 22928 24840
rect 22980 24828 22986 24880
rect 36446 24868 36452 24880
rect 34822 24840 36452 24868
rect 36446 24828 36452 24840
rect 36504 24828 36510 24880
rect 18138 24800 18144 24812
rect 13219 24772 18000 24800
rect 18099 24772 18144 24800
rect 13219 24769 13231 24772
rect 13173 24763 13231 24769
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 19518 24760 19524 24812
rect 19576 24760 19582 24812
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24800 22063 24803
rect 29822 24800 29828 24812
rect 22051 24772 22784 24800
rect 29670 24772 29828 24800
rect 22051 24769 22063 24772
rect 22005 24763 22063 24769
rect 13265 24735 13323 24741
rect 13265 24732 13277 24735
rect 12728 24704 13277 24732
rect 12069 24695 12127 24701
rect 13265 24701 13277 24704
rect 13311 24701 13323 24735
rect 13265 24695 13323 24701
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 18414 24732 18420 24744
rect 15620 24704 18420 24732
rect 15620 24692 15626 24704
rect 18414 24692 18420 24704
rect 18472 24692 18478 24744
rect 19426 24692 19432 24744
rect 19484 24732 19490 24744
rect 22756 24732 22784 24772
rect 29822 24760 29828 24772
rect 29880 24760 29886 24812
rect 27614 24732 27620 24744
rect 19484 24704 22094 24732
rect 22756 24704 27620 24732
rect 19484 24692 19490 24704
rect 3881 24667 3939 24673
rect 3881 24633 3893 24667
rect 3927 24633 3939 24667
rect 3881 24627 3939 24633
rect 4525 24667 4583 24673
rect 4525 24633 4537 24667
rect 4571 24664 4583 24667
rect 5534 24664 5540 24676
rect 4571 24636 5540 24664
rect 4571 24633 4583 24636
rect 4525 24627 4583 24633
rect 5534 24624 5540 24636
rect 5592 24624 5598 24676
rect 5994 24624 6000 24676
rect 6052 24664 6058 24676
rect 7193 24667 7251 24673
rect 7193 24664 7205 24667
rect 6052 24636 7205 24664
rect 6052 24624 6058 24636
rect 7193 24633 7205 24636
rect 7239 24633 7251 24667
rect 7193 24627 7251 24633
rect 9858 24624 9864 24676
rect 9916 24664 9922 24676
rect 12621 24667 12679 24673
rect 12621 24664 12633 24667
rect 9916 24636 12633 24664
rect 9916 24624 9922 24636
rect 12621 24633 12633 24636
rect 12667 24664 12679 24667
rect 13170 24664 13176 24676
rect 12667 24636 13176 24664
rect 12667 24633 12679 24636
rect 12621 24627 12679 24633
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 14550 24624 14556 24676
rect 14608 24664 14614 24676
rect 20070 24664 20076 24676
rect 14608 24636 18276 24664
rect 14608 24624 14614 24636
rect 1762 24596 1768 24608
rect 1723 24568 1768 24596
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 5905 24599 5963 24605
rect 5905 24565 5917 24599
rect 5951 24596 5963 24599
rect 6730 24596 6736 24608
rect 5951 24568 6736 24596
rect 5951 24565 5963 24568
rect 5905 24559 5963 24565
rect 6730 24556 6736 24568
rect 6788 24556 6794 24608
rect 8018 24596 8024 24608
rect 7979 24568 8024 24596
rect 8018 24556 8024 24568
rect 8076 24556 8082 24608
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 18046 24596 18052 24608
rect 15896 24568 18052 24596
rect 15896 24556 15902 24568
rect 18046 24556 18052 24568
rect 18104 24556 18110 24608
rect 18248 24596 18276 24636
rect 19812 24636 20076 24664
rect 19812 24596 19840 24636
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 22066 24664 22094 24704
rect 27614 24692 27620 24704
rect 27672 24692 27678 24744
rect 28261 24735 28319 24741
rect 28261 24701 28273 24735
rect 28307 24701 28319 24735
rect 28534 24732 28540 24744
rect 28495 24704 28540 24732
rect 28261 24695 28319 24701
rect 22278 24664 22284 24676
rect 22066 24636 22284 24664
rect 22278 24624 22284 24636
rect 22336 24664 22342 24676
rect 22922 24664 22928 24676
rect 22336 24636 22928 24664
rect 22336 24624 22342 24636
rect 22922 24624 22928 24636
rect 22980 24624 22986 24676
rect 18248 24568 19840 24596
rect 19889 24599 19947 24605
rect 19889 24565 19901 24599
rect 19935 24596 19947 24599
rect 20162 24596 20168 24608
rect 19935 24568 20168 24596
rect 19935 24565 19947 24568
rect 19889 24559 19947 24565
rect 20162 24556 20168 24568
rect 20220 24556 20226 24608
rect 28276 24596 28304 24695
rect 28534 24692 28540 24704
rect 28592 24692 28598 24744
rect 31938 24692 31944 24744
rect 31996 24732 32002 24744
rect 33042 24732 33048 24744
rect 31996 24704 33048 24732
rect 31996 24692 32002 24704
rect 33042 24692 33048 24704
rect 33100 24732 33106 24744
rect 33321 24735 33379 24741
rect 33321 24732 33333 24735
rect 33100 24704 33333 24732
rect 33100 24692 33106 24704
rect 33321 24701 33333 24704
rect 33367 24701 33379 24735
rect 33321 24695 33379 24701
rect 33597 24735 33655 24741
rect 33597 24701 33609 24735
rect 33643 24732 33655 24735
rect 33962 24732 33968 24744
rect 33643 24704 33968 24732
rect 33643 24701 33655 24704
rect 33597 24695 33655 24701
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 35345 24735 35403 24741
rect 35345 24701 35357 24735
rect 35391 24701 35403 24735
rect 35345 24695 35403 24701
rect 29638 24624 29644 24676
rect 29696 24664 29702 24676
rect 29696 24636 31754 24664
rect 29696 24624 29702 24636
rect 28994 24596 29000 24608
rect 28276 24568 29000 24596
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 30006 24596 30012 24608
rect 29967 24568 30012 24596
rect 30006 24556 30012 24568
rect 30064 24556 30070 24608
rect 31726 24596 31754 24636
rect 35360 24596 35388 24695
rect 31726 24568 35388 24596
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 15838 24392 15844 24404
rect 8628 24364 15844 24392
rect 8628 24352 8634 24364
rect 15838 24352 15844 24364
rect 15896 24352 15902 24404
rect 16022 24401 16028 24404
rect 16012 24395 16028 24401
rect 16012 24392 16024 24395
rect 15935 24364 16024 24392
rect 16012 24361 16024 24364
rect 16080 24392 16086 24404
rect 16080 24364 17908 24392
rect 16012 24355 16028 24361
rect 16022 24352 16028 24355
rect 16080 24352 16086 24364
rect 8386 24324 8392 24336
rect 2746 24296 8392 24324
rect 1857 24259 1915 24265
rect 1857 24225 1869 24259
rect 1903 24256 1915 24259
rect 2746 24256 2774 24296
rect 8386 24284 8392 24296
rect 8444 24284 8450 24336
rect 17880 24324 17908 24364
rect 18414 24352 18420 24404
rect 18472 24392 18478 24404
rect 21177 24395 21235 24401
rect 21177 24392 21189 24395
rect 18472 24364 21189 24392
rect 18472 24352 18478 24364
rect 21177 24361 21189 24364
rect 21223 24361 21235 24395
rect 21177 24355 21235 24361
rect 26510 24352 26516 24404
rect 26568 24392 26574 24404
rect 30006 24392 30012 24404
rect 26568 24364 30012 24392
rect 26568 24352 26574 24364
rect 30006 24352 30012 24364
rect 30064 24352 30070 24404
rect 34422 24352 34428 24404
rect 34480 24392 34486 24404
rect 35802 24392 35808 24404
rect 34480 24364 35808 24392
rect 34480 24352 34486 24364
rect 35802 24352 35808 24364
rect 35860 24352 35866 24404
rect 18690 24324 18696 24336
rect 17880 24296 18696 24324
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 26694 24284 26700 24336
rect 26752 24324 26758 24336
rect 29638 24324 29644 24336
rect 26752 24296 29644 24324
rect 26752 24284 26758 24296
rect 29638 24284 29644 24296
rect 29696 24284 29702 24336
rect 1903 24228 2774 24256
rect 1903 24225 1915 24228
rect 1857 24219 1915 24225
rect 5810 24216 5816 24268
rect 5868 24256 5874 24268
rect 6825 24259 6883 24265
rect 6825 24256 6837 24259
rect 5868 24228 6837 24256
rect 5868 24216 5874 24228
rect 6825 24225 6837 24228
rect 6871 24256 6883 24259
rect 9858 24256 9864 24268
rect 6871 24228 9864 24256
rect 6871 24225 6883 24228
rect 6825 24219 6883 24225
rect 9858 24216 9864 24228
rect 9916 24216 9922 24268
rect 10778 24216 10784 24268
rect 10836 24256 10842 24268
rect 12437 24259 12495 24265
rect 12437 24256 12449 24259
rect 10836 24228 12449 24256
rect 10836 24216 10842 24228
rect 12437 24225 12449 24228
rect 12483 24225 12495 24259
rect 19426 24256 19432 24268
rect 19387 24228 19432 24256
rect 12437 24219 12495 24225
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 27614 24216 27620 24268
rect 27672 24256 27678 24268
rect 27672 24228 31754 24256
rect 27672 24216 27678 24228
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 7282 24188 7288 24200
rect 7243 24160 7288 24188
rect 7282 24148 7288 24160
rect 7340 24148 7346 24200
rect 9769 24191 9827 24197
rect 9769 24157 9781 24191
rect 9815 24188 9827 24191
rect 10134 24188 10140 24200
rect 9815 24160 10140 24188
rect 9815 24157 9827 24160
rect 9769 24151 9827 24157
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 13265 24191 13323 24197
rect 13265 24157 13277 24191
rect 13311 24188 13323 24191
rect 15562 24188 15568 24200
rect 13311 24160 15568 24188
rect 13311 24157 13323 24160
rect 13265 24151 13323 24157
rect 15562 24148 15568 24160
rect 15620 24148 15626 24200
rect 15746 24188 15752 24200
rect 15707 24160 15752 24188
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 20806 24148 20812 24200
rect 20864 24148 20870 24200
rect 28276 24197 28304 24228
rect 28261 24191 28319 24197
rect 28261 24157 28273 24191
rect 28307 24157 28319 24191
rect 28261 24151 28319 24157
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24157 29791 24191
rect 31726 24188 31754 24228
rect 33042 24216 33048 24268
rect 33100 24256 33106 24268
rect 34149 24259 34207 24265
rect 34149 24256 34161 24259
rect 33100 24228 34161 24256
rect 33100 24216 33106 24228
rect 34149 24225 34161 24228
rect 34195 24256 34207 24259
rect 34606 24256 34612 24268
rect 34195 24228 34612 24256
rect 34195 24225 34207 24228
rect 34149 24219 34207 24225
rect 34606 24216 34612 24228
rect 34664 24256 34670 24268
rect 34885 24259 34943 24265
rect 34885 24256 34897 24259
rect 34664 24228 34897 24256
rect 34664 24216 34670 24228
rect 34885 24225 34897 24228
rect 34931 24225 34943 24259
rect 34885 24219 34943 24225
rect 35161 24259 35219 24265
rect 35161 24225 35173 24259
rect 35207 24256 35219 24259
rect 35250 24256 35256 24268
rect 35207 24228 35256 24256
rect 35207 24225 35219 24228
rect 35161 24219 35219 24225
rect 35250 24216 35256 24228
rect 35308 24216 35314 24268
rect 33413 24191 33471 24197
rect 33413 24188 33425 24191
rect 31726 24160 33425 24188
rect 29733 24151 29791 24157
rect 33413 24157 33425 24160
rect 33459 24188 33471 24191
rect 34514 24188 34520 24200
rect 33459 24160 34520 24188
rect 33459 24157 33471 24160
rect 33413 24151 33471 24157
rect 4890 24080 4896 24132
rect 4948 24120 4954 24132
rect 6181 24123 6239 24129
rect 6181 24120 6193 24123
rect 4948 24092 6193 24120
rect 4948 24080 4954 24092
rect 6181 24089 6193 24092
rect 6227 24089 6239 24123
rect 6181 24083 6239 24089
rect 6270 24080 6276 24132
rect 6328 24120 6334 24132
rect 7377 24123 7435 24129
rect 6328 24092 6373 24120
rect 6328 24080 6334 24092
rect 7377 24089 7389 24123
rect 7423 24120 7435 24123
rect 9490 24120 9496 24132
rect 7423 24092 9496 24120
rect 7423 24089 7435 24092
rect 7377 24083 7435 24089
rect 9490 24080 9496 24092
rect 9548 24080 9554 24132
rect 11974 24080 11980 24132
rect 12032 24120 12038 24132
rect 12161 24123 12219 24129
rect 12161 24120 12173 24123
rect 12032 24092 12173 24120
rect 12032 24080 12038 24092
rect 12161 24089 12173 24092
rect 12207 24089 12219 24123
rect 12161 24083 12219 24089
rect 12250 24080 12256 24132
rect 12308 24120 12314 24132
rect 12308 24092 12353 24120
rect 12406 24092 13492 24120
rect 12308 24080 12314 24092
rect 8294 24012 8300 24064
rect 8352 24052 8358 24064
rect 9861 24055 9919 24061
rect 9861 24052 9873 24055
rect 8352 24024 9873 24052
rect 8352 24012 8358 24024
rect 9861 24021 9873 24024
rect 9907 24021 9919 24055
rect 9861 24015 9919 24021
rect 10778 24012 10784 24064
rect 10836 24052 10842 24064
rect 12406 24052 12434 24092
rect 13354 24052 13360 24064
rect 10836 24024 12434 24052
rect 13315 24024 13360 24052
rect 10836 24012 10842 24024
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 13464 24052 13492 24092
rect 14366 24080 14372 24132
rect 14424 24120 14430 24132
rect 16298 24120 16304 24132
rect 14424 24092 16304 24120
rect 14424 24080 14430 24092
rect 16298 24080 16304 24092
rect 16356 24080 16362 24132
rect 17678 24120 17684 24132
rect 17250 24092 17684 24120
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 17773 24123 17831 24129
rect 17773 24089 17785 24123
rect 17819 24120 17831 24123
rect 18322 24120 18328 24132
rect 17819 24092 18328 24120
rect 17819 24089 17831 24092
rect 17773 24083 17831 24089
rect 18322 24080 18328 24092
rect 18380 24080 18386 24132
rect 19705 24123 19763 24129
rect 19705 24120 19717 24123
rect 18432 24092 19717 24120
rect 16666 24052 16672 24064
rect 13464 24024 16672 24052
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 17494 24012 17500 24064
rect 17552 24052 17558 24064
rect 18432 24052 18460 24092
rect 19705 24089 19717 24092
rect 19751 24089 19763 24123
rect 28994 24120 29000 24132
rect 28955 24092 29000 24120
rect 19705 24083 19763 24089
rect 28994 24080 29000 24092
rect 29052 24120 29058 24132
rect 29748 24120 29776 24151
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 38286 24188 38292 24200
rect 38247 24160 38292 24188
rect 38286 24148 38292 24160
rect 38344 24148 38350 24200
rect 29052 24092 29776 24120
rect 30009 24123 30067 24129
rect 29052 24080 29058 24092
rect 30009 24089 30021 24123
rect 30055 24089 30067 24123
rect 30009 24083 30067 24089
rect 17552 24024 18460 24052
rect 17552 24012 17558 24024
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19518 24052 19524 24064
rect 19392 24024 19524 24052
rect 19392 24012 19398 24024
rect 19518 24012 19524 24024
rect 19576 24012 19582 24064
rect 24302 24012 24308 24064
rect 24360 24052 24366 24064
rect 30024 24052 30052 24083
rect 30558 24080 30564 24132
rect 30616 24080 30622 24132
rect 35894 24080 35900 24132
rect 35952 24080 35958 24132
rect 31478 24052 31484 24064
rect 24360 24024 30052 24052
rect 31439 24024 31484 24052
rect 24360 24012 24366 24024
rect 31478 24012 31484 24024
rect 31536 24012 31542 24064
rect 33226 24012 33232 24064
rect 33284 24052 33290 24064
rect 36633 24055 36691 24061
rect 36633 24052 36645 24055
rect 33284 24024 36645 24052
rect 33284 24012 33290 24024
rect 36633 24021 36645 24024
rect 36679 24021 36691 24055
rect 36633 24015 36691 24021
rect 38105 24055 38163 24061
rect 38105 24021 38117 24055
rect 38151 24052 38163 24055
rect 38194 24052 38200 24064
rect 38151 24024 38200 24052
rect 38151 24021 38163 24024
rect 38105 24015 38163 24021
rect 38194 24012 38200 24024
rect 38252 24012 38258 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 6270 23808 6276 23860
rect 6328 23848 6334 23860
rect 10505 23851 10563 23857
rect 10505 23848 10517 23851
rect 6328 23820 10517 23848
rect 6328 23808 6334 23820
rect 10505 23817 10517 23820
rect 10551 23817 10563 23851
rect 10505 23811 10563 23817
rect 12250 23808 12256 23860
rect 12308 23848 12314 23860
rect 12897 23851 12955 23857
rect 12897 23848 12909 23851
rect 12308 23820 12909 23848
rect 12308 23808 12314 23820
rect 12897 23817 12909 23820
rect 12943 23817 12955 23851
rect 15746 23848 15752 23860
rect 12897 23811 12955 23817
rect 14660 23820 15752 23848
rect 8294 23780 8300 23792
rect 8255 23752 8300 23780
rect 8294 23740 8300 23752
rect 8352 23740 8358 23792
rect 9953 23783 10011 23789
rect 9953 23749 9965 23783
rect 9999 23780 10011 23783
rect 10962 23780 10968 23792
rect 9999 23752 10968 23780
rect 9999 23749 10011 23752
rect 9953 23743 10011 23749
rect 10962 23740 10968 23752
rect 11020 23740 11026 23792
rect 14660 23780 14688 23820
rect 15746 23808 15752 23820
rect 15804 23848 15810 23860
rect 18138 23848 18144 23860
rect 15804 23820 18144 23848
rect 15804 23808 15810 23820
rect 16206 23780 16212 23792
rect 14568 23752 14688 23780
rect 16054 23752 16212 23780
rect 1946 23672 1952 23724
rect 2004 23712 2010 23724
rect 5537 23715 5595 23721
rect 5537 23712 5549 23715
rect 2004 23684 5549 23712
rect 2004 23672 2010 23684
rect 5537 23681 5549 23684
rect 5583 23681 5595 23715
rect 6730 23712 6736 23724
rect 6691 23684 6736 23712
rect 5537 23675 5595 23681
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 10413 23715 10471 23721
rect 10413 23681 10425 23715
rect 10459 23712 10471 23715
rect 12805 23715 12863 23721
rect 10459 23684 12434 23712
rect 10459 23681 10471 23684
rect 10413 23675 10471 23681
rect 8113 23647 8171 23653
rect 8113 23613 8125 23647
rect 8159 23644 8171 23647
rect 9122 23644 9128 23656
rect 8159 23616 9128 23644
rect 8159 23613 8171 23616
rect 8113 23607 8171 23613
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 3970 23536 3976 23588
rect 4028 23576 4034 23588
rect 6549 23579 6607 23585
rect 6549 23576 6561 23579
rect 4028 23548 6561 23576
rect 4028 23536 4034 23548
rect 6549 23545 6561 23548
rect 6595 23545 6607 23579
rect 12406 23576 12434 23684
rect 12805 23681 12817 23715
rect 12851 23712 12863 23715
rect 14366 23712 14372 23724
rect 12851 23684 14372 23712
rect 12851 23681 12863 23684
rect 12805 23675 12863 23681
rect 14366 23672 14372 23684
rect 14424 23672 14430 23724
rect 14568 23721 14596 23752
rect 16206 23740 16212 23752
rect 16264 23740 16270 23792
rect 16868 23721 16896 23820
rect 18138 23808 18144 23820
rect 18196 23808 18202 23860
rect 18598 23848 18604 23860
rect 18559 23820 18604 23848
rect 18598 23808 18604 23820
rect 18656 23808 18662 23860
rect 18690 23808 18696 23860
rect 18748 23848 18754 23860
rect 24854 23848 24860 23860
rect 18748 23820 21496 23848
rect 18748 23808 18754 23820
rect 20714 23740 20720 23792
rect 20772 23740 20778 23792
rect 21468 23789 21496 23820
rect 22066 23820 24860 23848
rect 21453 23783 21511 23789
rect 21453 23749 21465 23783
rect 21499 23749 21511 23783
rect 21453 23743 21511 23749
rect 14553 23715 14611 23721
rect 14553 23681 14565 23715
rect 14599 23681 14611 23715
rect 14553 23675 14611 23681
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 18230 23672 18236 23724
rect 18288 23672 18294 23724
rect 14829 23647 14887 23653
rect 14829 23613 14841 23647
rect 14875 23644 14887 23647
rect 16758 23644 16764 23656
rect 14875 23616 16764 23644
rect 14875 23613 14887 23616
rect 14829 23607 14887 23613
rect 16758 23604 16764 23616
rect 16816 23604 16822 23656
rect 17494 23644 17500 23656
rect 16868 23616 17500 23644
rect 14550 23576 14556 23588
rect 12406 23548 14556 23576
rect 6549 23539 6607 23545
rect 14550 23536 14556 23548
rect 14608 23536 14614 23588
rect 16301 23579 16359 23585
rect 16301 23545 16313 23579
rect 16347 23576 16359 23579
rect 16868 23576 16896 23616
rect 17494 23604 17500 23616
rect 17552 23604 17558 23656
rect 18138 23604 18144 23656
rect 18196 23644 18202 23656
rect 19429 23647 19487 23653
rect 19429 23644 19441 23647
rect 18196 23616 19441 23644
rect 18196 23604 18202 23616
rect 19429 23613 19441 23616
rect 19475 23613 19487 23647
rect 19429 23607 19487 23613
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23644 19763 23647
rect 20162 23644 20168 23656
rect 19751 23616 20168 23644
rect 19751 23613 19763 23616
rect 19705 23607 19763 23613
rect 20162 23604 20168 23616
rect 20220 23604 20226 23656
rect 20254 23604 20260 23656
rect 20312 23644 20318 23656
rect 22066 23644 22094 23820
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 26970 23808 26976 23860
rect 27028 23848 27034 23860
rect 32674 23848 32680 23860
rect 27028 23820 32680 23848
rect 27028 23808 27034 23820
rect 32674 23808 32680 23820
rect 32732 23808 32738 23860
rect 33502 23808 33508 23860
rect 33560 23848 33566 23860
rect 33962 23848 33968 23860
rect 33560 23820 33968 23848
rect 33560 23808 33566 23820
rect 33962 23808 33968 23820
rect 34020 23848 34026 23860
rect 34057 23851 34115 23857
rect 34057 23848 34069 23851
rect 34020 23820 34069 23848
rect 34020 23808 34026 23820
rect 34057 23817 34069 23820
rect 34103 23817 34115 23851
rect 34057 23811 34115 23817
rect 23934 23780 23940 23792
rect 23895 23752 23940 23780
rect 23934 23740 23940 23752
rect 23992 23740 23998 23792
rect 25682 23780 25688 23792
rect 25162 23752 25688 23780
rect 25682 23740 25688 23752
rect 25740 23740 25746 23792
rect 30282 23780 30288 23792
rect 30130 23752 30288 23780
rect 30282 23740 30288 23752
rect 30340 23740 30346 23792
rect 34330 23780 34336 23792
rect 33810 23752 34336 23780
rect 34330 23740 34336 23752
rect 34388 23740 34394 23792
rect 37458 23780 37464 23792
rect 36018 23752 37464 23780
rect 37458 23740 37464 23752
rect 37516 23740 37522 23792
rect 22278 23672 22284 23724
rect 22336 23712 22342 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 22336 23684 23673 23712
rect 22336 23672 22342 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 34514 23712 34520 23724
rect 34475 23684 34520 23712
rect 23661 23675 23719 23681
rect 34514 23672 34520 23684
rect 34572 23672 34578 23724
rect 20312 23616 22094 23644
rect 20312 23604 20318 23616
rect 25498 23604 25504 23656
rect 25556 23644 25562 23656
rect 25685 23647 25743 23653
rect 25685 23644 25697 23647
rect 25556 23616 25697 23644
rect 25556 23604 25562 23616
rect 25685 23613 25697 23616
rect 25731 23613 25743 23647
rect 25685 23607 25743 23613
rect 28629 23647 28687 23653
rect 28629 23613 28641 23647
rect 28675 23613 28687 23647
rect 28902 23644 28908 23656
rect 28863 23616 28908 23644
rect 28629 23607 28687 23613
rect 16347 23548 16896 23576
rect 18156 23548 18736 23576
rect 16347 23545 16359 23548
rect 16301 23539 16359 23545
rect 5629 23511 5687 23517
rect 5629 23477 5641 23511
rect 5675 23508 5687 23511
rect 9950 23508 9956 23520
rect 5675 23480 9956 23508
rect 5675 23477 5687 23480
rect 5629 23471 5687 23477
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 14366 23468 14372 23520
rect 14424 23508 14430 23520
rect 16316 23508 16344 23539
rect 14424 23480 16344 23508
rect 14424 23468 14430 23480
rect 16666 23468 16672 23520
rect 16724 23508 16730 23520
rect 17116 23511 17174 23517
rect 17116 23508 17128 23511
rect 16724 23480 17128 23508
rect 16724 23468 16730 23480
rect 17116 23477 17128 23480
rect 17162 23508 17174 23511
rect 18156 23508 18184 23548
rect 17162 23480 18184 23508
rect 18708 23508 18736 23548
rect 20990 23508 20996 23520
rect 18708 23480 20996 23508
rect 17162 23477 17174 23480
rect 17116 23471 17174 23477
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 28644 23508 28672 23607
rect 28902 23604 28908 23616
rect 28960 23604 28966 23656
rect 31938 23604 31944 23656
rect 31996 23644 32002 23656
rect 32309 23647 32367 23653
rect 32309 23644 32321 23647
rect 31996 23616 32321 23644
rect 31996 23604 32002 23616
rect 32309 23613 32321 23616
rect 32355 23613 32367 23647
rect 32309 23607 32367 23613
rect 32585 23647 32643 23653
rect 32585 23613 32597 23647
rect 32631 23644 32643 23647
rect 33318 23644 33324 23656
rect 32631 23616 33324 23644
rect 32631 23613 32643 23616
rect 32585 23607 32643 23613
rect 33318 23604 33324 23616
rect 33376 23604 33382 23656
rect 34793 23647 34851 23653
rect 34793 23613 34805 23647
rect 34839 23644 34851 23647
rect 36722 23644 36728 23656
rect 34839 23616 36728 23644
rect 34839 23613 34851 23616
rect 34793 23607 34851 23613
rect 36722 23604 36728 23616
rect 36780 23604 36786 23656
rect 28994 23508 29000 23520
rect 28644 23480 29000 23508
rect 28994 23468 29000 23480
rect 29052 23468 29058 23520
rect 30374 23508 30380 23520
rect 30335 23480 30380 23508
rect 30374 23468 30380 23480
rect 30432 23468 30438 23520
rect 30650 23468 30656 23520
rect 30708 23508 30714 23520
rect 32582 23508 32588 23520
rect 30708 23480 32588 23508
rect 30708 23468 30714 23480
rect 32582 23468 32588 23480
rect 32640 23468 32646 23520
rect 32674 23468 32680 23520
rect 32732 23508 32738 23520
rect 36265 23511 36323 23517
rect 36265 23508 36277 23511
rect 32732 23480 36277 23508
rect 32732 23468 32738 23480
rect 36265 23477 36277 23480
rect 36311 23508 36323 23511
rect 36354 23508 36360 23520
rect 36311 23480 36360 23508
rect 36311 23477 36323 23480
rect 36265 23471 36323 23477
rect 36354 23468 36360 23480
rect 36412 23468 36418 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 9766 23264 9772 23316
rect 9824 23304 9830 23316
rect 13354 23304 13360 23316
rect 9824 23276 13360 23304
rect 9824 23264 9830 23276
rect 13354 23264 13360 23276
rect 13412 23264 13418 23316
rect 15378 23264 15384 23316
rect 15436 23304 15442 23316
rect 16758 23304 16764 23316
rect 15436 23276 16344 23304
rect 16719 23276 16764 23304
rect 15436 23264 15442 23276
rect 8386 23196 8392 23248
rect 8444 23236 8450 23248
rect 16316 23236 16344 23276
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 37826 23304 37832 23316
rect 22020 23276 36952 23304
rect 37787 23276 37832 23304
rect 8444 23208 12480 23236
rect 16316 23208 19932 23236
rect 8444 23196 8450 23208
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9548 23140 9689 23168
rect 9548 23128 9554 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 10318 23168 10324 23180
rect 10279 23140 10324 23168
rect 9677 23131 9735 23137
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 8110 23060 8116 23112
rect 8168 23100 8174 23112
rect 8389 23103 8447 23109
rect 8389 23100 8401 23103
rect 8168 23072 8401 23100
rect 8168 23060 8174 23072
rect 8389 23069 8401 23072
rect 8435 23069 8447 23103
rect 8389 23063 8447 23069
rect 11333 23103 11391 23109
rect 11333 23069 11345 23103
rect 11379 23100 11391 23103
rect 11790 23100 11796 23112
rect 11379 23072 11796 23100
rect 11379 23069 11391 23072
rect 11333 23063 11391 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 12452 23109 12480 23208
rect 15013 23171 15071 23177
rect 15013 23137 15025 23171
rect 15059 23168 15071 23171
rect 15746 23168 15752 23180
rect 15059 23140 15752 23168
rect 15059 23137 15071 23140
rect 15013 23131 15071 23137
rect 15746 23128 15752 23140
rect 15804 23128 15810 23180
rect 19426 23128 19432 23180
rect 19484 23168 19490 23180
rect 19797 23171 19855 23177
rect 19797 23168 19809 23171
rect 19484 23140 19809 23168
rect 19484 23128 19490 23140
rect 19797 23137 19809 23140
rect 19843 23137 19855 23171
rect 19904 23168 19932 23208
rect 21821 23171 21879 23177
rect 21821 23168 21833 23171
rect 19904 23140 21833 23168
rect 19797 23131 19855 23137
rect 21821 23137 21833 23140
rect 21867 23137 21879 23171
rect 21821 23131 21879 23137
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 13081 23103 13139 23109
rect 13081 23069 13093 23103
rect 13127 23100 13139 23103
rect 13127 23072 15056 23100
rect 13127 23069 13139 23072
rect 13081 23063 13139 23069
rect 9766 23032 9772 23044
rect 9727 23004 9772 23032
rect 9766 22992 9772 23004
rect 9824 22992 9830 23044
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 13173 23035 13231 23041
rect 13173 23032 13185 23035
rect 11940 23004 13185 23032
rect 11940 22992 11946 23004
rect 13173 23001 13185 23004
rect 13219 23001 13231 23035
rect 13173 22995 13231 23001
rect 8481 22967 8539 22973
rect 8481 22933 8493 22967
rect 8527 22964 8539 22967
rect 9398 22964 9404 22976
rect 8527 22936 9404 22964
rect 8527 22933 8539 22936
rect 8481 22927 8539 22933
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 11238 22924 11244 22976
rect 11296 22964 11302 22976
rect 11425 22967 11483 22973
rect 11425 22964 11437 22967
rect 11296 22936 11437 22964
rect 11296 22924 11302 22936
rect 11425 22933 11437 22936
rect 11471 22933 11483 22967
rect 11425 22927 11483 22933
rect 11790 22924 11796 22976
rect 11848 22964 11854 22976
rect 12158 22964 12164 22976
rect 11848 22936 12164 22964
rect 11848 22924 11854 22936
rect 12158 22924 12164 22936
rect 12216 22924 12222 22976
rect 12526 22924 12532 22976
rect 12584 22964 12590 22976
rect 15028 22964 15056 23072
rect 15286 23032 15292 23044
rect 15247 23004 15292 23032
rect 15286 22992 15292 23004
rect 15344 22992 15350 23044
rect 17402 23032 17408 23044
rect 16514 23004 17408 23032
rect 17402 22992 17408 23004
rect 17460 22992 17466 23044
rect 17678 22992 17684 23044
rect 17736 23032 17742 23044
rect 18690 23032 18696 23044
rect 17736 23004 18696 23032
rect 17736 22992 17742 23004
rect 18690 22992 18696 23004
rect 18748 22992 18754 23044
rect 20070 23032 20076 23044
rect 20031 23004 20076 23032
rect 20070 22992 20076 23004
rect 20128 22992 20134 23044
rect 21358 23032 21364 23044
rect 21298 23004 21364 23032
rect 21358 22992 21364 23004
rect 21416 22992 21422 23044
rect 21818 22992 21824 23044
rect 21876 23032 21882 23044
rect 22020 23032 22048 23276
rect 33318 23196 33324 23248
rect 33376 23236 33382 23248
rect 33686 23236 33692 23248
rect 33376 23208 33692 23236
rect 33376 23196 33382 23208
rect 33686 23196 33692 23208
rect 33744 23196 33750 23248
rect 22278 23168 22284 23180
rect 22239 23140 22284 23168
rect 22278 23128 22284 23140
rect 22336 23128 22342 23180
rect 23750 23128 23756 23180
rect 23808 23168 23814 23180
rect 24029 23171 24087 23177
rect 24029 23168 24041 23171
rect 23808 23140 24041 23168
rect 23808 23128 23814 23140
rect 24029 23137 24041 23140
rect 24075 23168 24087 23171
rect 26053 23171 26111 23177
rect 26053 23168 26065 23171
rect 24075 23140 26065 23168
rect 24075 23137 24087 23140
rect 24029 23131 24087 23137
rect 26053 23137 26065 23140
rect 26099 23137 26111 23171
rect 26053 23131 26111 23137
rect 28994 23128 29000 23180
rect 29052 23168 29058 23180
rect 29733 23171 29791 23177
rect 29733 23168 29745 23171
rect 29052 23140 29745 23168
rect 29052 23128 29058 23140
rect 29733 23137 29745 23140
rect 29779 23137 29791 23171
rect 29733 23131 29791 23137
rect 30466 23128 30472 23180
rect 30524 23168 30530 23180
rect 30650 23168 30656 23180
rect 30524 23140 30656 23168
rect 30524 23128 30530 23140
rect 30650 23128 30656 23140
rect 30708 23168 30714 23180
rect 31481 23171 31539 23177
rect 31481 23168 31493 23171
rect 30708 23140 31493 23168
rect 30708 23128 30714 23140
rect 31481 23137 31493 23140
rect 31527 23137 31539 23171
rect 31481 23131 31539 23137
rect 32217 23171 32275 23177
rect 32217 23137 32229 23171
rect 32263 23168 32275 23171
rect 33226 23168 33232 23180
rect 32263 23140 33232 23168
rect 32263 23137 32275 23140
rect 32217 23131 32275 23137
rect 33226 23128 33232 23140
rect 33284 23128 33290 23180
rect 34606 23128 34612 23180
rect 34664 23168 34670 23180
rect 34885 23171 34943 23177
rect 34885 23168 34897 23171
rect 34664 23140 34897 23168
rect 34664 23128 34670 23140
rect 34885 23137 34897 23140
rect 34931 23137 34943 23171
rect 34885 23131 34943 23137
rect 35161 23171 35219 23177
rect 35161 23137 35173 23171
rect 35207 23168 35219 23171
rect 35618 23168 35624 23180
rect 35207 23140 35624 23168
rect 35207 23137 35219 23140
rect 35161 23131 35219 23137
rect 35618 23128 35624 23140
rect 35676 23168 35682 23180
rect 35802 23168 35808 23180
rect 35676 23140 35808 23168
rect 35676 23128 35682 23140
rect 35802 23128 35808 23140
rect 35860 23128 35866 23180
rect 36924 23177 36952 23276
rect 37826 23264 37832 23276
rect 37884 23264 37890 23316
rect 36909 23171 36967 23177
rect 36909 23137 36921 23171
rect 36955 23137 36967 23171
rect 36909 23131 36967 23137
rect 25774 23100 25780 23112
rect 25735 23072 25780 23100
rect 25774 23060 25780 23072
rect 25832 23060 25838 23112
rect 31570 23100 31576 23112
rect 31142 23072 31576 23100
rect 31570 23060 31576 23072
rect 31628 23060 31634 23112
rect 31938 23100 31944 23112
rect 31899 23072 31944 23100
rect 31938 23060 31944 23072
rect 31996 23060 32002 23112
rect 38013 23103 38071 23109
rect 38013 23069 38025 23103
rect 38059 23100 38071 23103
rect 38194 23100 38200 23112
rect 38059 23072 38200 23100
rect 38059 23069 38071 23072
rect 38013 23063 38071 23069
rect 38194 23060 38200 23072
rect 38252 23100 38258 23112
rect 39022 23100 39028 23112
rect 38252 23072 39028 23100
rect 38252 23060 38258 23072
rect 39022 23060 39028 23072
rect 39080 23060 39086 23112
rect 22557 23035 22615 23041
rect 22557 23032 22569 23035
rect 21876 23004 22569 23032
rect 21876 22992 21882 23004
rect 22557 23001 22569 23004
rect 22603 23001 22615 23035
rect 25958 23032 25964 23044
rect 23782 23004 25964 23032
rect 22557 22995 22615 23001
rect 25958 22992 25964 23004
rect 26016 22992 26022 23044
rect 27062 22992 27068 23044
rect 27120 22992 27126 23044
rect 27801 23035 27859 23041
rect 27801 23001 27813 23035
rect 27847 23001 27859 23035
rect 27801 22995 27859 23001
rect 21450 22964 21456 22976
rect 12584 22936 12629 22964
rect 15028 22936 21456 22964
rect 12584 22924 12590 22936
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 27816 22964 27844 22995
rect 29362 22992 29368 23044
rect 29420 23032 29426 23044
rect 29914 23032 29920 23044
rect 29420 23004 29920 23032
rect 29420 22992 29426 23004
rect 29914 22992 29920 23004
rect 29972 23032 29978 23044
rect 30009 23035 30067 23041
rect 30009 23032 30021 23035
rect 29972 23004 30021 23032
rect 29972 22992 29978 23004
rect 30009 23001 30021 23004
rect 30055 23001 30067 23035
rect 33870 23032 33876 23044
rect 30009 22995 30067 23001
rect 31404 23004 31754 23032
rect 33442 23004 33876 23032
rect 31404 22964 31432 23004
rect 27816 22936 31432 22964
rect 31726 22964 31754 23004
rect 33870 22992 33876 23004
rect 33928 22992 33934 23044
rect 37826 23032 37832 23044
rect 36386 23004 37832 23032
rect 37826 22992 37832 23004
rect 37884 22992 37890 23044
rect 32030 22964 32036 22976
rect 31726 22936 32036 22964
rect 32030 22924 32036 22936
rect 32088 22964 32094 22976
rect 32490 22964 32496 22976
rect 32088 22936 32496 22964
rect 32088 22924 32094 22936
rect 32490 22924 32496 22936
rect 32548 22924 32554 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 7282 22760 7288 22772
rect 1627 22732 7288 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 8662 22760 8668 22772
rect 8444 22732 8668 22760
rect 8444 22720 8450 22732
rect 8662 22720 8668 22732
rect 8720 22720 8726 22772
rect 12989 22763 13047 22769
rect 12989 22729 13001 22763
rect 13035 22760 13047 22763
rect 15194 22760 15200 22772
rect 13035 22732 15200 22760
rect 13035 22729 13047 22732
rect 12989 22723 13047 22729
rect 15194 22720 15200 22732
rect 15252 22720 15258 22772
rect 20990 22760 20996 22772
rect 17604 22732 20996 22760
rect 9398 22692 9404 22704
rect 9359 22664 9404 22692
rect 9398 22652 9404 22664
rect 9456 22652 9462 22704
rect 11882 22692 11888 22704
rect 11843 22664 11888 22692
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 17604 22692 17632 22732
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 21358 22720 21364 22772
rect 21416 22760 21422 22772
rect 22097 22763 22155 22769
rect 22097 22760 22109 22763
rect 21416 22732 22109 22760
rect 21416 22720 21422 22732
rect 22097 22729 22109 22732
rect 22143 22729 22155 22763
rect 22097 22723 22155 22729
rect 22370 22720 22376 22772
rect 22428 22760 22434 22772
rect 26510 22760 26516 22772
rect 22428 22732 26516 22760
rect 22428 22720 22434 22732
rect 26510 22720 26516 22732
rect 26568 22720 26574 22772
rect 28994 22760 29000 22772
rect 27172 22732 29000 22760
rect 17862 22692 17868 22704
rect 12584 22664 17632 22692
rect 17696 22664 17868 22692
rect 12584 22652 12590 22664
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 11054 22624 11060 22636
rect 10827 22596 11060 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 12802 22584 12808 22636
rect 12860 22624 12866 22636
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12860 22596 12909 22624
rect 12860 22584 12866 22596
rect 12897 22593 12909 22596
rect 12943 22624 12955 22627
rect 12986 22624 12992 22636
rect 12943 22596 12992 22624
rect 12943 22593 12955 22596
rect 12897 22587 12955 22593
rect 12986 22584 12992 22596
rect 13044 22584 13050 22636
rect 17696 22633 17724 22664
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 19426 22692 19432 22704
rect 19182 22664 19432 22692
rect 19426 22652 19432 22664
rect 19484 22652 19490 22704
rect 19705 22695 19763 22701
rect 19705 22661 19717 22695
rect 19751 22692 19763 22695
rect 20254 22692 20260 22704
rect 19751 22664 20260 22692
rect 19751 22661 19763 22664
rect 19705 22655 19763 22661
rect 20254 22652 20260 22664
rect 20312 22652 20318 22704
rect 24486 22692 24492 22704
rect 24150 22664 24492 22692
rect 24486 22652 24492 22664
rect 24544 22652 24550 22704
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 22002 22624 22008 22636
rect 21963 22596 22008 22624
rect 17681 22587 17739 22593
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 22278 22584 22284 22636
rect 22336 22624 22342 22636
rect 22649 22627 22707 22633
rect 22649 22624 22661 22627
rect 22336 22596 22661 22624
rect 22336 22584 22342 22596
rect 22649 22593 22661 22596
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 24302 22584 24308 22636
rect 24360 22624 24366 22636
rect 24673 22627 24731 22633
rect 24673 22624 24685 22627
rect 24360 22596 24685 22624
rect 24360 22584 24366 22596
rect 24673 22593 24685 22596
rect 24719 22593 24731 22627
rect 24673 22587 24731 22593
rect 25774 22584 25780 22636
rect 25832 22624 25838 22636
rect 27172 22633 27200 22732
rect 28994 22720 29000 22732
rect 29052 22720 29058 22772
rect 36078 22760 36084 22772
rect 35636 22732 36084 22760
rect 27430 22692 27436 22704
rect 27391 22664 27436 22692
rect 27430 22652 27436 22664
rect 27488 22652 27494 22704
rect 28442 22652 28448 22704
rect 28500 22652 28506 22704
rect 35636 22692 35664 22732
rect 36078 22720 36084 22732
rect 36136 22720 36142 22772
rect 36538 22720 36544 22772
rect 36596 22760 36602 22772
rect 36722 22760 36728 22772
rect 36596 22732 36728 22760
rect 36596 22720 36602 22732
rect 36722 22720 36728 22732
rect 36780 22720 36786 22772
rect 37550 22692 37556 22704
rect 34270 22664 35664 22692
rect 36478 22664 37556 22692
rect 37550 22652 37556 22664
rect 37608 22652 37614 22704
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 25832 22596 27169 22624
rect 25832 22584 25838 22596
rect 27157 22593 27169 22596
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 31938 22584 31944 22636
rect 31996 22624 32002 22636
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 31996 22596 32781 22624
rect 31996 22584 32002 22596
rect 32769 22593 32781 22596
rect 32815 22593 32827 22627
rect 32769 22587 32827 22593
rect 34606 22584 34612 22636
rect 34664 22624 34670 22636
rect 34977 22627 35035 22633
rect 34977 22624 34989 22627
rect 34664 22596 34989 22624
rect 34664 22584 34670 22596
rect 34977 22593 34989 22596
rect 35023 22593 35035 22627
rect 34977 22587 35035 22593
rect 37642 22584 37648 22636
rect 37700 22624 37706 22636
rect 38013 22627 38071 22633
rect 38013 22624 38025 22627
rect 37700 22596 38025 22624
rect 37700 22584 37706 22596
rect 38013 22593 38025 22596
rect 38059 22593 38071 22627
rect 38013 22587 38071 22593
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22556 4583 22559
rect 4614 22556 4620 22568
rect 4571 22528 4620 22556
rect 4571 22525 4583 22528
rect 4525 22519 4583 22525
rect 4614 22516 4620 22528
rect 4672 22516 4678 22568
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 9309 22559 9367 22565
rect 9309 22556 9321 22559
rect 9180 22528 9321 22556
rect 9180 22516 9186 22528
rect 9309 22525 9321 22528
rect 9355 22525 9367 22559
rect 9309 22519 9367 22525
rect 10321 22559 10379 22565
rect 10321 22525 10333 22559
rect 10367 22556 10379 22559
rect 11146 22556 11152 22568
rect 10367 22528 11152 22556
rect 10367 22525 10379 22528
rect 10321 22519 10379 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 11790 22556 11796 22568
rect 11751 22528 11796 22556
rect 11790 22516 11796 22528
rect 11848 22516 11854 22568
rect 12069 22559 12127 22565
rect 12069 22525 12081 22559
rect 12115 22525 12127 22559
rect 12069 22519 12127 22525
rect 17957 22559 18015 22565
rect 17957 22525 17969 22559
rect 18003 22556 18015 22559
rect 18046 22556 18052 22568
rect 18003 22528 18052 22556
rect 18003 22525 18015 22528
rect 17957 22519 18015 22525
rect 11698 22448 11704 22500
rect 11756 22488 11762 22500
rect 12084 22488 12112 22519
rect 18046 22516 18052 22528
rect 18104 22556 18110 22568
rect 18322 22556 18328 22568
rect 18104 22528 18328 22556
rect 18104 22516 18110 22528
rect 18322 22516 18328 22528
rect 18380 22516 18386 22568
rect 22925 22559 22983 22565
rect 19812 22528 22692 22556
rect 11756 22460 12112 22488
rect 11756 22448 11762 22460
rect 12342 22448 12348 22500
rect 12400 22488 12406 22500
rect 12802 22488 12808 22500
rect 12400 22460 12808 22488
rect 12400 22448 12406 22460
rect 12802 22448 12808 22460
rect 12860 22448 12866 22500
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 10873 22423 10931 22429
rect 10873 22420 10885 22423
rect 9732 22392 10885 22420
rect 9732 22380 9738 22392
rect 10873 22389 10885 22392
rect 10919 22389 10931 22423
rect 10873 22383 10931 22389
rect 13630 22380 13636 22432
rect 13688 22420 13694 22432
rect 19812 22420 19840 22528
rect 20070 22448 20076 22500
rect 20128 22488 20134 22500
rect 22370 22488 22376 22500
rect 20128 22460 22376 22488
rect 20128 22448 20134 22460
rect 22370 22448 22376 22460
rect 22428 22448 22434 22500
rect 13688 22392 19840 22420
rect 22664 22420 22692 22528
rect 22925 22525 22937 22559
rect 22971 22556 22983 22559
rect 28902 22556 28908 22568
rect 22971 22528 24624 22556
rect 28863 22528 28908 22556
rect 22971 22525 22983 22528
rect 22925 22519 22983 22525
rect 24596 22488 24624 22528
rect 28902 22516 28908 22528
rect 28960 22516 28966 22568
rect 31478 22516 31484 22568
rect 31536 22556 31542 22568
rect 31662 22556 31668 22568
rect 31536 22528 31668 22556
rect 31536 22516 31542 22528
rect 31662 22516 31668 22528
rect 31720 22556 31726 22568
rect 33045 22559 33103 22565
rect 33045 22556 33057 22559
rect 31720 22528 33057 22556
rect 31720 22516 31726 22528
rect 33045 22525 33057 22528
rect 33091 22525 33103 22559
rect 33045 22519 33103 22525
rect 33134 22516 33140 22568
rect 33192 22556 33198 22568
rect 35253 22559 35311 22565
rect 35253 22556 35265 22559
rect 33192 22528 35265 22556
rect 33192 22516 33198 22528
rect 35253 22525 35265 22528
rect 35299 22525 35311 22559
rect 35253 22519 35311 22525
rect 25498 22488 25504 22500
rect 24596 22460 25504 22488
rect 25498 22448 25504 22460
rect 25556 22448 25562 22500
rect 38194 22488 38200 22500
rect 38155 22460 38200 22488
rect 38194 22448 38200 22460
rect 38252 22448 38258 22500
rect 23382 22420 23388 22432
rect 22664 22392 23388 22420
rect 13688 22380 13694 22392
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 33134 22380 33140 22432
rect 33192 22420 33198 22432
rect 34517 22423 34575 22429
rect 34517 22420 34529 22423
rect 33192 22392 34529 22420
rect 33192 22380 33198 22392
rect 34517 22389 34529 22392
rect 34563 22389 34575 22423
rect 34517 22383 34575 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 18414 22216 18420 22228
rect 15620 22188 18420 22216
rect 15620 22176 15626 22188
rect 18414 22176 18420 22188
rect 18472 22176 18478 22228
rect 18690 22216 18696 22228
rect 18651 22188 18696 22216
rect 18690 22176 18696 22188
rect 18748 22176 18754 22228
rect 20070 22176 20076 22228
rect 20128 22216 20134 22228
rect 20254 22216 20260 22228
rect 20128 22188 20260 22216
rect 20128 22176 20134 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 25590 22176 25596 22228
rect 25648 22216 25654 22228
rect 25758 22219 25816 22225
rect 25758 22216 25770 22219
rect 25648 22188 25770 22216
rect 25648 22176 25654 22188
rect 25758 22185 25770 22188
rect 25804 22185 25816 22219
rect 25758 22179 25816 22185
rect 34698 22176 34704 22228
rect 34756 22216 34762 22228
rect 34882 22216 34888 22228
rect 34756 22188 34888 22216
rect 34756 22176 34762 22188
rect 34882 22176 34888 22188
rect 34940 22176 34946 22228
rect 36446 22176 36452 22228
rect 36504 22216 36510 22228
rect 36817 22219 36875 22225
rect 36817 22216 36829 22219
rect 36504 22188 36829 22216
rect 36504 22176 36510 22188
rect 36817 22185 36829 22188
rect 36863 22185 36875 22219
rect 36817 22179 36875 22185
rect 4614 22148 4620 22160
rect 4448 22120 4620 22148
rect 4448 22089 4476 22120
rect 4614 22108 4620 22120
rect 4672 22108 4678 22160
rect 12066 22108 12072 22160
rect 12124 22148 12130 22160
rect 12124 22120 22232 22148
rect 12124 22108 12130 22120
rect 4433 22083 4491 22089
rect 4433 22049 4445 22083
rect 4479 22049 4491 22083
rect 9214 22080 9220 22092
rect 4433 22043 4491 22049
rect 9048 22052 9220 22080
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 22012 4675 22015
rect 4798 22012 4804 22024
rect 4663 21984 4804 22012
rect 4663 21981 4675 21984
rect 4617 21975 4675 21981
rect 4798 21972 4804 21984
rect 4856 21972 4862 22024
rect 8386 22012 8392 22024
rect 8299 21984 8392 22012
rect 8386 21972 8392 21984
rect 8444 22012 8450 22024
rect 9048 22012 9076 22052
rect 9214 22040 9220 22052
rect 9272 22040 9278 22092
rect 9861 22083 9919 22089
rect 9861 22049 9873 22083
rect 9907 22080 9919 22083
rect 10594 22080 10600 22092
rect 9907 22052 10600 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 10594 22040 10600 22052
rect 10652 22040 10658 22092
rect 10870 22040 10876 22092
rect 10928 22080 10934 22092
rect 12526 22080 12532 22092
rect 10928 22052 12532 22080
rect 10928 22040 10934 22052
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 12802 22080 12808 22092
rect 12763 22052 12808 22080
rect 12802 22040 12808 22052
rect 12860 22040 12866 22092
rect 16209 22083 16267 22089
rect 16209 22080 16221 22083
rect 13188 22052 16221 22080
rect 8444 21984 9076 22012
rect 13188 22006 13216 22052
rect 16209 22049 16221 22052
rect 16255 22049 16267 22083
rect 20714 22080 20720 22092
rect 20675 22052 20720 22080
rect 16209 22043 16267 22049
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 22204 22089 22232 22120
rect 24486 22108 24492 22160
rect 24544 22148 24550 22160
rect 24762 22148 24768 22160
rect 24544 22120 24768 22148
rect 24544 22108 24550 22120
rect 24762 22108 24768 22120
rect 24820 22108 24826 22160
rect 22189 22083 22247 22089
rect 22189 22049 22201 22083
rect 22235 22080 22247 22083
rect 23014 22080 23020 22092
rect 22235 22052 22876 22080
rect 22975 22052 23020 22080
rect 22235 22049 22247 22052
rect 22189 22043 22247 22049
rect 8444 21972 8450 21984
rect 13004 21978 13216 22006
rect 16117 22015 16175 22021
rect 16117 21981 16129 22015
rect 16163 22012 16175 22015
rect 18625 22015 18683 22021
rect 16163 21984 17724 22012
rect 16163 21981 16175 21984
rect 8018 21904 8024 21956
rect 8076 21944 8082 21956
rect 8076 21916 8616 21944
rect 8076 21904 8082 21916
rect 5077 21879 5135 21885
rect 5077 21845 5089 21879
rect 5123 21876 5135 21879
rect 5626 21876 5632 21888
rect 5123 21848 5632 21876
rect 5123 21845 5135 21848
rect 5077 21839 5135 21845
rect 5626 21836 5632 21848
rect 5684 21836 5690 21888
rect 7558 21836 7564 21888
rect 7616 21876 7622 21888
rect 8481 21879 8539 21885
rect 8481 21876 8493 21879
rect 7616 21848 8493 21876
rect 7616 21836 7622 21848
rect 8481 21845 8493 21848
rect 8527 21845 8539 21879
rect 8588 21876 8616 21916
rect 9030 21904 9036 21956
rect 9088 21944 9094 21956
rect 9217 21947 9275 21953
rect 9217 21944 9229 21947
rect 9088 21916 9229 21944
rect 9088 21904 9094 21916
rect 9217 21913 9229 21916
rect 9263 21913 9275 21947
rect 9217 21907 9275 21913
rect 9309 21947 9367 21953
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 9674 21944 9680 21956
rect 9355 21916 9680 21944
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 10410 21904 10416 21956
rect 10468 21944 10474 21956
rect 10962 21944 10968 21956
rect 10468 21916 10968 21944
rect 10468 21904 10474 21916
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 12342 21944 12348 21956
rect 12303 21916 12348 21944
rect 12342 21904 12348 21916
rect 12400 21904 12406 21956
rect 12437 21947 12495 21953
rect 12437 21913 12449 21947
rect 12483 21944 12495 21947
rect 13004 21944 13032 21978
rect 16117 21975 16175 21981
rect 12483 21916 13032 21944
rect 14645 21947 14703 21953
rect 12483 21913 12495 21916
rect 12437 21907 12495 21913
rect 14645 21913 14657 21947
rect 14691 21913 14703 21947
rect 14645 21907 14703 21913
rect 12250 21876 12256 21888
rect 8588 21848 12256 21876
rect 8481 21839 8539 21845
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 12526 21836 12532 21888
rect 12584 21876 12590 21888
rect 14660 21876 14688 21907
rect 14734 21904 14740 21956
rect 14792 21944 14798 21956
rect 15657 21947 15715 21953
rect 14792 21916 14837 21944
rect 14792 21904 14798 21916
rect 15657 21913 15669 21947
rect 15703 21944 15715 21947
rect 16758 21944 16764 21956
rect 15703 21916 16764 21944
rect 15703 21913 15715 21916
rect 15657 21907 15715 21913
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 16942 21904 16948 21956
rect 17000 21944 17006 21956
rect 17126 21944 17132 21956
rect 17000 21916 17132 21944
rect 17000 21904 17006 21916
rect 17126 21904 17132 21916
rect 17184 21904 17190 21956
rect 12584 21848 14688 21876
rect 17696 21876 17724 21984
rect 18625 21981 18637 22015
rect 18671 22012 18683 22015
rect 19242 22012 19248 22024
rect 18671 21984 19248 22012
rect 18671 21981 18683 21984
rect 18625 21975 18683 21981
rect 19242 21972 19248 21984
rect 19300 22012 19306 22024
rect 20438 22012 20444 22024
rect 19300 21984 20444 22012
rect 19300 21972 19306 21984
rect 20438 21972 20444 21984
rect 20496 22012 20502 22024
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 20496 21984 20637 22012
rect 20496 21972 20502 21984
rect 20625 21981 20637 21984
rect 20671 21981 20683 22015
rect 22741 22015 22799 22021
rect 22741 22012 22753 22015
rect 20625 21975 20683 21981
rect 22204 21984 22753 22012
rect 22204 21956 22232 21984
rect 22741 21981 22753 21984
rect 22787 21981 22799 22015
rect 22848 22012 22876 22052
rect 23014 22040 23020 22052
rect 23072 22040 23078 22092
rect 25501 22083 25559 22089
rect 25501 22049 25513 22083
rect 25547 22080 25559 22083
rect 25774 22080 25780 22092
rect 25547 22052 25780 22080
rect 25547 22049 25559 22052
rect 25501 22043 25559 22049
rect 25774 22040 25780 22052
rect 25832 22040 25838 22092
rect 31021 22083 31079 22089
rect 31021 22049 31033 22083
rect 31067 22080 31079 22083
rect 31938 22080 31944 22092
rect 31067 22052 31944 22080
rect 31067 22049 31079 22052
rect 31021 22043 31079 22049
rect 31938 22040 31944 22052
rect 31996 22040 32002 22092
rect 32306 22040 32312 22092
rect 32364 22080 32370 22092
rect 32858 22080 32864 22092
rect 32364 22052 32864 22080
rect 32364 22040 32370 22052
rect 32858 22040 32864 22052
rect 32916 22040 32922 22092
rect 37458 22080 37464 22092
rect 37419 22052 37464 22080
rect 37458 22040 37464 22052
rect 37516 22040 37522 22092
rect 23290 22012 23296 22024
rect 22848 21984 23296 22012
rect 22741 21975 22799 21981
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 36446 21972 36452 22024
rect 36504 22012 36510 22024
rect 36725 22015 36783 22021
rect 36725 22012 36737 22015
rect 36504 21984 36737 22012
rect 36504 21972 36510 21984
rect 36725 21981 36737 21984
rect 36771 22012 36783 22015
rect 37182 22012 37188 22024
rect 36771 21984 37188 22012
rect 36771 21981 36783 21984
rect 36725 21975 36783 21981
rect 37182 21972 37188 21984
rect 37240 22012 37246 22024
rect 37369 22015 37427 22021
rect 37369 22012 37381 22015
rect 37240 21984 37381 22012
rect 37240 21972 37246 21984
rect 37369 21981 37381 21984
rect 37415 21981 37427 22015
rect 38010 22012 38016 22024
rect 37971 21984 38016 22012
rect 37369 21975 37427 21981
rect 38010 21972 38016 21984
rect 38068 21972 38074 22024
rect 21361 21947 21419 21953
rect 21361 21913 21373 21947
rect 21407 21944 21419 21947
rect 22186 21944 22192 21956
rect 21407 21916 22192 21944
rect 21407 21913 21419 21916
rect 21361 21907 21419 21913
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 27430 21944 27436 21956
rect 27002 21916 27436 21944
rect 27430 21904 27436 21916
rect 27488 21904 27494 21956
rect 31202 21904 31208 21956
rect 31260 21944 31266 21956
rect 31297 21947 31355 21953
rect 31297 21944 31309 21947
rect 31260 21916 31309 21944
rect 31260 21904 31266 21916
rect 31297 21913 31309 21916
rect 31343 21913 31355 21947
rect 34790 21944 34796 21956
rect 32522 21916 34796 21944
rect 31297 21907 31355 21913
rect 34790 21904 34796 21916
rect 34848 21904 34854 21956
rect 34974 21944 34980 21956
rect 34935 21916 34980 21944
rect 34974 21904 34980 21916
rect 35032 21904 35038 21956
rect 35066 21904 35072 21956
rect 35124 21944 35130 21956
rect 35124 21916 35169 21944
rect 35124 21904 35130 21916
rect 35434 21904 35440 21956
rect 35492 21944 35498 21956
rect 35989 21947 36047 21953
rect 35989 21944 36001 21947
rect 35492 21916 36001 21944
rect 35492 21904 35498 21916
rect 35989 21913 36001 21916
rect 36035 21913 36047 21947
rect 35989 21907 36047 21913
rect 21266 21876 21272 21888
rect 17696 21848 21272 21876
rect 12584 21836 12590 21848
rect 21266 21836 21272 21848
rect 21324 21836 21330 21888
rect 26786 21836 26792 21888
rect 26844 21876 26850 21888
rect 27154 21876 27160 21888
rect 26844 21848 27160 21876
rect 26844 21836 26850 21848
rect 27154 21836 27160 21848
rect 27212 21876 27218 21888
rect 27249 21879 27307 21885
rect 27249 21876 27261 21879
rect 27212 21848 27261 21876
rect 27212 21836 27218 21848
rect 27249 21845 27261 21848
rect 27295 21845 27307 21879
rect 27249 21839 27307 21845
rect 32769 21879 32827 21885
rect 32769 21845 32781 21879
rect 32815 21876 32827 21879
rect 32858 21876 32864 21888
rect 32815 21848 32864 21876
rect 32815 21845 32827 21848
rect 32769 21839 32827 21845
rect 32858 21836 32864 21848
rect 32916 21836 32922 21888
rect 36538 21836 36544 21888
rect 36596 21876 36602 21888
rect 36906 21876 36912 21888
rect 36596 21848 36912 21876
rect 36596 21836 36602 21848
rect 36906 21836 36912 21848
rect 36964 21836 36970 21888
rect 38194 21876 38200 21888
rect 38155 21848 38200 21876
rect 38194 21836 38200 21848
rect 38252 21836 38258 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 4798 21672 4804 21684
rect 4759 21644 4804 21672
rect 4798 21632 4804 21644
rect 4856 21632 4862 21684
rect 5445 21675 5503 21681
rect 5445 21641 5457 21675
rect 5491 21641 5503 21675
rect 12250 21672 12256 21684
rect 5445 21635 5503 21641
rect 5552 21644 12256 21672
rect 1670 21536 1676 21548
rect 1631 21508 1676 21536
rect 1670 21496 1676 21508
rect 1728 21496 1734 21548
rect 1946 21496 1952 21548
rect 2004 21536 2010 21548
rect 2501 21539 2559 21545
rect 2501 21536 2513 21539
rect 2004 21508 2513 21536
rect 2004 21496 2010 21508
rect 2501 21505 2513 21508
rect 2547 21505 2559 21539
rect 2501 21499 2559 21505
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21536 5043 21539
rect 5460 21536 5488 21635
rect 5031 21508 5488 21536
rect 5031 21505 5043 21508
rect 4985 21499 5043 21505
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21400 1915 21403
rect 5552 21400 5580 21644
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 23934 21672 23940 21684
rect 16816 21644 23940 21672
rect 16816 21632 16822 21644
rect 23934 21632 23940 21644
rect 23992 21632 23998 21684
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25041 21675 25099 21681
rect 25041 21672 25053 21675
rect 24820 21644 25053 21672
rect 24820 21632 24826 21644
rect 25041 21641 25053 21644
rect 25087 21641 25099 21675
rect 25041 21635 25099 21641
rect 30469 21675 30527 21681
rect 30469 21641 30481 21675
rect 30515 21672 30527 21675
rect 30558 21672 30564 21684
rect 30515 21644 30564 21672
rect 30515 21641 30527 21644
rect 30469 21635 30527 21641
rect 30558 21632 30564 21644
rect 30616 21632 30622 21684
rect 31665 21675 31723 21681
rect 31665 21641 31677 21675
rect 31711 21672 31723 21675
rect 35066 21672 35072 21684
rect 31711 21644 35072 21672
rect 31711 21641 31723 21644
rect 31665 21635 31723 21641
rect 35066 21632 35072 21644
rect 35124 21632 35130 21684
rect 35710 21672 35716 21684
rect 35671 21644 35716 21672
rect 35710 21632 35716 21644
rect 35768 21632 35774 21684
rect 36633 21675 36691 21681
rect 36633 21672 36645 21675
rect 35820 21644 36645 21672
rect 8570 21604 8576 21616
rect 5644 21576 8576 21604
rect 5644 21545 5672 21576
rect 8570 21564 8576 21576
rect 8628 21564 8634 21616
rect 9217 21607 9275 21613
rect 9217 21573 9229 21607
rect 9263 21604 9275 21607
rect 12158 21604 12164 21616
rect 9263 21576 12164 21604
rect 9263 21573 9275 21576
rect 9217 21567 9275 21573
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 13173 21607 13231 21613
rect 13173 21573 13185 21607
rect 13219 21604 13231 21607
rect 13630 21604 13636 21616
rect 13219 21576 13636 21604
rect 13219 21573 13231 21576
rect 13173 21567 13231 21573
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 16206 21564 16212 21616
rect 16264 21604 16270 21616
rect 17773 21607 17831 21613
rect 17773 21604 17785 21607
rect 16264 21576 17785 21604
rect 16264 21564 16270 21576
rect 17773 21573 17785 21576
rect 17819 21573 17831 21607
rect 21269 21607 21327 21613
rect 21269 21604 21281 21607
rect 17773 21567 17831 21573
rect 19168 21576 21281 21604
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 7650 21496 7656 21548
rect 7708 21536 7714 21548
rect 7708 21508 7753 21536
rect 7708 21496 7714 21508
rect 10502 21496 10508 21548
rect 10560 21536 10566 21548
rect 10597 21539 10655 21545
rect 10597 21536 10609 21539
rect 10560 21508 10609 21536
rect 10560 21496 10566 21508
rect 10597 21505 10609 21508
rect 10643 21536 10655 21539
rect 11790 21536 11796 21548
rect 10643 21508 11796 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 11790 21496 11796 21508
rect 11848 21496 11854 21548
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21536 12403 21539
rect 12526 21536 12532 21548
rect 12391 21508 12532 21536
rect 12391 21505 12403 21508
rect 12345 21499 12403 21505
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 13081 21539 13139 21545
rect 13081 21534 13093 21539
rect 13004 21506 13093 21534
rect 8389 21471 8447 21477
rect 8389 21437 8401 21471
rect 8435 21468 8447 21471
rect 9125 21471 9183 21477
rect 9125 21468 9137 21471
rect 8435 21440 9137 21468
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 9125 21437 9137 21440
rect 9171 21437 9183 21471
rect 9125 21431 9183 21437
rect 9214 21428 9220 21480
rect 9272 21468 9278 21480
rect 9766 21468 9772 21480
rect 9272 21440 9772 21468
rect 9272 21428 9278 21440
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 10134 21468 10140 21480
rect 10095 21440 10140 21468
rect 10134 21428 10140 21440
rect 10192 21428 10198 21480
rect 1903 21372 5580 21400
rect 7745 21403 7803 21409
rect 1903 21369 1915 21372
rect 1857 21363 1915 21369
rect 7745 21369 7757 21403
rect 7791 21400 7803 21403
rect 12250 21400 12256 21412
rect 7791 21372 12256 21400
rect 7791 21369 7803 21372
rect 7745 21363 7803 21369
rect 12250 21360 12256 21372
rect 12308 21360 12314 21412
rect 13004 21344 13032 21506
rect 13081 21505 13093 21506
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 16853 21539 16911 21545
rect 16853 21505 16865 21539
rect 16899 21536 16911 21539
rect 16942 21536 16948 21548
rect 16899 21508 16948 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17678 21536 17684 21548
rect 17591 21508 17684 21536
rect 17678 21496 17684 21508
rect 17736 21536 17742 21548
rect 19168 21536 19196 21576
rect 21269 21573 21281 21576
rect 21315 21604 21327 21607
rect 28902 21604 28908 21616
rect 21315 21576 24992 21604
rect 21315 21573 21327 21576
rect 21269 21567 21327 21573
rect 17736 21508 19196 21536
rect 20993 21539 21051 21545
rect 17736 21496 17742 21508
rect 20993 21505 21005 21539
rect 21039 21536 21051 21539
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21039 21508 22017 21536
rect 21039 21505 21051 21508
rect 20993 21499 21051 21505
rect 22005 21505 22017 21508
rect 22051 21536 22063 21539
rect 22186 21536 22192 21548
rect 22051 21508 22192 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22186 21496 22192 21508
rect 22244 21496 22250 21548
rect 24964 21545 24992 21576
rect 25608 21576 28908 21604
rect 25608 21545 25636 21576
rect 28902 21564 28908 21576
rect 28960 21564 28966 21616
rect 33318 21604 33324 21616
rect 33279 21576 33324 21604
rect 33318 21564 33324 21576
rect 33376 21564 33382 21616
rect 34054 21564 34060 21616
rect 34112 21604 34118 21616
rect 35820 21604 35848 21644
rect 36633 21641 36645 21644
rect 36679 21641 36691 21675
rect 37550 21672 37556 21684
rect 37511 21644 37556 21672
rect 36633 21635 36691 21641
rect 37550 21632 37556 21644
rect 37608 21632 37614 21684
rect 34112 21576 35848 21604
rect 34112 21564 34118 21576
rect 36354 21564 36360 21616
rect 36412 21604 36418 21616
rect 38197 21607 38255 21613
rect 38197 21604 38209 21607
rect 36412 21576 38209 21604
rect 36412 21564 36418 21576
rect 38197 21573 38209 21576
rect 38243 21573 38255 21607
rect 38197 21567 38255 21573
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 25593 21539 25651 21545
rect 25593 21505 25605 21539
rect 25639 21505 25651 21539
rect 30377 21539 30435 21545
rect 30377 21536 30389 21539
rect 25593 21499 25651 21505
rect 28920 21508 30389 21536
rect 15838 21428 15844 21480
rect 15896 21468 15902 21480
rect 19978 21468 19984 21480
rect 15896 21440 19984 21468
rect 15896 21428 15902 21440
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 22646 21428 22652 21480
rect 22704 21468 22710 21480
rect 22830 21468 22836 21480
rect 22704 21440 22836 21468
rect 22704 21428 22710 21440
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 24964 21468 24992 21499
rect 28920 21480 28948 21508
rect 30377 21505 30389 21508
rect 30423 21536 30435 21539
rect 31018 21536 31024 21548
rect 30423 21508 31024 21536
rect 30423 21505 30435 21508
rect 30377 21499 30435 21505
rect 31018 21496 31024 21508
rect 31076 21496 31082 21548
rect 31202 21496 31208 21548
rect 31260 21536 31266 21548
rect 31573 21539 31631 21545
rect 31573 21536 31585 21539
rect 31260 21508 31585 21536
rect 31260 21496 31266 21508
rect 31573 21505 31585 21508
rect 31619 21505 31631 21539
rect 31573 21499 31631 21505
rect 34146 21496 34152 21548
rect 34204 21536 34210 21548
rect 34701 21539 34759 21545
rect 34701 21536 34713 21539
rect 34204 21508 34713 21536
rect 34204 21496 34210 21508
rect 34701 21505 34713 21508
rect 34747 21505 34759 21539
rect 34701 21499 34759 21505
rect 35621 21539 35679 21545
rect 35621 21505 35633 21539
rect 35667 21505 35679 21539
rect 36538 21536 36544 21548
rect 36499 21508 36544 21536
rect 35621 21499 35679 21505
rect 28902 21468 28908 21480
rect 24964 21440 28908 21468
rect 28902 21428 28908 21440
rect 28960 21428 28966 21480
rect 32674 21428 32680 21480
rect 32732 21468 32738 21480
rect 33229 21471 33287 21477
rect 33229 21468 33241 21471
rect 32732 21440 33241 21468
rect 32732 21428 32738 21440
rect 33229 21437 33241 21440
rect 33275 21437 33287 21471
rect 33229 21431 33287 21437
rect 33505 21471 33563 21477
rect 33505 21437 33517 21471
rect 33551 21468 33563 21471
rect 34974 21468 34980 21480
rect 33551 21440 34980 21468
rect 33551 21437 33563 21440
rect 33505 21431 33563 21437
rect 13446 21360 13452 21412
rect 13504 21400 13510 21412
rect 13504 21372 17908 21400
rect 13504 21360 13510 21372
rect 1946 21292 1952 21344
rect 2004 21332 2010 21344
rect 2317 21335 2375 21341
rect 2317 21332 2329 21335
rect 2004 21304 2329 21332
rect 2004 21292 2010 21304
rect 2317 21301 2329 21304
rect 2363 21301 2375 21335
rect 10686 21332 10692 21344
rect 10647 21304 10692 21332
rect 2317 21295 2375 21301
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 12437 21335 12495 21341
rect 12437 21301 12449 21335
rect 12483 21332 12495 21335
rect 12526 21332 12532 21344
rect 12483 21304 12532 21332
rect 12483 21301 12495 21304
rect 12437 21295 12495 21301
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 12986 21292 12992 21344
rect 13044 21292 13050 21344
rect 16945 21335 17003 21341
rect 16945 21301 16957 21335
rect 16991 21332 17003 21335
rect 17126 21332 17132 21344
rect 16991 21304 17132 21332
rect 16991 21301 17003 21304
rect 16945 21295 17003 21301
rect 17126 21292 17132 21304
rect 17184 21292 17190 21344
rect 17880 21332 17908 21372
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 26234 21400 26240 21412
rect 19208 21372 26240 21400
rect 19208 21360 19214 21372
rect 26234 21360 26240 21372
rect 26292 21360 26298 21412
rect 30466 21360 30472 21412
rect 30524 21400 30530 21412
rect 33520 21400 33548 21431
rect 34974 21428 34980 21440
rect 35032 21428 35038 21480
rect 35636 21400 35664 21499
rect 36538 21496 36544 21508
rect 36596 21536 36602 21548
rect 37090 21536 37096 21548
rect 36596 21508 37096 21536
rect 36596 21496 36602 21508
rect 37090 21496 37096 21508
rect 37148 21496 37154 21548
rect 37182 21496 37188 21548
rect 37240 21536 37246 21548
rect 37461 21539 37519 21545
rect 37461 21536 37473 21539
rect 37240 21508 37473 21536
rect 37240 21496 37246 21508
rect 37461 21505 37473 21508
rect 37507 21505 37519 21539
rect 37461 21499 37519 21505
rect 38105 21539 38163 21545
rect 38105 21505 38117 21539
rect 38151 21505 38163 21539
rect 38105 21499 38163 21505
rect 37108 21468 37136 21496
rect 38120 21468 38148 21499
rect 37108 21440 38148 21468
rect 30524 21372 33548 21400
rect 33612 21372 35664 21400
rect 30524 21360 30530 21372
rect 22370 21332 22376 21344
rect 17880 21304 22376 21332
rect 22370 21292 22376 21304
rect 22428 21332 22434 21344
rect 23198 21332 23204 21344
rect 22428 21304 23204 21332
rect 22428 21292 22434 21304
rect 23198 21292 23204 21304
rect 23256 21292 23262 21344
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 25685 21335 25743 21341
rect 25685 21332 25697 21335
rect 25188 21304 25697 21332
rect 25188 21292 25194 21304
rect 25685 21301 25697 21304
rect 25731 21301 25743 21335
rect 25685 21295 25743 21301
rect 31938 21292 31944 21344
rect 31996 21332 32002 21344
rect 33612 21332 33640 21372
rect 31996 21304 33640 21332
rect 31996 21292 32002 21304
rect 34514 21292 34520 21344
rect 34572 21332 34578 21344
rect 34701 21335 34759 21341
rect 34701 21332 34713 21335
rect 34572 21304 34713 21332
rect 34572 21292 34578 21304
rect 34701 21301 34713 21304
rect 34747 21301 34759 21335
rect 34701 21295 34759 21301
rect 34882 21292 34888 21344
rect 34940 21332 34946 21344
rect 35526 21332 35532 21344
rect 34940 21304 35532 21332
rect 34940 21292 34946 21304
rect 35526 21292 35532 21304
rect 35584 21292 35590 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1765 21131 1823 21137
rect 1765 21097 1777 21131
rect 1811 21128 1823 21131
rect 10870 21128 10876 21140
rect 1811 21100 10876 21128
rect 1811 21097 1823 21100
rect 1765 21091 1823 21097
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 14734 21128 14740 21140
rect 12308 21100 14740 21128
rect 12308 21088 12314 21100
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 17034 21128 17040 21140
rect 15252 21100 17040 21128
rect 15252 21088 15258 21100
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 18141 21131 18199 21137
rect 18141 21097 18153 21131
rect 18187 21128 18199 21131
rect 19334 21128 19340 21140
rect 18187 21100 19340 21128
rect 18187 21097 18199 21100
rect 18141 21091 18199 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 19426 21088 19432 21140
rect 19484 21128 19490 21140
rect 19521 21131 19579 21137
rect 19521 21128 19533 21131
rect 19484 21100 19533 21128
rect 19484 21088 19490 21100
rect 19521 21097 19533 21100
rect 19567 21097 19579 21131
rect 21174 21128 21180 21140
rect 21135 21100 21180 21128
rect 19521 21091 19579 21097
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 28997 21131 29055 21137
rect 28997 21097 29009 21131
rect 29043 21128 29055 21131
rect 29086 21128 29092 21140
rect 29043 21100 29092 21128
rect 29043 21097 29055 21100
rect 28997 21091 29055 21097
rect 29086 21088 29092 21100
rect 29144 21088 29150 21140
rect 29822 21128 29828 21140
rect 29783 21100 29828 21128
rect 29822 21088 29828 21100
rect 29880 21088 29886 21140
rect 30742 21128 30748 21140
rect 30703 21100 30748 21128
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 31846 21088 31852 21140
rect 31904 21128 31910 21140
rect 32033 21131 32091 21137
rect 32033 21128 32045 21131
rect 31904 21100 32045 21128
rect 31904 21088 31910 21100
rect 32033 21097 32045 21100
rect 32079 21097 32091 21131
rect 34146 21128 34152 21140
rect 34107 21100 34152 21128
rect 32033 21091 32091 21097
rect 34146 21088 34152 21100
rect 34204 21088 34210 21140
rect 34790 21088 34796 21140
rect 34848 21128 34854 21140
rect 36541 21131 36599 21137
rect 36541 21128 36553 21131
rect 34848 21100 36553 21128
rect 34848 21088 34854 21100
rect 36541 21097 36553 21100
rect 36587 21097 36599 21131
rect 36541 21091 36599 21097
rect 37366 21088 37372 21140
rect 37424 21128 37430 21140
rect 37829 21131 37887 21137
rect 37829 21128 37841 21131
rect 37424 21100 37841 21128
rect 37424 21088 37430 21100
rect 37829 21097 37841 21100
rect 37875 21097 37887 21131
rect 37829 21091 37887 21097
rect 12618 21020 12624 21072
rect 12676 21060 12682 21072
rect 12676 21032 19564 21060
rect 12676 21020 12682 21032
rect 8113 20995 8171 21001
rect 8113 20961 8125 20995
rect 8159 20992 8171 20995
rect 8478 20992 8484 21004
rect 8159 20964 8484 20992
rect 8159 20961 8171 20964
rect 8113 20955 8171 20961
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 10226 20992 10232 21004
rect 9600 20964 10232 20992
rect 1670 20856 1676 20868
rect 1631 20828 1676 20856
rect 1670 20816 1676 20828
rect 1728 20816 1734 20868
rect 7466 20856 7472 20868
rect 7427 20828 7472 20856
rect 7466 20816 7472 20828
rect 7524 20816 7530 20868
rect 7558 20816 7564 20868
rect 7616 20856 7622 20868
rect 7616 20828 7661 20856
rect 7616 20816 7622 20828
rect 9122 20816 9128 20868
rect 9180 20856 9186 20868
rect 9600 20856 9628 20964
rect 10226 20952 10232 20964
rect 10284 20952 10290 21004
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 10376 20964 10421 20992
rect 10376 20952 10382 20964
rect 10594 20952 10600 21004
rect 10652 20992 10658 21004
rect 11333 20995 11391 21001
rect 11333 20992 11345 20995
rect 10652 20964 11345 20992
rect 10652 20952 10658 20964
rect 11333 20961 11345 20964
rect 11379 20961 11391 20995
rect 11333 20955 11391 20961
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 15028 21001 15240 21004
rect 15028 20995 15255 21001
rect 15028 20992 15209 20995
rect 11848 20976 15209 20992
rect 11848 20964 15056 20976
rect 11848 20952 11854 20964
rect 15197 20961 15209 20976
rect 15243 20961 15255 20995
rect 15378 20992 15384 21004
rect 15339 20964 15384 20992
rect 15197 20955 15255 20961
rect 15378 20952 15384 20964
rect 15436 20952 15442 21004
rect 11054 20884 11060 20936
rect 11112 20924 11118 20936
rect 11241 20927 11299 20933
rect 11241 20924 11253 20927
rect 11112 20896 11253 20924
rect 11112 20884 11118 20896
rect 11241 20893 11253 20896
rect 11287 20893 11299 20927
rect 11241 20887 11299 20893
rect 11422 20884 11428 20936
rect 11480 20924 11486 20936
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 11480 20896 12173 20924
rect 11480 20884 11486 20896
rect 12161 20893 12173 20896
rect 12207 20893 12219 20927
rect 12161 20887 12219 20893
rect 13081 20927 13139 20933
rect 13081 20893 13093 20927
rect 13127 20924 13139 20927
rect 13446 20924 13452 20936
rect 13127 20896 13452 20924
rect 13127 20893 13139 20896
rect 13081 20887 13139 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20924 13599 20927
rect 14366 20924 14372 20936
rect 13587 20896 14372 20924
rect 13587 20893 13599 20896
rect 13541 20887 13599 20893
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20893 14611 20927
rect 14553 20887 14611 20893
rect 9769 20859 9827 20865
rect 9769 20856 9781 20859
rect 9180 20828 9781 20856
rect 9180 20816 9186 20828
rect 9769 20825 9781 20828
rect 9815 20825 9827 20859
rect 9769 20819 9827 20825
rect 9861 20859 9919 20865
rect 9861 20825 9873 20859
rect 9907 20825 9919 20859
rect 13633 20859 13691 20865
rect 13633 20856 13645 20859
rect 9861 20819 9919 20825
rect 11164 20828 13645 20856
rect 9876 20788 9904 20819
rect 11164 20788 11192 20828
rect 13633 20825 13645 20828
rect 13679 20825 13691 20859
rect 13633 20819 13691 20825
rect 12250 20788 12256 20800
rect 9876 20760 11192 20788
rect 12211 20760 12256 20788
rect 12250 20748 12256 20760
rect 12308 20748 12314 20800
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 12897 20791 12955 20797
rect 12897 20788 12909 20791
rect 12676 20760 12909 20788
rect 12676 20748 12682 20760
rect 12897 20757 12909 20760
rect 12943 20757 12955 20791
rect 12897 20751 12955 20757
rect 12986 20748 12992 20800
rect 13044 20788 13050 20800
rect 14090 20788 14096 20800
rect 13044 20760 14096 20788
rect 13044 20748 13050 20760
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 14568 20788 14596 20887
rect 14642 20884 14648 20936
rect 14700 20924 14706 20936
rect 18046 20924 18052 20936
rect 14700 20896 14745 20924
rect 18007 20896 18052 20924
rect 14700 20884 14706 20896
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 18690 20924 18696 20936
rect 18651 20896 18696 20924
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19300 20896 19441 20924
rect 19300 20884 19306 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19536 20924 19564 21032
rect 21082 21020 21088 21072
rect 21140 21060 21146 21072
rect 23385 21063 23443 21069
rect 23385 21060 23397 21063
rect 21140 21032 23397 21060
rect 21140 21020 21146 21032
rect 23385 21029 23397 21032
rect 23431 21029 23443 21063
rect 26418 21060 26424 21072
rect 23385 21023 23443 21029
rect 23492 21032 26424 21060
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 20496 20964 21680 20992
rect 20496 20952 20502 20964
rect 21358 20924 21364 20936
rect 19536 20896 21364 20924
rect 19429 20887 19487 20893
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 17034 20856 17040 20868
rect 16995 20828 17040 20856
rect 17034 20816 17040 20828
rect 17092 20816 17098 20868
rect 17218 20816 17224 20868
rect 17276 20856 17282 20868
rect 21266 20856 21272 20868
rect 17276 20828 21272 20856
rect 17276 20816 17282 20828
rect 21266 20816 21272 20828
rect 21324 20816 21330 20868
rect 17862 20788 17868 20800
rect 14568 20760 17868 20788
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 18785 20791 18843 20797
rect 18785 20757 18797 20791
rect 18831 20788 18843 20791
rect 21542 20788 21548 20800
rect 18831 20760 21548 20788
rect 18831 20757 18843 20760
rect 18785 20751 18843 20757
rect 21542 20748 21548 20760
rect 21600 20748 21606 20800
rect 21652 20788 21680 20964
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 22097 20995 22155 21001
rect 22097 20992 22109 20995
rect 22060 20964 22109 20992
rect 22060 20952 22066 20964
rect 22097 20961 22109 20964
rect 22143 20992 22155 20995
rect 23492 20992 23520 21032
rect 26418 21020 26424 21032
rect 26476 21020 26482 21072
rect 33410 21060 33416 21072
rect 31312 21032 33416 21060
rect 22143 20964 23520 20992
rect 22143 20961 22155 20964
rect 22097 20955 22155 20961
rect 23934 20952 23940 21004
rect 23992 20992 23998 21004
rect 30466 20992 30472 21004
rect 23992 20964 30472 20992
rect 23992 20952 23998 20964
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20924 21879 20927
rect 22186 20924 22192 20936
rect 21867 20896 22192 20924
rect 21867 20893 21879 20896
rect 21821 20887 21879 20893
rect 22186 20884 22192 20896
rect 22244 20924 22250 20936
rect 22646 20924 22652 20936
rect 22244 20896 22652 20924
rect 22244 20884 22250 20896
rect 22646 20884 22652 20896
rect 22704 20884 22710 20936
rect 23290 20924 23296 20936
rect 23251 20896 23296 20924
rect 23290 20884 23296 20896
rect 23348 20884 23354 20936
rect 26050 20884 26056 20936
rect 26108 20924 26114 20936
rect 26237 20927 26295 20933
rect 26237 20924 26249 20927
rect 26108 20896 26249 20924
rect 26108 20884 26114 20896
rect 26237 20893 26249 20896
rect 26283 20893 26295 20927
rect 26237 20887 26295 20893
rect 26326 20884 26332 20936
rect 26384 20924 26390 20936
rect 27157 20927 27215 20933
rect 27157 20924 27169 20927
rect 26384 20896 27169 20924
rect 26384 20884 26390 20896
rect 27157 20893 27169 20896
rect 27203 20893 27215 20927
rect 28902 20924 28908 20936
rect 28863 20896 28908 20924
rect 27157 20887 27215 20893
rect 28902 20884 28908 20896
rect 28960 20884 28966 20936
rect 29730 20924 29736 20936
rect 29691 20896 29736 20924
rect 29730 20884 29736 20896
rect 29788 20924 29794 20936
rect 31312 20933 31340 21032
rect 33410 21020 33416 21032
rect 33468 21020 33474 21072
rect 33778 21020 33784 21072
rect 33836 21060 33842 21072
rect 37185 21063 37243 21069
rect 37185 21060 37197 21063
rect 33836 21032 37197 21060
rect 33836 21020 33842 21032
rect 37185 21029 37197 21032
rect 37231 21029 37243 21063
rect 37185 21023 37243 21029
rect 31389 20995 31447 21001
rect 31389 20961 31401 20995
rect 31435 20992 31447 20995
rect 33134 20992 33140 21004
rect 31435 20964 33140 20992
rect 31435 20961 31447 20964
rect 31389 20955 31447 20961
rect 33134 20952 33140 20964
rect 33192 20952 33198 21004
rect 34790 20952 34796 21004
rect 34848 20952 34854 21004
rect 35250 20992 35256 21004
rect 35211 20964 35256 20992
rect 35250 20952 35256 20964
rect 35308 20992 35314 21004
rect 35434 20992 35440 21004
rect 35308 20964 35440 20992
rect 35308 20952 35314 20964
rect 35434 20952 35440 20964
rect 35492 20952 35498 21004
rect 30653 20927 30711 20933
rect 30653 20924 30665 20927
rect 29788 20896 30665 20924
rect 29788 20884 29794 20896
rect 30653 20893 30665 20896
rect 30699 20893 30711 20927
rect 30653 20887 30711 20893
rect 31297 20927 31355 20933
rect 31297 20893 31309 20927
rect 31343 20893 31355 20927
rect 31938 20924 31944 20936
rect 31297 20887 31355 20893
rect 31726 20896 31944 20924
rect 24486 20816 24492 20868
rect 24544 20856 24550 20868
rect 24673 20859 24731 20865
rect 24673 20856 24685 20859
rect 24544 20828 24685 20856
rect 24544 20816 24550 20828
rect 24673 20825 24685 20828
rect 24719 20825 24731 20859
rect 24673 20819 24731 20825
rect 24765 20859 24823 20865
rect 24765 20825 24777 20859
rect 24811 20856 24823 20859
rect 25130 20856 25136 20868
rect 24811 20828 25136 20856
rect 24811 20825 24823 20828
rect 24765 20819 24823 20825
rect 25130 20816 25136 20828
rect 25188 20816 25194 20868
rect 25685 20859 25743 20865
rect 25685 20825 25697 20859
rect 25731 20856 25743 20859
rect 25774 20856 25780 20868
rect 25731 20828 25780 20856
rect 25731 20825 25743 20828
rect 25685 20819 25743 20825
rect 25774 20816 25780 20828
rect 25832 20816 25838 20868
rect 25866 20816 25872 20868
rect 25924 20856 25930 20868
rect 26513 20859 26571 20865
rect 26513 20856 26525 20859
rect 25924 20828 26525 20856
rect 25924 20816 25930 20828
rect 26513 20825 26525 20828
rect 26559 20856 26571 20859
rect 27890 20856 27896 20868
rect 26559 20828 27896 20856
rect 26559 20825 26571 20828
rect 26513 20819 26571 20825
rect 27890 20816 27896 20828
rect 27948 20816 27954 20868
rect 30668 20856 30696 20887
rect 31726 20856 31754 20896
rect 31938 20884 31944 20896
rect 31996 20884 32002 20936
rect 34333 20927 34391 20933
rect 34333 20893 34345 20927
rect 34379 20924 34391 20927
rect 34606 20924 34612 20936
rect 34379 20896 34612 20924
rect 34379 20893 34391 20896
rect 34333 20887 34391 20893
rect 34606 20884 34612 20896
rect 34664 20884 34670 20936
rect 32674 20856 32680 20868
rect 30668 20828 31754 20856
rect 31956 20828 32168 20856
rect 32635 20828 32680 20856
rect 25884 20788 25912 20816
rect 21652 20760 25912 20788
rect 27249 20791 27307 20797
rect 27249 20757 27261 20791
rect 27295 20788 27307 20791
rect 29914 20788 29920 20800
rect 27295 20760 29920 20788
rect 27295 20757 27307 20760
rect 27249 20751 27307 20757
rect 29914 20748 29920 20760
rect 29972 20748 29978 20800
rect 30006 20748 30012 20800
rect 30064 20788 30070 20800
rect 31956 20788 31984 20828
rect 30064 20760 31984 20788
rect 32140 20788 32168 20828
rect 32674 20816 32680 20828
rect 32732 20816 32738 20868
rect 32769 20859 32827 20865
rect 32769 20825 32781 20859
rect 32815 20825 32827 20859
rect 32769 20819 32827 20825
rect 33321 20859 33379 20865
rect 33321 20825 33333 20859
rect 33367 20856 33379 20859
rect 34054 20856 34060 20868
rect 33367 20828 34060 20856
rect 33367 20825 33379 20828
rect 33321 20819 33379 20825
rect 32784 20788 32812 20819
rect 34054 20816 34060 20828
rect 34112 20816 34118 20868
rect 34808 20856 34836 20952
rect 36446 20924 36452 20936
rect 36407 20896 36452 20924
rect 36446 20884 36452 20896
rect 36504 20884 36510 20936
rect 36538 20884 36544 20936
rect 36596 20924 36602 20936
rect 37093 20927 37151 20933
rect 37093 20924 37105 20927
rect 36596 20896 37105 20924
rect 36596 20884 36602 20896
rect 37093 20893 37105 20896
rect 37139 20924 37151 20927
rect 37737 20927 37795 20933
rect 37737 20924 37749 20927
rect 37139 20896 37749 20924
rect 37139 20893 37151 20896
rect 37093 20887 37151 20893
rect 37737 20893 37749 20896
rect 37783 20893 37795 20927
rect 37737 20887 37795 20893
rect 34977 20859 35035 20865
rect 34977 20856 34989 20859
rect 34808 20828 34989 20856
rect 34977 20825 34989 20828
rect 35023 20825 35035 20859
rect 34977 20819 35035 20825
rect 35069 20859 35127 20865
rect 35069 20825 35081 20859
rect 35115 20825 35127 20859
rect 35069 20819 35127 20825
rect 32140 20760 32812 20788
rect 30064 20748 30070 20760
rect 34698 20748 34704 20800
rect 34756 20788 34762 20800
rect 35084 20788 35112 20819
rect 34756 20760 35112 20788
rect 34756 20748 34762 20760
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 1765 20587 1823 20593
rect 1765 20553 1777 20587
rect 1811 20584 1823 20587
rect 1854 20584 1860 20596
rect 1811 20556 1860 20584
rect 1811 20553 1823 20556
rect 1765 20547 1823 20553
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 5408 20556 12112 20584
rect 5408 20544 5414 20556
rect 6638 20476 6644 20528
rect 6696 20516 6702 20528
rect 6733 20519 6791 20525
rect 6733 20516 6745 20519
rect 6696 20488 6745 20516
rect 6696 20476 6702 20488
rect 6733 20485 6745 20488
rect 6779 20485 6791 20519
rect 6733 20479 6791 20485
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 11790 20516 11796 20528
rect 10008 20488 11796 20516
rect 10008 20476 10014 20488
rect 1854 20408 1860 20460
rect 1912 20448 1918 20460
rect 1949 20451 2007 20457
rect 1949 20448 1961 20451
rect 1912 20420 1961 20448
rect 1912 20408 1918 20420
rect 1949 20417 1961 20420
rect 1995 20417 2007 20451
rect 1949 20411 2007 20417
rect 7834 20408 7840 20460
rect 7892 20448 7898 20460
rect 10244 20457 10272 20488
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 8021 20451 8079 20457
rect 8021 20448 8033 20451
rect 7892 20420 8033 20448
rect 7892 20408 7898 20420
rect 8021 20417 8033 20420
rect 8067 20417 8079 20451
rect 8021 20411 8079 20417
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20448 10471 20451
rect 10686 20448 10692 20460
rect 10459 20420 10692 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 5626 20340 5632 20392
rect 5684 20380 5690 20392
rect 6641 20383 6699 20389
rect 6641 20380 6653 20383
rect 5684 20352 6653 20380
rect 5684 20340 5690 20352
rect 6641 20349 6653 20352
rect 6687 20349 6699 20383
rect 7282 20380 7288 20392
rect 7243 20352 7288 20380
rect 6641 20343 6699 20349
rect 7282 20340 7288 20352
rect 7340 20340 7346 20392
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20380 9643 20383
rect 10042 20380 10048 20392
rect 9631 20352 10048 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 12084 20380 12112 20556
rect 12158 20544 12164 20596
rect 12216 20584 12222 20596
rect 12345 20587 12403 20593
rect 12345 20584 12357 20587
rect 12216 20556 12357 20584
rect 12216 20544 12222 20556
rect 12345 20553 12357 20556
rect 12391 20553 12403 20587
rect 16390 20584 16396 20596
rect 12345 20547 12403 20553
rect 12452 20556 16396 20584
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12452 20448 12480 20556
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 17497 20587 17555 20593
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 18230 20584 18236 20596
rect 17543 20556 18236 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 18230 20544 18236 20556
rect 18288 20544 18294 20596
rect 18874 20584 18880 20596
rect 18835 20556 18880 20584
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 22830 20584 22836 20596
rect 19812 20556 22836 20584
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 13170 20516 13176 20528
rect 12860 20488 13176 20516
rect 12860 20476 12866 20488
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 13449 20519 13507 20525
rect 13449 20485 13461 20519
rect 13495 20516 13507 20519
rect 14550 20516 14556 20528
rect 13495 20488 14556 20516
rect 13495 20485 13507 20488
rect 13449 20479 13507 20485
rect 14550 20476 14556 20488
rect 14608 20476 14614 20528
rect 14734 20476 14740 20528
rect 14792 20516 14798 20528
rect 15289 20519 15347 20525
rect 15289 20516 15301 20519
rect 14792 20488 15301 20516
rect 14792 20476 14798 20488
rect 15289 20485 15301 20488
rect 15335 20485 15347 20519
rect 15289 20479 15347 20485
rect 15381 20519 15439 20525
rect 15381 20485 15393 20519
rect 15427 20516 15439 20519
rect 16758 20516 16764 20528
rect 15427 20488 16764 20516
rect 15427 20485 15439 20488
rect 15381 20479 15439 20485
rect 16758 20476 16764 20488
rect 16816 20476 16822 20528
rect 17586 20476 17592 20528
rect 17644 20516 17650 20528
rect 19812 20516 19840 20556
rect 22830 20544 22836 20556
rect 22888 20584 22894 20596
rect 23382 20584 23388 20596
rect 22888 20556 23388 20584
rect 22888 20544 22894 20556
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 25406 20584 25412 20596
rect 24596 20556 25412 20584
rect 17644 20488 19840 20516
rect 17644 20476 17650 20488
rect 20990 20476 20996 20528
rect 21048 20516 21054 20528
rect 22925 20519 22983 20525
rect 22925 20516 22937 20519
rect 21048 20488 22937 20516
rect 21048 20476 21054 20488
rect 22925 20485 22937 20488
rect 22971 20485 22983 20519
rect 22925 20479 22983 20485
rect 23017 20519 23075 20525
rect 23017 20485 23029 20519
rect 23063 20516 23075 20519
rect 23566 20516 23572 20528
rect 23063 20488 23572 20516
rect 23063 20485 23075 20488
rect 23017 20479 23075 20485
rect 23566 20476 23572 20488
rect 23624 20476 23630 20528
rect 23934 20476 23940 20528
rect 23992 20516 23998 20528
rect 23992 20488 24037 20516
rect 23992 20476 23998 20488
rect 17405 20451 17463 20457
rect 12299 20420 12480 20448
rect 12544 20420 13216 20448
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12544 20380 12572 20420
rect 12802 20380 12808 20392
rect 12084 20352 12572 20380
rect 12636 20352 12808 20380
rect 7742 20272 7748 20324
rect 7800 20312 7806 20324
rect 10870 20312 10876 20324
rect 7800 20284 8892 20312
rect 10783 20284 10876 20312
rect 7800 20272 7806 20284
rect 5074 20204 5080 20256
rect 5132 20244 5138 20256
rect 8018 20244 8024 20256
rect 5132 20216 8024 20244
rect 5132 20204 5138 20216
rect 8018 20204 8024 20216
rect 8076 20204 8082 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8754 20244 8760 20256
rect 8159 20216 8760 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 8864 20244 8892 20284
rect 10870 20272 10876 20284
rect 10928 20312 10934 20324
rect 12636 20312 12664 20352
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 10928 20284 12664 20312
rect 13188 20312 13216 20420
rect 17405 20417 17417 20451
rect 17451 20448 17463 20451
rect 17678 20448 17684 20460
rect 17451 20420 17684 20448
rect 17451 20417 17463 20420
rect 17405 20411 17463 20417
rect 17678 20408 17684 20420
rect 17736 20408 17742 20460
rect 18046 20408 18052 20460
rect 18104 20448 18110 20460
rect 18141 20451 18199 20457
rect 18141 20448 18153 20451
rect 18104 20420 18153 20448
rect 18104 20408 18110 20420
rect 18141 20417 18153 20420
rect 18187 20417 18199 20451
rect 18141 20411 18199 20417
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20448 18843 20451
rect 22002 20448 22008 20460
rect 18831 20420 22008 20448
rect 18831 20417 18843 20420
rect 18785 20411 18843 20417
rect 13357 20383 13415 20389
rect 13357 20349 13369 20383
rect 13403 20380 13415 20383
rect 13446 20380 13452 20392
rect 13403 20352 13452 20380
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 14366 20380 14372 20392
rect 14327 20352 14372 20380
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20349 15623 20383
rect 18156 20380 18184 20411
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 24118 20408 24124 20460
rect 24176 20448 24182 20460
rect 24596 20448 24624 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 25682 20544 25688 20596
rect 25740 20584 25746 20596
rect 25777 20587 25835 20593
rect 25777 20584 25789 20587
rect 25740 20556 25789 20584
rect 25740 20544 25746 20556
rect 25777 20553 25789 20556
rect 25823 20553 25835 20587
rect 25777 20547 25835 20553
rect 26510 20544 26516 20596
rect 26568 20584 26574 20596
rect 27154 20584 27160 20596
rect 26568 20556 27160 20584
rect 26568 20544 26574 20556
rect 27154 20544 27160 20556
rect 27212 20544 27218 20596
rect 28166 20544 28172 20596
rect 28224 20584 28230 20596
rect 29181 20587 29239 20593
rect 29181 20584 29193 20587
rect 28224 20556 29193 20584
rect 28224 20544 28230 20556
rect 29181 20553 29193 20556
rect 29227 20553 29239 20587
rect 29181 20547 29239 20553
rect 29730 20544 29736 20596
rect 29788 20584 29794 20596
rect 31110 20584 31116 20596
rect 29788 20556 30512 20584
rect 31071 20556 31116 20584
rect 29788 20544 29794 20556
rect 24670 20476 24676 20528
rect 24728 20516 24734 20528
rect 26421 20519 26479 20525
rect 26421 20516 26433 20519
rect 24728 20488 26433 20516
rect 24728 20476 24734 20488
rect 26421 20485 26433 20488
rect 26467 20485 26479 20519
rect 28534 20516 28540 20528
rect 28495 20488 28540 20516
rect 26421 20479 26479 20485
rect 28534 20476 28540 20488
rect 28592 20476 28598 20528
rect 28626 20476 28632 20528
rect 28684 20516 28690 20528
rect 29825 20519 29883 20525
rect 29825 20516 29837 20519
rect 28684 20488 29837 20516
rect 28684 20476 28690 20488
rect 29825 20485 29837 20488
rect 29871 20485 29883 20519
rect 29825 20479 29883 20485
rect 24765 20451 24823 20457
rect 24765 20448 24777 20451
rect 24176 20420 24777 20448
rect 24176 20408 24182 20420
rect 24765 20417 24777 20420
rect 24811 20417 24823 20451
rect 25682 20448 25688 20460
rect 24765 20411 24823 20417
rect 24872 20420 25688 20448
rect 23198 20380 23204 20392
rect 18156 20352 23204 20380
rect 15565 20343 15623 20349
rect 15580 20312 15608 20343
rect 23198 20340 23204 20352
rect 23256 20340 23262 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 24872 20380 24900 20420
rect 25682 20408 25688 20420
rect 25740 20408 25746 20460
rect 26329 20451 26387 20457
rect 26329 20417 26341 20451
rect 26375 20448 26387 20451
rect 26510 20448 26516 20460
rect 26375 20420 26516 20448
rect 26375 20417 26387 20420
rect 26329 20411 26387 20417
rect 26510 20408 26516 20420
rect 26568 20408 26574 20460
rect 27157 20451 27215 20457
rect 27157 20417 27169 20451
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 28445 20451 28503 20457
rect 28445 20417 28457 20451
rect 28491 20448 28503 20451
rect 28810 20448 28816 20460
rect 28491 20420 28816 20448
rect 28491 20417 28503 20420
rect 28445 20411 28503 20417
rect 23348 20352 24900 20380
rect 25041 20383 25099 20389
rect 23348 20340 23354 20352
rect 25041 20349 25053 20383
rect 25087 20380 25099 20383
rect 25130 20380 25136 20392
rect 25087 20352 25136 20380
rect 25087 20349 25099 20352
rect 25041 20343 25099 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 25406 20340 25412 20392
rect 25464 20380 25470 20392
rect 26050 20380 26056 20392
rect 25464 20352 26056 20380
rect 25464 20340 25470 20352
rect 26050 20340 26056 20352
rect 26108 20380 26114 20392
rect 26234 20380 26240 20392
rect 26108 20352 26240 20380
rect 26108 20340 26114 20352
rect 26234 20340 26240 20352
rect 26292 20380 26298 20392
rect 27172 20380 27200 20411
rect 26292 20352 27200 20380
rect 27433 20383 27491 20389
rect 26292 20340 26298 20352
rect 27433 20349 27445 20383
rect 27479 20380 27491 20383
rect 28166 20380 28172 20392
rect 27479 20352 28172 20380
rect 27479 20349 27491 20352
rect 27433 20343 27491 20349
rect 28166 20340 28172 20352
rect 28224 20340 28230 20392
rect 16666 20312 16672 20324
rect 13188 20284 16672 20312
rect 10928 20272 10934 20284
rect 16666 20272 16672 20284
rect 16724 20272 16730 20324
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20312 18291 20315
rect 20806 20312 20812 20324
rect 18279 20284 20812 20312
rect 18279 20281 18291 20284
rect 18233 20275 18291 20281
rect 20806 20272 20812 20284
rect 20864 20272 20870 20324
rect 23014 20272 23020 20324
rect 23072 20312 23078 20324
rect 28460 20312 28488 20411
rect 28810 20408 28816 20420
rect 28868 20448 28874 20460
rect 29089 20451 29147 20457
rect 29089 20448 29101 20451
rect 28868 20420 29101 20448
rect 28868 20408 28874 20420
rect 29089 20417 29101 20420
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 29454 20408 29460 20460
rect 29512 20448 29518 20460
rect 29733 20451 29791 20457
rect 29733 20448 29745 20451
rect 29512 20420 29745 20448
rect 29512 20408 29518 20420
rect 29733 20417 29745 20420
rect 29779 20417 29791 20451
rect 30374 20448 30380 20460
rect 30335 20420 30380 20448
rect 29733 20411 29791 20417
rect 30374 20408 30380 20420
rect 30432 20408 30438 20460
rect 30484 20448 30512 20556
rect 31110 20544 31116 20556
rect 31168 20544 31174 20596
rect 32582 20544 32588 20596
rect 32640 20584 32646 20596
rect 33045 20587 33103 20593
rect 33045 20584 33057 20587
rect 32640 20556 33057 20584
rect 32640 20544 32646 20556
rect 33045 20553 33057 20556
rect 33091 20553 33103 20587
rect 33045 20547 33103 20553
rect 33134 20544 33140 20596
rect 33192 20584 33198 20596
rect 35713 20587 35771 20593
rect 33192 20556 34652 20584
rect 33192 20544 33198 20556
rect 31938 20476 31944 20528
rect 31996 20516 32002 20528
rect 32401 20519 32459 20525
rect 32401 20516 32413 20519
rect 31996 20488 32413 20516
rect 31996 20476 32002 20488
rect 32401 20485 32413 20488
rect 32447 20485 32459 20519
rect 34514 20516 34520 20528
rect 34475 20488 34520 20516
rect 32401 20479 32459 20485
rect 34514 20476 34520 20488
rect 34572 20476 34578 20528
rect 34624 20525 34652 20556
rect 35713 20553 35725 20587
rect 35759 20584 35771 20587
rect 35894 20584 35900 20596
rect 35759 20556 35900 20584
rect 35759 20553 35771 20556
rect 35713 20547 35771 20553
rect 35894 20544 35900 20556
rect 35952 20544 35958 20596
rect 36078 20544 36084 20596
rect 36136 20584 36142 20596
rect 36357 20587 36415 20593
rect 36357 20584 36369 20587
rect 36136 20556 36369 20584
rect 36136 20544 36142 20556
rect 36357 20553 36369 20556
rect 36403 20553 36415 20587
rect 36357 20547 36415 20553
rect 37274 20544 37280 20596
rect 37332 20584 37338 20596
rect 37553 20587 37611 20593
rect 37553 20584 37565 20587
rect 37332 20556 37565 20584
rect 37332 20544 37338 20556
rect 37553 20553 37565 20556
rect 37599 20553 37611 20587
rect 37553 20547 37611 20553
rect 37734 20544 37740 20596
rect 37792 20584 37798 20596
rect 38197 20587 38255 20593
rect 38197 20584 38209 20587
rect 37792 20556 38209 20584
rect 37792 20544 37798 20556
rect 38197 20553 38209 20556
rect 38243 20553 38255 20587
rect 38197 20547 38255 20553
rect 34609 20519 34667 20525
rect 34609 20485 34621 20519
rect 34655 20485 34667 20519
rect 34609 20479 34667 20485
rect 31021 20451 31079 20457
rect 31021 20448 31033 20451
rect 30484 20420 31033 20448
rect 31021 20417 31033 20420
rect 31067 20417 31079 20451
rect 32309 20451 32367 20457
rect 32309 20448 32321 20451
rect 31021 20411 31079 20417
rect 31726 20420 32321 20448
rect 28902 20340 28908 20392
rect 28960 20380 28966 20392
rect 31726 20380 31754 20420
rect 32309 20417 32321 20420
rect 32355 20448 32367 20451
rect 32953 20451 33011 20457
rect 32953 20448 32965 20451
rect 32355 20420 32965 20448
rect 32355 20417 32367 20420
rect 32309 20411 32367 20417
rect 32953 20417 32965 20420
rect 32999 20448 33011 20451
rect 33042 20448 33048 20460
rect 32999 20420 33048 20448
rect 32999 20417 33011 20420
rect 32953 20411 33011 20417
rect 33042 20408 33048 20420
rect 33100 20408 33106 20460
rect 33597 20451 33655 20457
rect 33597 20417 33609 20451
rect 33643 20417 33655 20451
rect 33597 20411 33655 20417
rect 35621 20451 35679 20457
rect 35621 20417 35633 20451
rect 35667 20417 35679 20451
rect 36262 20448 36268 20460
rect 36223 20420 36268 20448
rect 35621 20411 35679 20417
rect 28960 20352 31754 20380
rect 33612 20380 33640 20411
rect 35342 20380 35348 20392
rect 33612 20352 35348 20380
rect 28960 20340 28966 20352
rect 35342 20340 35348 20352
rect 35400 20340 35406 20392
rect 23072 20284 28488 20312
rect 23072 20272 23078 20284
rect 31294 20272 31300 20324
rect 31352 20312 31358 20324
rect 35069 20315 35127 20321
rect 31352 20284 35020 20312
rect 31352 20272 31358 20284
rect 18782 20244 18788 20256
rect 8864 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 23382 20204 23388 20256
rect 23440 20244 23446 20256
rect 26418 20244 26424 20256
rect 23440 20216 26424 20244
rect 23440 20204 23446 20216
rect 26418 20204 26424 20216
rect 26476 20204 26482 20256
rect 26510 20204 26516 20256
rect 26568 20244 26574 20256
rect 29730 20244 29736 20256
rect 26568 20216 29736 20244
rect 26568 20204 26574 20216
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 30469 20247 30527 20253
rect 30469 20213 30481 20247
rect 30515 20244 30527 20247
rect 31202 20244 31208 20256
rect 30515 20216 31208 20244
rect 30515 20213 30527 20216
rect 30469 20207 30527 20213
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 33689 20247 33747 20253
rect 33689 20213 33701 20247
rect 33735 20244 33747 20247
rect 34790 20244 34796 20256
rect 33735 20216 34796 20244
rect 33735 20213 33747 20216
rect 33689 20207 33747 20213
rect 34790 20204 34796 20216
rect 34848 20204 34854 20256
rect 34992 20244 35020 20284
rect 35069 20281 35081 20315
rect 35115 20312 35127 20315
rect 35434 20312 35440 20324
rect 35115 20284 35440 20312
rect 35115 20281 35127 20284
rect 35069 20275 35127 20281
rect 35434 20272 35440 20284
rect 35492 20272 35498 20324
rect 35636 20244 35664 20411
rect 36262 20408 36268 20420
rect 36320 20408 36326 20460
rect 37182 20408 37188 20460
rect 37240 20448 37246 20460
rect 37461 20451 37519 20457
rect 37461 20448 37473 20451
rect 37240 20420 37473 20448
rect 37240 20408 37246 20420
rect 37461 20417 37473 20420
rect 37507 20448 37519 20451
rect 38105 20451 38163 20457
rect 38105 20448 38117 20451
rect 37507 20420 38117 20448
rect 37507 20417 37519 20420
rect 37461 20411 37519 20417
rect 38105 20417 38117 20420
rect 38151 20417 38163 20451
rect 38105 20411 38163 20417
rect 36078 20244 36084 20256
rect 34992 20216 36084 20244
rect 36078 20204 36084 20216
rect 36136 20204 36142 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 6638 20040 6644 20052
rect 6599 20012 6644 20040
rect 6638 20000 6644 20012
rect 6696 20000 6702 20052
rect 10229 20043 10287 20049
rect 10229 20009 10241 20043
rect 10275 20040 10287 20043
rect 10870 20040 10876 20052
rect 10275 20012 10876 20040
rect 10275 20009 10287 20012
rect 10229 20003 10287 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 14645 20043 14703 20049
rect 11204 20012 14412 20040
rect 11204 20000 11210 20012
rect 14384 19984 14412 20012
rect 14645 20009 14657 20043
rect 14691 20040 14703 20043
rect 14826 20040 14832 20052
rect 14691 20012 14832 20040
rect 14691 20009 14703 20012
rect 14645 20003 14703 20009
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 16758 20040 16764 20052
rect 16719 20012 16764 20040
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 17402 20040 17408 20052
rect 17363 20012 17408 20040
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 22554 20000 22560 20052
rect 22612 20040 22618 20052
rect 22741 20043 22799 20049
rect 22741 20040 22753 20043
rect 22612 20012 22753 20040
rect 22612 20000 22618 20012
rect 22741 20009 22753 20012
rect 22787 20009 22799 20043
rect 22741 20003 22799 20009
rect 23198 20000 23204 20052
rect 23256 20040 23262 20052
rect 25130 20040 25136 20052
rect 23256 20012 25136 20040
rect 23256 20000 23262 20012
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 27522 20000 27528 20052
rect 27580 20040 27586 20052
rect 27617 20043 27675 20049
rect 27617 20040 27629 20043
rect 27580 20012 27629 20040
rect 27580 20000 27586 20012
rect 27617 20009 27629 20012
rect 27663 20009 27675 20043
rect 28902 20040 28908 20052
rect 28863 20012 28908 20040
rect 27617 20003 27675 20009
rect 28902 20000 28908 20012
rect 28960 20000 28966 20052
rect 31386 20040 31392 20052
rect 31347 20012 31392 20040
rect 31386 20000 31392 20012
rect 31444 20000 31450 20052
rect 32033 20043 32091 20049
rect 32033 20009 32045 20043
rect 32079 20040 32091 20043
rect 32674 20040 32680 20052
rect 32079 20012 32680 20040
rect 32079 20009 32091 20012
rect 32033 20003 32091 20009
rect 32674 20000 32680 20012
rect 32732 20000 32738 20052
rect 33318 20000 33324 20052
rect 33376 20040 33382 20052
rect 33781 20043 33839 20049
rect 33781 20040 33793 20043
rect 33376 20012 33793 20040
rect 33376 20000 33382 20012
rect 33781 20009 33793 20012
rect 33827 20009 33839 20043
rect 33781 20003 33839 20009
rect 34054 20000 34060 20052
rect 34112 20040 34118 20052
rect 35434 20040 35440 20052
rect 34112 20012 35440 20040
rect 34112 20000 34118 20012
rect 35434 20000 35440 20012
rect 35492 20040 35498 20052
rect 35710 20040 35716 20052
rect 35492 20012 35716 20040
rect 35492 20000 35498 20012
rect 35710 20000 35716 20012
rect 35768 20000 35774 20052
rect 36170 20040 36176 20052
rect 36131 20012 36176 20040
rect 36170 20000 36176 20012
rect 36228 20000 36234 20052
rect 36722 20000 36728 20052
rect 36780 20040 36786 20052
rect 36817 20043 36875 20049
rect 36817 20040 36829 20043
rect 36780 20012 36829 20040
rect 36780 20000 36786 20012
rect 36817 20009 36829 20012
rect 36863 20009 36875 20043
rect 36817 20003 36875 20009
rect 37918 20000 37924 20052
rect 37976 20040 37982 20052
rect 38013 20043 38071 20049
rect 38013 20040 38025 20043
rect 37976 20012 38025 20040
rect 37976 20000 37982 20012
rect 38013 20009 38025 20012
rect 38059 20009 38071 20043
rect 38013 20003 38071 20009
rect 5442 19932 5448 19984
rect 5500 19972 5506 19984
rect 8389 19975 8447 19981
rect 8389 19972 8401 19975
rect 5500 19944 8401 19972
rect 5500 19932 5506 19944
rect 8389 19941 8401 19944
rect 8435 19941 8447 19975
rect 8389 19935 8447 19941
rect 10318 19932 10324 19984
rect 10376 19972 10382 19984
rect 10376 19944 14320 19972
rect 10376 19932 10382 19944
rect 1854 19864 1860 19916
rect 1912 19904 1918 19916
rect 1912 19876 7328 19904
rect 1912 19864 1918 19876
rect 6822 19836 6828 19848
rect 6783 19808 6828 19836
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 7300 19845 7328 19876
rect 8018 19864 8024 19916
rect 8076 19904 8082 19916
rect 12066 19904 12072 19916
rect 8076 19876 12072 19904
rect 8076 19864 8082 19876
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 13078 19904 13084 19916
rect 12584 19876 13084 19904
rect 12584 19864 12590 19876
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 13170 19864 13176 19916
rect 13228 19904 13234 19916
rect 13265 19907 13323 19913
rect 13265 19904 13277 19907
rect 13228 19876 13277 19904
rect 13228 19864 13234 19876
rect 13265 19873 13277 19876
rect 13311 19873 13323 19907
rect 14292 19904 14320 19944
rect 14366 19932 14372 19984
rect 14424 19972 14430 19984
rect 20438 19972 20444 19984
rect 14424 19944 20444 19972
rect 14424 19932 14430 19944
rect 20438 19932 20444 19944
rect 20496 19932 20502 19984
rect 21358 19972 21364 19984
rect 21319 19944 21364 19972
rect 21358 19932 21364 19944
rect 21416 19932 21422 19984
rect 27430 19932 27436 19984
rect 27488 19972 27494 19984
rect 28261 19975 28319 19981
rect 28261 19972 28273 19975
rect 27488 19944 28273 19972
rect 27488 19932 27494 19944
rect 28261 19941 28273 19944
rect 28307 19941 28319 19975
rect 28261 19935 28319 19941
rect 28350 19932 28356 19984
rect 28408 19972 28414 19984
rect 29730 19972 29736 19984
rect 28408 19944 29736 19972
rect 28408 19932 28414 19944
rect 29730 19932 29736 19944
rect 29788 19932 29794 19984
rect 31938 19932 31944 19984
rect 31996 19972 32002 19984
rect 34422 19972 34428 19984
rect 31996 19944 34428 19972
rect 31996 19932 32002 19944
rect 34422 19932 34428 19944
rect 34480 19972 34486 19984
rect 36446 19972 36452 19984
rect 34480 19944 36452 19972
rect 34480 19932 34486 19944
rect 36446 19932 36452 19944
rect 36504 19932 36510 19984
rect 37461 19975 37519 19981
rect 37461 19941 37473 19975
rect 37507 19972 37519 19975
rect 39206 19972 39212 19984
rect 37507 19944 39212 19972
rect 37507 19941 37519 19944
rect 37461 19935 37519 19941
rect 39206 19932 39212 19944
rect 39264 19932 39270 19984
rect 16298 19904 16304 19916
rect 14292 19876 16304 19904
rect 13265 19867 13323 19873
rect 16298 19864 16304 19876
rect 16356 19864 16362 19916
rect 19150 19904 19156 19916
rect 16684 19876 19156 19904
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 9398 19836 9404 19848
rect 8619 19808 9404 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 9398 19796 9404 19808
rect 9456 19796 9462 19848
rect 9582 19836 9588 19848
rect 9543 19808 9588 19836
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 9766 19836 9772 19848
rect 9727 19808 9772 19836
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 11333 19839 11391 19845
rect 11333 19805 11345 19839
rect 11379 19836 11391 19839
rect 12618 19836 12624 19848
rect 11379 19808 12624 19836
rect 11379 19805 11391 19808
rect 11333 19799 11391 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 14090 19796 14096 19848
rect 14148 19836 14154 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14148 19808 14565 19836
rect 14148 19796 14154 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19836 15255 19839
rect 15930 19836 15936 19848
rect 15243 19808 15936 19836
rect 15243 19805 15255 19808
rect 15197 19799 15255 19805
rect 1486 19728 1492 19780
rect 1544 19768 1550 19780
rect 11882 19768 11888 19780
rect 1544 19740 11284 19768
rect 11843 19740 11888 19768
rect 1544 19728 1550 19740
rect 7377 19703 7435 19709
rect 7377 19669 7389 19703
rect 7423 19700 7435 19703
rect 9858 19700 9864 19712
rect 7423 19672 9864 19700
rect 7423 19669 7435 19672
rect 7377 19663 7435 19669
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 11146 19700 11152 19712
rect 11107 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11256 19700 11284 19740
rect 11882 19728 11888 19740
rect 11940 19728 11946 19780
rect 12986 19768 12992 19780
rect 12947 19740 12992 19768
rect 12986 19728 12992 19740
rect 13044 19728 13050 19780
rect 13078 19728 13084 19780
rect 13136 19768 13142 19780
rect 14568 19768 14596 19799
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19836 16083 19839
rect 16574 19836 16580 19848
rect 16071 19808 16580 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 16684 19845 16712 19876
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 20809 19907 20867 19913
rect 20809 19873 20821 19907
rect 20855 19904 20867 19907
rect 20990 19904 20996 19916
rect 20855 19876 20996 19904
rect 20855 19873 20867 19876
rect 20809 19867 20867 19873
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 23014 19864 23020 19916
rect 23072 19904 23078 19916
rect 23661 19907 23719 19913
rect 23661 19904 23673 19907
rect 23072 19876 23673 19904
rect 23072 19864 23078 19876
rect 23661 19873 23673 19876
rect 23707 19873 23719 19907
rect 23661 19867 23719 19873
rect 25314 19864 25320 19916
rect 25372 19904 25378 19916
rect 25409 19907 25467 19913
rect 25409 19904 25421 19907
rect 25372 19876 25421 19904
rect 25372 19864 25378 19876
rect 25409 19873 25421 19876
rect 25455 19904 25467 19907
rect 29454 19904 29460 19916
rect 25455 19876 29460 19904
rect 25455 19873 25467 19876
rect 25409 19867 25467 19873
rect 29454 19864 29460 19876
rect 29512 19864 29518 19916
rect 29822 19904 29828 19916
rect 29783 19876 29828 19904
rect 29822 19864 29828 19876
rect 29880 19864 29886 19916
rect 30466 19904 30472 19916
rect 30427 19876 30472 19904
rect 30466 19864 30472 19876
rect 30524 19864 30530 19916
rect 31018 19864 31024 19916
rect 31076 19904 31082 19916
rect 32508 19904 32720 19916
rect 36262 19904 36268 19916
rect 31076 19888 36268 19904
rect 31076 19876 32536 19888
rect 32692 19876 36268 19888
rect 31076 19864 31082 19876
rect 32609 19849 32667 19855
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 17678 19836 17684 19848
rect 17359 19808 17684 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 22649 19839 22707 19845
rect 22649 19805 22661 19839
rect 22695 19836 22707 19839
rect 25133 19839 25191 19845
rect 22695 19808 23244 19836
rect 22695 19805 22707 19808
rect 22649 19799 22707 19805
rect 16758 19768 16764 19780
rect 13136 19740 13181 19768
rect 14568 19740 16764 19768
rect 13136 19728 13142 19740
rect 16758 19728 16764 19740
rect 16816 19768 16822 19780
rect 16942 19768 16948 19780
rect 16816 19740 16948 19768
rect 16816 19728 16822 19740
rect 16942 19728 16948 19740
rect 17000 19768 17006 19780
rect 20806 19768 20812 19780
rect 17000 19740 20812 19768
rect 17000 19728 17006 19740
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 20901 19771 20959 19777
rect 20901 19737 20913 19771
rect 20947 19737 20959 19771
rect 20901 19731 20959 19737
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 11256 19672 11989 19700
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 11977 19663 12035 19669
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 13906 19700 13912 19712
rect 12124 19672 13912 19700
rect 12124 19660 12130 19672
rect 13906 19660 13912 19672
rect 13964 19660 13970 19712
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 15436 19672 16129 19700
rect 15436 19660 15442 19672
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 16117 19663 16175 19669
rect 20254 19660 20260 19712
rect 20312 19700 20318 19712
rect 20916 19700 20944 19731
rect 20312 19672 20944 19700
rect 23216 19700 23244 19808
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25866 19836 25872 19848
rect 25179 19808 25872 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 25866 19796 25872 19808
rect 25924 19796 25930 19848
rect 26234 19796 26240 19848
rect 26292 19836 26298 19848
rect 26605 19839 26663 19845
rect 26605 19836 26617 19839
rect 26292 19808 26617 19836
rect 26292 19796 26298 19808
rect 26605 19805 26617 19808
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 26881 19839 26939 19845
rect 26881 19805 26893 19839
rect 26927 19836 26939 19839
rect 27525 19839 27583 19845
rect 27525 19836 27537 19839
rect 26927 19808 27537 19836
rect 26927 19805 26939 19808
rect 26881 19799 26939 19805
rect 27525 19805 27537 19808
rect 27571 19836 27583 19839
rect 28169 19839 28227 19845
rect 28169 19836 28181 19839
rect 27571 19808 28181 19836
rect 27571 19805 27583 19808
rect 27525 19799 27583 19805
rect 28169 19805 28181 19808
rect 28215 19805 28227 19839
rect 28810 19836 28816 19848
rect 28771 19808 28816 19836
rect 28169 19799 28227 19805
rect 23382 19768 23388 19780
rect 23343 19740 23388 19768
rect 23382 19728 23388 19740
rect 23440 19728 23446 19780
rect 23474 19728 23480 19780
rect 23532 19768 23538 19780
rect 23532 19740 23577 19768
rect 23532 19728 23538 19740
rect 25406 19728 25412 19780
rect 25464 19768 25470 19780
rect 26896 19768 26924 19799
rect 25464 19740 26924 19768
rect 28184 19768 28212 19799
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 30742 19796 30748 19848
rect 30800 19836 30806 19848
rect 31294 19836 31300 19848
rect 30800 19808 31300 19836
rect 30800 19796 30806 19808
rect 31294 19796 31300 19808
rect 31352 19796 31358 19848
rect 31478 19796 31484 19848
rect 31536 19836 31542 19848
rect 31941 19839 31999 19845
rect 31941 19836 31953 19839
rect 31536 19808 31953 19836
rect 31536 19796 31542 19808
rect 31941 19805 31953 19808
rect 31987 19805 31999 19839
rect 32609 19815 32621 19849
rect 32655 19846 32667 19849
rect 32784 19846 32812 19876
rect 36262 19864 36268 19876
rect 36320 19864 36326 19916
rect 32655 19818 32812 19846
rect 32655 19815 32667 19818
rect 32609 19809 32667 19815
rect 31941 19799 31999 19805
rect 33410 19796 33416 19848
rect 33468 19836 33474 19848
rect 33689 19839 33747 19845
rect 33689 19836 33701 19839
rect 33468 19808 33701 19836
rect 33468 19796 33474 19808
rect 33689 19805 33701 19808
rect 33735 19805 33747 19839
rect 36078 19836 36084 19848
rect 36039 19808 36084 19836
rect 33689 19799 33747 19805
rect 36078 19796 36084 19808
rect 36136 19796 36142 19848
rect 36538 19796 36544 19848
rect 36596 19836 36602 19848
rect 36725 19839 36783 19845
rect 36725 19836 36737 19839
rect 36596 19808 36737 19836
rect 36596 19796 36602 19808
rect 36725 19805 36737 19808
rect 36771 19805 36783 19839
rect 36725 19799 36783 19805
rect 37182 19796 37188 19848
rect 37240 19836 37246 19848
rect 37369 19839 37427 19845
rect 37369 19836 37381 19839
rect 37240 19808 37381 19836
rect 37240 19796 37246 19808
rect 37369 19805 37381 19808
rect 37415 19805 37427 19839
rect 37369 19799 37427 19805
rect 37458 19796 37464 19848
rect 37516 19836 37522 19848
rect 38197 19839 38255 19845
rect 38197 19836 38209 19839
rect 37516 19808 38209 19836
rect 37516 19796 37522 19808
rect 38197 19805 38209 19808
rect 38243 19805 38255 19839
rect 38197 19799 38255 19805
rect 28994 19768 29000 19780
rect 28184 19740 29000 19768
rect 25464 19728 25470 19740
rect 28994 19728 29000 19740
rect 29052 19728 29058 19780
rect 29914 19768 29920 19780
rect 29875 19740 29920 19768
rect 29914 19728 29920 19740
rect 29972 19728 29978 19780
rect 32674 19768 32680 19780
rect 32635 19740 32680 19768
rect 32674 19728 32680 19740
rect 32732 19728 32738 19780
rect 34977 19771 35035 19777
rect 34977 19768 34989 19771
rect 34900 19740 34989 19768
rect 34900 19712 34928 19740
rect 34977 19737 34989 19740
rect 35023 19737 35035 19771
rect 34977 19731 35035 19737
rect 35066 19728 35072 19780
rect 35124 19768 35130 19780
rect 35124 19740 35169 19768
rect 35124 19728 35130 19740
rect 35434 19728 35440 19780
rect 35492 19768 35498 19780
rect 35621 19771 35679 19777
rect 35621 19768 35633 19771
rect 35492 19740 35633 19768
rect 35492 19728 35498 19740
rect 35621 19737 35633 19740
rect 35667 19737 35679 19771
rect 35621 19731 35679 19737
rect 24854 19700 24860 19712
rect 23216 19672 24860 19700
rect 20312 19660 20318 19672
rect 24854 19660 24860 19672
rect 24912 19660 24918 19712
rect 28626 19660 28632 19712
rect 28684 19700 28690 19712
rect 33226 19700 33232 19712
rect 28684 19672 33232 19700
rect 28684 19660 28690 19672
rect 33226 19660 33232 19672
rect 33284 19660 33290 19712
rect 33870 19660 33876 19712
rect 33928 19700 33934 19712
rect 34238 19700 34244 19712
rect 33928 19672 34244 19700
rect 33928 19660 33934 19672
rect 34238 19660 34244 19672
rect 34296 19660 34302 19712
rect 34882 19660 34888 19712
rect 34940 19660 34946 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 1596 19428 1624 19459
rect 6822 19456 6828 19508
rect 6880 19496 6886 19508
rect 7469 19499 7527 19505
rect 7469 19496 7481 19499
rect 6880 19468 7481 19496
rect 6880 19456 6886 19468
rect 7469 19465 7481 19468
rect 7515 19465 7527 19499
rect 7469 19459 7527 19465
rect 7650 19456 7656 19508
rect 7708 19456 7714 19508
rect 12161 19499 12219 19505
rect 10152 19468 11100 19496
rect 7668 19428 7696 19456
rect 8754 19428 8760 19440
rect 1596 19400 7696 19428
rect 8715 19400 8760 19428
rect 8754 19388 8760 19400
rect 8812 19388 8818 19440
rect 10152 19437 10180 19468
rect 10137 19431 10195 19437
rect 10137 19397 10149 19431
rect 10183 19397 10195 19431
rect 10137 19391 10195 19397
rect 10229 19431 10287 19437
rect 10229 19397 10241 19431
rect 10275 19428 10287 19431
rect 10962 19428 10968 19440
rect 10275 19400 10968 19428
rect 10275 19397 10287 19400
rect 10229 19391 10287 19397
rect 10962 19388 10968 19400
rect 11020 19388 11026 19440
rect 1762 19360 1768 19372
rect 1723 19332 1768 19360
rect 1762 19320 1768 19332
rect 1820 19320 1826 19372
rect 7653 19363 7711 19369
rect 7653 19329 7665 19363
rect 7699 19360 7711 19363
rect 7742 19360 7748 19372
rect 7699 19332 7748 19360
rect 7699 19329 7711 19332
rect 7653 19323 7711 19329
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 8110 19320 8116 19372
rect 8168 19360 8174 19372
rect 8168 19332 8524 19360
rect 8168 19320 8174 19332
rect 8496 19292 8524 19332
rect 8665 19295 8723 19301
rect 8665 19292 8677 19295
rect 8496 19264 8677 19292
rect 8665 19261 8677 19264
rect 8711 19261 8723 19295
rect 9122 19292 9128 19304
rect 9083 19264 9128 19292
rect 8665 19255 8723 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 11072 19156 11100 19468
rect 12161 19465 12173 19499
rect 12207 19496 12219 19499
rect 13078 19496 13084 19508
rect 12207 19468 13084 19496
rect 12207 19465 12219 19468
rect 12161 19459 12219 19465
rect 13078 19456 13084 19468
rect 13136 19496 13142 19508
rect 13446 19496 13452 19508
rect 13136 19468 13452 19496
rect 13136 19456 13142 19468
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 14182 19496 14188 19508
rect 14143 19468 14188 19496
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 16945 19499 17003 19505
rect 16945 19465 16957 19499
rect 16991 19496 17003 19499
rect 17494 19496 17500 19508
rect 16991 19468 17500 19496
rect 16991 19465 17003 19468
rect 16945 19459 17003 19465
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 17681 19499 17739 19505
rect 17681 19465 17693 19499
rect 17727 19496 17739 19499
rect 17770 19496 17776 19508
rect 17727 19468 17776 19496
rect 17727 19465 17739 19468
rect 17681 19459 17739 19465
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 18969 19499 19027 19505
rect 18969 19465 18981 19499
rect 19015 19496 19027 19499
rect 19058 19496 19064 19508
rect 19015 19468 19064 19496
rect 19015 19465 19027 19468
rect 18969 19459 19027 19465
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 20254 19496 20260 19508
rect 20215 19468 20260 19496
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 20898 19496 20904 19508
rect 20859 19468 20904 19496
rect 20898 19456 20904 19468
rect 20956 19456 20962 19508
rect 24578 19496 24584 19508
rect 24539 19468 24584 19496
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 24946 19456 24952 19508
rect 25004 19496 25010 19508
rect 25501 19499 25559 19505
rect 25501 19496 25513 19499
rect 25004 19468 25513 19496
rect 25004 19456 25010 19468
rect 25501 19465 25513 19468
rect 25547 19465 25559 19499
rect 25501 19459 25559 19465
rect 25958 19456 25964 19508
rect 26016 19496 26022 19508
rect 26145 19499 26203 19505
rect 26145 19496 26157 19499
rect 26016 19468 26157 19496
rect 26016 19456 26022 19468
rect 26145 19465 26157 19468
rect 26191 19465 26203 19499
rect 27893 19499 27951 19505
rect 27893 19496 27905 19499
rect 26145 19459 26203 19465
rect 26436 19468 27905 19496
rect 11146 19388 11152 19440
rect 11204 19428 11210 19440
rect 12897 19431 12955 19437
rect 12897 19428 12909 19431
rect 11204 19400 12909 19428
rect 11204 19388 11210 19400
rect 12897 19397 12909 19400
rect 12943 19397 12955 19431
rect 12897 19391 12955 19397
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 13538 19428 13544 19440
rect 13228 19400 13544 19428
rect 13228 19388 13234 19400
rect 13538 19388 13544 19400
rect 13596 19428 13602 19440
rect 15378 19428 15384 19440
rect 13596 19400 15148 19428
rect 15339 19400 15384 19428
rect 13596 19388 13602 19400
rect 12066 19360 12072 19372
rect 12027 19332 12072 19360
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 14090 19360 14096 19372
rect 14051 19332 14096 19360
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 11149 19295 11207 19301
rect 11149 19261 11161 19295
rect 11195 19292 11207 19295
rect 12802 19292 12808 19304
rect 11195 19264 12434 19292
rect 12763 19264 12808 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 12406 19236 12434 19264
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 15120 19292 15148 19400
rect 15378 19388 15384 19400
rect 15436 19388 15442 19440
rect 16298 19428 16304 19440
rect 16211 19400 16304 19428
rect 16298 19388 16304 19400
rect 16356 19428 16362 19440
rect 20714 19428 20720 19440
rect 16356 19400 20720 19428
rect 16356 19388 16362 19400
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 25314 19428 25320 19440
rect 20916 19400 25320 19428
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16816 19332 16865 19360
rect 16816 19320 16822 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 17586 19360 17592 19372
rect 17547 19332 17592 19360
rect 16853 19323 16911 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 17678 19320 17684 19372
rect 17736 19360 17742 19372
rect 18877 19363 18935 19369
rect 18877 19360 18889 19363
rect 17736 19332 18889 19360
rect 17736 19320 17742 19332
rect 18877 19329 18889 19332
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 20165 19363 20223 19369
rect 20165 19360 20177 19363
rect 19484 19332 20177 19360
rect 19484 19320 19490 19332
rect 20165 19329 20177 19332
rect 20211 19360 20223 19363
rect 20530 19360 20536 19372
rect 20211 19332 20536 19360
rect 20211 19329 20223 19332
rect 20165 19323 20223 19329
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20806 19360 20812 19372
rect 20719 19332 20812 19360
rect 20806 19320 20812 19332
rect 20864 19360 20870 19372
rect 20916 19360 20944 19400
rect 25314 19388 25320 19400
rect 25372 19388 25378 19440
rect 26436 19428 26464 19468
rect 27893 19465 27905 19468
rect 27939 19465 27951 19499
rect 27893 19459 27951 19465
rect 28994 19456 29000 19508
rect 29052 19496 29058 19508
rect 30190 19496 30196 19508
rect 29052 19468 30196 19496
rect 29052 19456 29058 19468
rect 30190 19456 30196 19468
rect 30248 19456 30254 19508
rect 30282 19456 30288 19508
rect 30340 19496 30346 19508
rect 32401 19499 32459 19505
rect 32401 19496 32413 19499
rect 30340 19468 32413 19496
rect 30340 19456 30346 19468
rect 32401 19465 32413 19468
rect 32447 19465 32459 19499
rect 33226 19496 33232 19508
rect 33187 19468 33232 19496
rect 32401 19459 32459 19465
rect 33226 19456 33232 19468
rect 33284 19456 33290 19508
rect 34330 19456 34336 19508
rect 34388 19496 34394 19508
rect 34701 19499 34759 19505
rect 34701 19496 34713 19499
rect 34388 19468 34713 19496
rect 34388 19456 34394 19468
rect 34701 19465 34713 19468
rect 34747 19465 34759 19499
rect 34701 19459 34759 19465
rect 34790 19456 34796 19508
rect 34848 19496 34854 19508
rect 35250 19496 35256 19508
rect 34848 19468 35256 19496
rect 34848 19456 34854 19468
rect 35250 19456 35256 19468
rect 35308 19456 35314 19508
rect 35986 19456 35992 19508
rect 36044 19496 36050 19508
rect 36173 19499 36231 19505
rect 36173 19496 36185 19499
rect 36044 19468 36185 19496
rect 36044 19456 36050 19468
rect 36173 19465 36185 19468
rect 36219 19465 36231 19499
rect 36814 19496 36820 19508
rect 36775 19468 36820 19496
rect 36173 19459 36231 19465
rect 36814 19456 36820 19468
rect 36872 19456 36878 19508
rect 25516 19400 26464 19428
rect 20864 19332 20944 19360
rect 20864 19320 20870 19332
rect 21634 19320 21640 19372
rect 21692 19360 21698 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21692 19332 22017 19360
rect 21692 19320 21698 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22005 19323 22063 19329
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 23569 19363 23627 19369
rect 23569 19360 23581 19363
rect 22704 19332 23581 19360
rect 22704 19320 22710 19332
rect 23569 19329 23581 19332
rect 23615 19360 23627 19363
rect 24118 19360 24124 19372
rect 23615 19332 24124 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24489 19363 24547 19369
rect 24489 19329 24501 19363
rect 24535 19360 24547 19363
rect 24535 19332 24716 19360
rect 24535 19329 24547 19332
rect 24489 19323 24547 19329
rect 15289 19295 15347 19301
rect 15289 19292 15301 19295
rect 15120 19264 15301 19292
rect 15289 19261 15301 19264
rect 15335 19261 15347 19295
rect 23014 19292 23020 19304
rect 15289 19255 15347 19261
rect 16500 19264 23020 19292
rect 12406 19196 12440 19236
rect 12434 19184 12440 19196
rect 12492 19224 12498 19236
rect 13357 19227 13415 19233
rect 12492 19196 13308 19224
rect 12492 19184 12498 19196
rect 12618 19156 12624 19168
rect 11072 19128 12624 19156
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 13280 19156 13308 19196
rect 13357 19193 13369 19227
rect 13403 19224 13415 19227
rect 13998 19224 14004 19236
rect 13403 19196 14004 19224
rect 13403 19193 13415 19196
rect 13357 19187 13415 19193
rect 13998 19184 14004 19196
rect 14056 19224 14062 19236
rect 16500 19224 16528 19264
rect 23014 19252 23020 19264
rect 23072 19252 23078 19304
rect 23845 19295 23903 19301
rect 23845 19261 23857 19295
rect 23891 19292 23903 19295
rect 23934 19292 23940 19304
rect 23891 19264 23940 19292
rect 23891 19261 23903 19264
rect 23845 19255 23903 19261
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 24688 19292 24716 19332
rect 24762 19320 24768 19372
rect 24820 19360 24826 19372
rect 25406 19360 25412 19372
rect 24820 19332 25268 19360
rect 25367 19332 25412 19360
rect 24820 19320 24826 19332
rect 24854 19292 24860 19304
rect 24688 19264 24860 19292
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 25240 19292 25268 19332
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 25516 19292 25544 19400
rect 26970 19388 26976 19440
rect 27028 19428 27034 19440
rect 27028 19400 28580 19428
rect 27028 19388 27034 19400
rect 26053 19363 26111 19369
rect 26053 19329 26065 19363
rect 26099 19329 26111 19363
rect 26053 19323 26111 19329
rect 25240 19264 25544 19292
rect 26068 19292 26096 19323
rect 26234 19320 26240 19372
rect 26292 19360 26298 19372
rect 26694 19360 26700 19372
rect 26292 19332 26700 19360
rect 26292 19320 26298 19332
rect 26694 19320 26700 19332
rect 26752 19360 26758 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26752 19332 27169 19360
rect 26752 19320 26758 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27246 19320 27252 19372
rect 27304 19360 27310 19372
rect 27304 19332 27349 19360
rect 27304 19320 27310 19332
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 28552 19369 28580 19400
rect 29270 19388 29276 19440
rect 29328 19428 29334 19440
rect 29328 19400 30880 19428
rect 29328 19388 29334 19400
rect 30852 19369 30880 19400
rect 31570 19388 31576 19440
rect 31628 19428 31634 19440
rect 33873 19431 33931 19437
rect 33873 19428 33885 19431
rect 31628 19400 33885 19428
rect 31628 19388 31634 19400
rect 33873 19397 33885 19400
rect 33919 19397 33931 19431
rect 33873 19391 33931 19397
rect 34238 19388 34244 19440
rect 34296 19428 34302 19440
rect 35345 19431 35403 19437
rect 35345 19428 35357 19431
rect 34296 19400 35357 19428
rect 34296 19388 34302 19400
rect 35345 19397 35357 19400
rect 35391 19397 35403 19431
rect 35345 19391 35403 19397
rect 35526 19388 35532 19440
rect 35584 19428 35590 19440
rect 35584 19400 38056 19428
rect 35584 19388 35590 19400
rect 27801 19363 27859 19369
rect 27801 19360 27813 19363
rect 27488 19332 27813 19360
rect 27488 19320 27494 19332
rect 27801 19329 27813 19332
rect 27847 19329 27859 19363
rect 27801 19323 27859 19329
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19329 28595 19363
rect 28537 19323 28595 19329
rect 30837 19363 30895 19369
rect 30837 19329 30849 19363
rect 30883 19329 30895 19363
rect 30837 19323 30895 19329
rect 31110 19320 31116 19372
rect 31168 19360 31174 19372
rect 31938 19360 31944 19372
rect 31168 19332 31944 19360
rect 31168 19320 31174 19332
rect 31938 19320 31944 19332
rect 31996 19320 32002 19372
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19360 32367 19363
rect 33137 19363 33195 19369
rect 33137 19360 33149 19363
rect 32355 19332 33149 19360
rect 32355 19329 32367 19332
rect 32309 19323 32367 19329
rect 33137 19329 33149 19332
rect 33183 19329 33195 19363
rect 33137 19323 33195 19329
rect 33781 19363 33839 19369
rect 33781 19329 33793 19363
rect 33827 19360 33839 19363
rect 34146 19360 34152 19372
rect 33827 19332 34152 19360
rect 33827 19329 33839 19332
rect 33781 19323 33839 19329
rect 28721 19295 28779 19301
rect 26068 19264 28212 19292
rect 22830 19224 22836 19236
rect 14056 19196 16528 19224
rect 16592 19196 22836 19224
rect 14056 19184 14062 19196
rect 16592 19156 16620 19196
rect 22830 19184 22836 19196
rect 22888 19184 22894 19236
rect 24872 19224 24900 19252
rect 25958 19224 25964 19236
rect 24872 19196 25964 19224
rect 25958 19184 25964 19196
rect 26016 19184 26022 19236
rect 13280 19128 16620 19156
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22152 19128 22197 19156
rect 22152 19116 22158 19128
rect 24578 19116 24584 19168
rect 24636 19156 24642 19168
rect 26068 19156 26096 19264
rect 28184 19236 28212 19264
rect 28721 19261 28733 19295
rect 28767 19292 28779 19295
rect 28902 19292 28908 19304
rect 28767 19264 28908 19292
rect 28767 19261 28779 19264
rect 28721 19255 28779 19261
rect 28902 19252 28908 19264
rect 28960 19252 28966 19304
rect 28994 19252 29000 19304
rect 29052 19292 29058 19304
rect 29052 19264 29097 19292
rect 29052 19252 29058 19264
rect 30558 19252 30564 19304
rect 30616 19292 30622 19304
rect 32324 19292 32352 19323
rect 30616 19264 32352 19292
rect 33152 19292 33180 19323
rect 34146 19320 34152 19332
rect 34204 19320 34210 19372
rect 34422 19320 34428 19372
rect 34480 19360 34486 19372
rect 34609 19363 34667 19369
rect 34609 19360 34621 19363
rect 34480 19332 34621 19360
rect 34480 19320 34486 19332
rect 34609 19329 34621 19332
rect 34655 19329 34667 19363
rect 34609 19323 34667 19329
rect 35253 19363 35311 19369
rect 35253 19329 35265 19363
rect 35299 19360 35311 19363
rect 35986 19360 35992 19372
rect 35299 19332 35992 19360
rect 35299 19329 35311 19332
rect 35253 19323 35311 19329
rect 35986 19320 35992 19332
rect 36044 19320 36050 19372
rect 36081 19363 36139 19369
rect 36081 19329 36093 19363
rect 36127 19360 36139 19363
rect 36170 19360 36176 19372
rect 36127 19332 36176 19360
rect 36127 19329 36139 19332
rect 36081 19323 36139 19329
rect 36170 19320 36176 19332
rect 36228 19360 36234 19372
rect 36725 19363 36783 19369
rect 36725 19360 36737 19363
rect 36228 19332 36737 19360
rect 36228 19320 36234 19332
rect 36725 19329 36737 19332
rect 36771 19360 36783 19363
rect 37182 19360 37188 19372
rect 36771 19332 37188 19360
rect 36771 19329 36783 19332
rect 36725 19323 36783 19329
rect 37182 19320 37188 19332
rect 37240 19320 37246 19372
rect 38028 19369 38056 19400
rect 38013 19363 38071 19369
rect 38013 19329 38025 19363
rect 38059 19329 38071 19363
rect 38013 19323 38071 19329
rect 36354 19292 36360 19304
rect 33152 19264 36360 19292
rect 30616 19252 30622 19264
rect 36354 19252 36360 19264
rect 36412 19252 36418 19304
rect 28166 19184 28172 19236
rect 28224 19224 28230 19236
rect 33226 19224 33232 19236
rect 28224 19196 33232 19224
rect 28224 19184 28230 19196
rect 33226 19184 33232 19196
rect 33284 19184 33290 19236
rect 24636 19128 26096 19156
rect 24636 19116 24642 19128
rect 26326 19116 26332 19168
rect 26384 19156 26390 19168
rect 28994 19156 29000 19168
rect 26384 19128 29000 19156
rect 26384 19116 26390 19128
rect 28994 19116 29000 19128
rect 29052 19116 29058 19168
rect 30929 19159 30987 19165
rect 30929 19125 30941 19159
rect 30975 19156 30987 19159
rect 31294 19156 31300 19168
rect 30975 19128 31300 19156
rect 30975 19125 30987 19128
rect 30929 19119 30987 19125
rect 31294 19116 31300 19128
rect 31352 19116 31358 19168
rect 38194 19156 38200 19168
rect 38155 19128 38200 19156
rect 38194 19116 38200 19128
rect 38252 19116 38258 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 15562 18952 15568 18964
rect 15523 18924 15568 18952
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 18325 18955 18383 18961
rect 18325 18921 18337 18955
rect 18371 18952 18383 18955
rect 18506 18952 18512 18964
rect 18371 18924 18512 18952
rect 18371 18921 18383 18924
rect 18325 18915 18383 18921
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 18616 18924 23520 18952
rect 10965 18887 11023 18893
rect 10965 18853 10977 18887
rect 11011 18884 11023 18887
rect 12894 18884 12900 18896
rect 11011 18856 12900 18884
rect 11011 18853 11023 18856
rect 10965 18847 11023 18853
rect 12894 18844 12900 18856
rect 12952 18884 12958 18896
rect 13722 18884 13728 18896
rect 12952 18856 13728 18884
rect 12952 18844 12958 18856
rect 13722 18844 13728 18856
rect 13780 18844 13786 18896
rect 16942 18844 16948 18896
rect 17000 18844 17006 18896
rect 17862 18844 17868 18896
rect 17920 18884 17926 18896
rect 18616 18884 18644 18924
rect 17920 18856 18644 18884
rect 17920 18844 17926 18856
rect 20898 18844 20904 18896
rect 20956 18884 20962 18896
rect 23382 18884 23388 18896
rect 20956 18856 23388 18884
rect 20956 18844 20962 18856
rect 23382 18844 23388 18856
rect 23440 18844 23446 18896
rect 23492 18884 23520 18924
rect 23566 18912 23572 18964
rect 23624 18952 23630 18964
rect 23661 18955 23719 18961
rect 23661 18952 23673 18955
rect 23624 18924 23673 18952
rect 23624 18912 23630 18924
rect 23661 18921 23673 18924
rect 23707 18921 23719 18955
rect 23661 18915 23719 18921
rect 24210 18912 24216 18964
rect 24268 18952 24274 18964
rect 24762 18952 24768 18964
rect 24268 18924 24768 18952
rect 24268 18912 24274 18924
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 26326 18952 26332 18964
rect 26287 18924 26332 18952
rect 26326 18912 26332 18924
rect 26384 18912 26390 18964
rect 27798 18912 27804 18964
rect 27856 18952 27862 18964
rect 28810 18952 28816 18964
rect 27856 18924 28816 18952
rect 27856 18912 27862 18924
rect 28810 18912 28816 18924
rect 28868 18912 28874 18964
rect 29546 18912 29552 18964
rect 29604 18952 29610 18964
rect 30469 18955 30527 18961
rect 30469 18952 30481 18955
rect 29604 18924 30481 18952
rect 29604 18912 29610 18924
rect 30469 18921 30481 18924
rect 30515 18921 30527 18955
rect 30469 18915 30527 18921
rect 31573 18955 31631 18961
rect 31573 18921 31585 18955
rect 31619 18952 31631 18955
rect 32306 18952 32312 18964
rect 31619 18924 32312 18952
rect 31619 18921 31631 18924
rect 31573 18915 31631 18921
rect 32306 18912 32312 18924
rect 32364 18912 32370 18964
rect 33502 18952 33508 18964
rect 32784 18924 33508 18952
rect 23492 18856 31340 18884
rect 9582 18816 9588 18828
rect 9543 18788 9588 18816
rect 9582 18776 9588 18788
rect 9640 18776 9646 18828
rect 10042 18776 10048 18828
rect 10100 18816 10106 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 10100 18788 10425 18816
rect 10100 18776 10106 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 10413 18779 10471 18785
rect 11974 18776 11980 18828
rect 12032 18816 12038 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 12032 18788 12173 18816
rect 12032 18776 12038 18788
rect 12161 18785 12173 18788
rect 12207 18816 12219 18819
rect 16960 18816 16988 18844
rect 12207 18788 14320 18816
rect 12207 18785 12219 18788
rect 12161 18779 12219 18785
rect 7742 18708 7748 18760
rect 7800 18748 7806 18760
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 7800 18720 8217 18748
rect 7800 18708 7806 18720
rect 8205 18717 8217 18720
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 10505 18683 10563 18689
rect 10505 18649 10517 18683
rect 10551 18680 10563 18683
rect 10594 18680 10600 18692
rect 10551 18652 10600 18680
rect 10551 18649 10563 18652
rect 10505 18643 10563 18649
rect 10594 18640 10600 18652
rect 10652 18640 10658 18692
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 13170 18680 13176 18692
rect 12308 18652 12353 18680
rect 13131 18652 13176 18680
rect 12308 18640 12314 18652
rect 13170 18640 13176 18652
rect 13228 18640 13234 18692
rect 8297 18615 8355 18621
rect 8297 18581 8309 18615
rect 8343 18612 8355 18615
rect 9306 18612 9312 18624
rect 8343 18584 9312 18612
rect 8343 18581 8355 18584
rect 8297 18575 8355 18581
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 14292 18612 14320 18788
rect 15488 18788 16988 18816
rect 19429 18819 19487 18825
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 15194 18748 15200 18760
rect 14691 18720 15200 18748
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 15488 18757 15516 18788
rect 19429 18785 19441 18819
rect 19475 18816 19487 18819
rect 19978 18816 19984 18828
rect 19475 18788 19984 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 21266 18816 21272 18828
rect 21227 18788 21272 18816
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 21542 18776 21548 18828
rect 21600 18816 21606 18828
rect 21821 18819 21879 18825
rect 21821 18816 21833 18819
rect 21600 18788 21833 18816
rect 21600 18776 21606 18788
rect 21821 18785 21833 18788
rect 21867 18785 21879 18819
rect 21821 18779 21879 18785
rect 22462 18776 22468 18828
rect 22520 18816 22526 18828
rect 24673 18819 24731 18825
rect 24673 18816 24685 18819
rect 22520 18788 24685 18816
rect 22520 18776 22526 18788
rect 24673 18785 24685 18788
rect 24719 18785 24731 18819
rect 26418 18816 26424 18828
rect 24673 18779 24731 18785
rect 26252 18788 26424 18816
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16942 18748 16948 18760
rect 16163 18720 16948 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17678 18708 17684 18760
rect 17736 18748 17742 18760
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 17736 18720 18245 18748
rect 17736 18708 17742 18720
rect 18233 18717 18245 18720
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 24578 18748 24584 18760
rect 23615 18720 23796 18748
rect 24539 18720 24584 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 14737 18683 14795 18689
rect 14737 18649 14749 18683
rect 14783 18680 14795 18683
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 14783 18652 19625 18680
rect 14783 18649 14795 18652
rect 14737 18643 14795 18649
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 19613 18643 19671 18649
rect 21913 18683 21971 18689
rect 21913 18649 21925 18683
rect 21959 18680 21971 18683
rect 22094 18680 22100 18692
rect 21959 18652 22100 18680
rect 21959 18649 21971 18652
rect 21913 18643 21971 18649
rect 22094 18640 22100 18652
rect 22152 18640 22158 18692
rect 22830 18680 22836 18692
rect 22791 18652 22836 18680
rect 22830 18640 22836 18652
rect 22888 18640 22894 18692
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 14292 18584 16221 18612
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16209 18575 16267 18581
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 23658 18612 23664 18624
rect 17092 18584 23664 18612
rect 17092 18572 17098 18584
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 23768 18612 23796 18720
rect 24578 18708 24584 18720
rect 24636 18708 24642 18760
rect 24762 18708 24768 18760
rect 24820 18748 24826 18760
rect 26252 18757 26280 18788
rect 26418 18776 26424 18788
rect 26476 18816 26482 18828
rect 27430 18816 27436 18828
rect 26476 18788 27436 18816
rect 26476 18776 26482 18788
rect 27430 18776 27436 18788
rect 27488 18776 27494 18828
rect 27982 18816 27988 18828
rect 27943 18788 27988 18816
rect 27982 18776 27988 18788
rect 28040 18776 28046 18828
rect 30558 18816 30564 18828
rect 28460 18788 30564 18816
rect 25225 18751 25283 18757
rect 25225 18748 25237 18751
rect 24820 18720 25237 18748
rect 24820 18708 24826 18720
rect 25225 18717 25237 18720
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 26237 18751 26295 18757
rect 26237 18717 26249 18751
rect 26283 18717 26295 18751
rect 26237 18711 26295 18717
rect 27890 18708 27896 18760
rect 27948 18748 27954 18760
rect 28460 18757 28488 18788
rect 30558 18776 30564 18788
rect 30616 18776 30622 18828
rect 31312 18816 31340 18856
rect 32784 18816 32812 18924
rect 33502 18912 33508 18924
rect 33560 18952 33566 18964
rect 34054 18952 34060 18964
rect 33560 18924 34060 18952
rect 33560 18912 33566 18924
rect 34054 18912 34060 18924
rect 34112 18912 34118 18964
rect 34149 18955 34207 18961
rect 34149 18921 34161 18955
rect 34195 18952 34207 18955
rect 34698 18952 34704 18964
rect 34195 18924 34704 18952
rect 34195 18921 34207 18924
rect 34149 18915 34207 18921
rect 34698 18912 34704 18924
rect 34756 18912 34762 18964
rect 35250 18912 35256 18964
rect 35308 18952 35314 18964
rect 35713 18955 35771 18961
rect 35713 18952 35725 18955
rect 35308 18924 35725 18952
rect 35308 18912 35314 18924
rect 35713 18921 35725 18924
rect 35759 18921 35771 18955
rect 35713 18915 35771 18921
rect 36357 18955 36415 18961
rect 36357 18921 36369 18955
rect 36403 18952 36415 18955
rect 38838 18952 38844 18964
rect 36403 18924 38844 18952
rect 36403 18921 36415 18924
rect 36357 18915 36415 18921
rect 38838 18912 38844 18924
rect 38896 18912 38902 18964
rect 33229 18887 33287 18893
rect 33229 18853 33241 18887
rect 33275 18884 33287 18887
rect 34606 18884 34612 18896
rect 33275 18856 34612 18884
rect 33275 18853 33287 18856
rect 33229 18847 33287 18853
rect 34606 18844 34612 18856
rect 34664 18844 34670 18896
rect 37550 18844 37556 18896
rect 37608 18884 37614 18896
rect 37608 18856 37872 18884
rect 37608 18844 37614 18856
rect 31312 18788 32812 18816
rect 32858 18776 32864 18828
rect 32916 18816 32922 18828
rect 37734 18816 37740 18828
rect 32916 18788 34100 18816
rect 32916 18776 32922 18788
rect 28445 18751 28503 18757
rect 28445 18748 28457 18751
rect 27948 18720 28457 18748
rect 27948 18708 27954 18720
rect 28445 18717 28457 18720
rect 28491 18717 28503 18751
rect 29730 18748 29736 18760
rect 29691 18720 29736 18748
rect 28445 18711 28503 18717
rect 29730 18708 29736 18720
rect 29788 18708 29794 18760
rect 30377 18751 30435 18757
rect 30377 18717 30389 18751
rect 30423 18748 30435 18751
rect 30742 18748 30748 18760
rect 30423 18720 30748 18748
rect 30423 18717 30435 18720
rect 30377 18711 30435 18717
rect 30742 18708 30748 18720
rect 30800 18708 30806 18760
rect 31110 18708 31116 18760
rect 31168 18748 31174 18760
rect 31473 18751 31531 18757
rect 31473 18748 31485 18751
rect 31168 18720 31485 18748
rect 31168 18708 31174 18720
rect 31473 18717 31485 18720
rect 31519 18717 31531 18751
rect 33134 18748 33140 18760
rect 33095 18720 33140 18748
rect 31473 18711 31531 18717
rect 33134 18708 33140 18720
rect 33192 18708 33198 18760
rect 34072 18757 34100 18788
rect 34992 18788 37740 18816
rect 34057 18751 34115 18757
rect 34057 18717 34069 18751
rect 34103 18717 34115 18751
rect 34057 18711 34115 18717
rect 34146 18708 34152 18760
rect 34204 18748 34210 18760
rect 34992 18757 35020 18788
rect 37734 18776 37740 18788
rect 37792 18776 37798 18828
rect 37844 18825 37872 18856
rect 37829 18819 37887 18825
rect 37829 18785 37841 18819
rect 37875 18785 37887 18819
rect 37829 18779 37887 18785
rect 34977 18751 35035 18757
rect 34977 18748 34989 18751
rect 34204 18720 34989 18748
rect 34204 18708 34210 18720
rect 34977 18717 34989 18720
rect 35023 18717 35035 18751
rect 34977 18711 35035 18717
rect 35621 18751 35679 18757
rect 35621 18717 35633 18751
rect 35667 18717 35679 18751
rect 35621 18711 35679 18717
rect 23842 18640 23848 18692
rect 23900 18680 23906 18692
rect 25317 18683 25375 18689
rect 25317 18680 25329 18683
rect 23900 18652 25329 18680
rect 23900 18640 23906 18652
rect 25317 18649 25329 18652
rect 25363 18649 25375 18683
rect 25317 18643 25375 18649
rect 25958 18640 25964 18692
rect 26016 18680 26022 18692
rect 26970 18680 26976 18692
rect 26016 18652 26372 18680
rect 26931 18652 26976 18680
rect 26016 18640 26022 18652
rect 26234 18612 26240 18624
rect 23768 18584 26240 18612
rect 26234 18572 26240 18584
rect 26292 18572 26298 18624
rect 26344 18612 26372 18652
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 27065 18683 27123 18689
rect 27065 18649 27077 18683
rect 27111 18680 27123 18683
rect 27430 18680 27436 18692
rect 27111 18652 27436 18680
rect 27111 18649 27123 18652
rect 27065 18643 27123 18649
rect 27430 18640 27436 18652
rect 27488 18640 27494 18692
rect 28721 18683 28779 18689
rect 28721 18649 28733 18683
rect 28767 18680 28779 18683
rect 32858 18680 32864 18692
rect 28767 18652 32864 18680
rect 28767 18649 28779 18652
rect 28721 18643 28779 18649
rect 28736 18612 28764 18643
rect 32858 18640 32864 18652
rect 32916 18640 32922 18692
rect 33042 18640 33048 18692
rect 33100 18680 33106 18692
rect 35636 18680 35664 18711
rect 35894 18708 35900 18760
rect 35952 18748 35958 18760
rect 36170 18748 36176 18760
rect 35952 18720 36176 18748
rect 35952 18708 35958 18720
rect 36170 18708 36176 18720
rect 36228 18748 36234 18760
rect 36265 18751 36323 18757
rect 36265 18748 36277 18751
rect 36228 18720 36277 18748
rect 36228 18708 36234 18720
rect 36265 18717 36277 18720
rect 36311 18717 36323 18751
rect 36265 18711 36323 18717
rect 37274 18680 37280 18692
rect 33100 18652 35664 18680
rect 37235 18652 37280 18680
rect 33100 18640 33106 18652
rect 37274 18640 37280 18652
rect 37332 18640 37338 18692
rect 37366 18640 37372 18692
rect 37424 18680 37430 18692
rect 37424 18652 37469 18680
rect 37424 18640 37430 18652
rect 26344 18584 28764 18612
rect 29825 18615 29883 18621
rect 29825 18581 29837 18615
rect 29871 18612 29883 18615
rect 30006 18612 30012 18624
rect 29871 18584 30012 18612
rect 29871 18581 29883 18584
rect 29825 18575 29883 18581
rect 30006 18572 30012 18584
rect 30064 18572 30070 18624
rect 32398 18572 32404 18624
rect 32456 18612 32462 18624
rect 35069 18615 35127 18621
rect 35069 18612 35081 18615
rect 32456 18584 35081 18612
rect 32456 18572 32462 18584
rect 35069 18581 35081 18584
rect 35115 18581 35127 18615
rect 37292 18612 37320 18640
rect 37918 18612 37924 18624
rect 37292 18584 37924 18612
rect 35069 18575 35127 18581
rect 37918 18572 37924 18584
rect 37976 18572 37982 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7653 18411 7711 18417
rect 7653 18408 7665 18411
rect 7524 18380 7665 18408
rect 7524 18368 7530 18380
rect 7653 18377 7665 18380
rect 7699 18377 7711 18411
rect 7653 18371 7711 18377
rect 9033 18411 9091 18417
rect 9033 18377 9045 18411
rect 9079 18408 9091 18411
rect 9766 18408 9772 18420
rect 9079 18380 9772 18408
rect 9079 18377 9091 18380
rect 9033 18371 9091 18377
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 10229 18411 10287 18417
rect 10229 18377 10241 18411
rect 10275 18408 10287 18411
rect 11514 18408 11520 18420
rect 10275 18380 11520 18408
rect 10275 18377 10287 18380
rect 10229 18371 10287 18377
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 19242 18408 19248 18420
rect 12360 18380 19248 18408
rect 10502 18340 10508 18352
rect 8588 18312 10508 18340
rect 4614 18232 4620 18284
rect 4672 18272 4678 18284
rect 8588 18281 8616 18312
rect 10502 18300 10508 18312
rect 10560 18300 10566 18352
rect 12360 18349 12388 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 22465 18411 22523 18417
rect 22465 18377 22477 18411
rect 22511 18408 22523 18411
rect 23474 18408 23480 18420
rect 22511 18380 23480 18408
rect 22511 18377 22523 18380
rect 22465 18371 22523 18377
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 24394 18408 24400 18420
rect 24355 18380 24400 18408
rect 24394 18368 24400 18380
rect 24452 18368 24458 18420
rect 26050 18408 26056 18420
rect 26011 18380 26056 18408
rect 26050 18368 26056 18380
rect 26108 18368 26114 18420
rect 27430 18408 27436 18420
rect 27391 18380 27436 18408
rect 27430 18368 27436 18380
rect 27488 18368 27494 18420
rect 28718 18408 28724 18420
rect 28679 18380 28724 18408
rect 28718 18368 28724 18380
rect 28776 18368 28782 18420
rect 28902 18368 28908 18420
rect 28960 18408 28966 18420
rect 29365 18411 29423 18417
rect 29365 18408 29377 18411
rect 28960 18380 29377 18408
rect 28960 18368 28966 18380
rect 29365 18377 29377 18380
rect 29411 18377 29423 18411
rect 29365 18371 29423 18377
rect 32122 18368 32128 18420
rect 32180 18408 32186 18420
rect 33594 18408 33600 18420
rect 32180 18380 33456 18408
rect 33555 18380 33600 18408
rect 32180 18368 32186 18380
rect 12345 18343 12403 18349
rect 12345 18309 12357 18343
rect 12391 18309 12403 18343
rect 13906 18340 13912 18352
rect 13867 18312 13912 18340
rect 12345 18303 12403 18309
rect 13906 18300 13912 18312
rect 13964 18300 13970 18352
rect 21910 18300 21916 18352
rect 21968 18340 21974 18352
rect 23753 18343 23811 18349
rect 23753 18340 23765 18343
rect 21968 18312 23765 18340
rect 21968 18300 21974 18312
rect 23753 18309 23765 18312
rect 23799 18309 23811 18343
rect 23753 18303 23811 18309
rect 24762 18300 24768 18352
rect 24820 18340 24826 18352
rect 24820 18312 26096 18340
rect 24820 18300 24826 18312
rect 7561 18275 7619 18281
rect 7561 18272 7573 18275
rect 4672 18244 7573 18272
rect 4672 18232 4678 18244
rect 7561 18241 7573 18244
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 1578 18204 1584 18216
rect 1539 18176 1584 18204
rect 1578 18164 1584 18176
rect 1636 18164 1642 18216
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 7926 18204 7932 18216
rect 1903 18176 7932 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9232 18204 9260 18235
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 9456 18244 10149 18272
rect 9456 18232 9462 18244
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10778 18272 10784 18284
rect 10739 18244 10784 18272
rect 10137 18235 10195 18241
rect 10778 18232 10784 18244
rect 10836 18232 10842 18284
rect 14550 18272 14556 18284
rect 14511 18244 14556 18272
rect 14550 18232 14556 18244
rect 14608 18232 14614 18284
rect 19426 18272 19432 18284
rect 19387 18244 19432 18272
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 22370 18272 22376 18284
rect 22331 18244 22376 18272
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 23017 18275 23075 18281
rect 23017 18241 23029 18275
rect 23063 18241 23075 18275
rect 23017 18235 23075 18241
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18272 23719 18275
rect 23934 18272 23940 18284
rect 23707 18244 23940 18272
rect 23707 18241 23719 18244
rect 23661 18235 23719 18241
rect 8404 18176 9260 18204
rect 12253 18207 12311 18213
rect 8404 18145 8432 18176
rect 12253 18173 12265 18207
rect 12299 18204 12311 18207
rect 12618 18204 12624 18216
rect 12299 18176 12624 18204
rect 12299 18173 12311 18176
rect 12253 18167 12311 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 13262 18204 13268 18216
rect 13223 18176 13268 18204
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 21634 18164 21640 18216
rect 21692 18204 21698 18216
rect 23032 18204 23060 18235
rect 23934 18232 23940 18244
rect 23992 18272 23998 18284
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 23992 18244 24317 18272
rect 23992 18232 23998 18244
rect 24305 18241 24317 18244
rect 24351 18272 24363 18275
rect 25133 18275 25191 18281
rect 25133 18272 25145 18275
rect 24351 18244 25145 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 25133 18241 25145 18244
rect 25179 18272 25191 18275
rect 25958 18272 25964 18284
rect 25179 18244 25820 18272
rect 25919 18244 25964 18272
rect 25179 18241 25191 18244
rect 25133 18235 25191 18241
rect 21692 18176 23060 18204
rect 21692 18164 21698 18176
rect 23382 18164 23388 18216
rect 23440 18204 23446 18216
rect 25792 18204 25820 18244
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26068 18272 26096 18312
rect 27062 18300 27068 18352
rect 27120 18340 27126 18352
rect 28077 18343 28135 18349
rect 28077 18340 28089 18343
rect 27120 18312 28089 18340
rect 27120 18300 27126 18312
rect 28077 18309 28089 18312
rect 28123 18309 28135 18343
rect 30742 18340 30748 18352
rect 28077 18303 28135 18309
rect 28644 18312 30748 18340
rect 27341 18275 27399 18281
rect 27341 18272 27353 18275
rect 26068 18244 27353 18272
rect 27341 18241 27353 18244
rect 27387 18241 27399 18275
rect 27341 18235 27399 18241
rect 27985 18275 28043 18281
rect 27985 18241 27997 18275
rect 28031 18272 28043 18275
rect 28166 18272 28172 18284
rect 28031 18244 28172 18272
rect 28031 18241 28043 18244
rect 27985 18235 28043 18241
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 28644 18281 28672 18312
rect 30742 18300 30748 18312
rect 30800 18300 30806 18352
rect 31202 18340 31208 18352
rect 31163 18312 31208 18340
rect 31202 18300 31208 18312
rect 31260 18300 31266 18352
rect 31294 18300 31300 18352
rect 31352 18340 31358 18352
rect 32493 18343 32551 18349
rect 32493 18340 32505 18343
rect 31352 18312 32505 18340
rect 31352 18300 31358 18312
rect 32493 18309 32505 18312
rect 32539 18309 32551 18343
rect 33428 18340 33456 18380
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 34606 18368 34612 18420
rect 34664 18408 34670 18420
rect 35434 18408 35440 18420
rect 34664 18380 35440 18408
rect 34664 18368 34670 18380
rect 35434 18368 35440 18380
rect 35492 18368 35498 18420
rect 36817 18411 36875 18417
rect 36817 18377 36829 18411
rect 36863 18408 36875 18411
rect 36998 18408 37004 18420
rect 36863 18380 37004 18408
rect 36863 18377 36875 18380
rect 36817 18371 36875 18377
rect 36998 18368 37004 18380
rect 37056 18368 37062 18420
rect 37826 18368 37832 18420
rect 37884 18408 37890 18420
rect 37921 18411 37979 18417
rect 37921 18408 37933 18411
rect 37884 18380 37933 18408
rect 37884 18368 37890 18380
rect 37921 18377 37933 18380
rect 37967 18377 37979 18411
rect 37921 18371 37979 18377
rect 35069 18343 35127 18349
rect 35069 18340 35081 18343
rect 33428 18312 35081 18340
rect 32493 18303 32551 18309
rect 35069 18309 35081 18312
rect 35115 18309 35127 18343
rect 36538 18340 36544 18352
rect 35069 18303 35127 18309
rect 35728 18312 36544 18340
rect 28629 18275 28687 18281
rect 28629 18241 28641 18275
rect 28675 18241 28687 18275
rect 28629 18235 28687 18241
rect 28644 18204 28672 18235
rect 28810 18232 28816 18284
rect 28868 18272 28874 18284
rect 29273 18275 29331 18281
rect 29273 18272 29285 18275
rect 28868 18244 29285 18272
rect 28868 18232 28874 18244
rect 29273 18241 29285 18244
rect 29319 18272 29331 18275
rect 30466 18272 30472 18284
rect 29319 18244 30472 18272
rect 29319 18241 29331 18244
rect 29273 18235 29331 18241
rect 30466 18232 30472 18244
rect 30524 18232 30530 18284
rect 33134 18232 33140 18284
rect 33192 18272 33198 18284
rect 33505 18275 33563 18281
rect 33505 18272 33517 18275
rect 33192 18244 33517 18272
rect 33192 18232 33198 18244
rect 33505 18241 33517 18244
rect 33551 18272 33563 18275
rect 34146 18272 34152 18284
rect 33551 18244 34152 18272
rect 33551 18241 33563 18244
rect 33505 18235 33563 18241
rect 34146 18232 34152 18244
rect 34204 18232 34210 18284
rect 34425 18275 34483 18281
rect 34425 18241 34437 18275
rect 34471 18272 34483 18275
rect 34606 18272 34612 18284
rect 34471 18244 34612 18272
rect 34471 18241 34483 18244
rect 34425 18235 34483 18241
rect 34606 18232 34612 18244
rect 34664 18232 34670 18284
rect 34977 18275 35035 18281
rect 34977 18241 34989 18275
rect 35023 18272 35035 18275
rect 35728 18272 35756 18312
rect 36538 18300 36544 18312
rect 36596 18300 36602 18352
rect 35023 18244 35756 18272
rect 35805 18275 35863 18281
rect 35023 18241 35035 18244
rect 34977 18235 35035 18241
rect 35805 18241 35817 18275
rect 35851 18241 35863 18275
rect 35805 18235 35863 18241
rect 23440 18176 25452 18204
rect 25792 18176 28672 18204
rect 31113 18207 31171 18213
rect 23440 18164 23446 18176
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18105 8447 18139
rect 25225 18139 25283 18145
rect 25225 18136 25237 18139
rect 8389 18099 8447 18105
rect 22388 18108 25237 18136
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 10873 18071 10931 18077
rect 10873 18068 10885 18071
rect 10468 18040 10885 18068
rect 10468 18028 10474 18040
rect 10873 18037 10885 18040
rect 10919 18037 10931 18071
rect 13998 18068 14004 18080
rect 13959 18040 14004 18068
rect 10873 18031 10931 18037
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 14090 18028 14096 18080
rect 14148 18068 14154 18080
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 14148 18040 14657 18068
rect 14148 18028 14154 18040
rect 14645 18037 14657 18040
rect 14691 18037 14703 18071
rect 14645 18031 14703 18037
rect 19245 18071 19303 18077
rect 19245 18037 19257 18071
rect 19291 18068 19303 18071
rect 19610 18068 19616 18080
rect 19291 18040 19616 18068
rect 19291 18037 19303 18040
rect 19245 18031 19303 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 21450 18028 21456 18080
rect 21508 18068 21514 18080
rect 22388 18068 22416 18108
rect 25225 18105 25237 18108
rect 25271 18105 25283 18139
rect 25225 18099 25283 18105
rect 21508 18040 22416 18068
rect 23109 18071 23167 18077
rect 21508 18028 21514 18040
rect 23109 18037 23121 18071
rect 23155 18068 23167 18071
rect 25314 18068 25320 18080
rect 23155 18040 25320 18068
rect 23155 18037 23167 18040
rect 23109 18031 23167 18037
rect 25314 18028 25320 18040
rect 25372 18028 25378 18080
rect 25424 18068 25452 18176
rect 31113 18173 31125 18207
rect 31159 18173 31171 18207
rect 31386 18204 31392 18216
rect 31347 18176 31392 18204
rect 31113 18167 31171 18173
rect 31128 18136 31156 18167
rect 31386 18164 31392 18176
rect 31444 18164 31450 18216
rect 32401 18207 32459 18213
rect 32401 18204 32413 18207
rect 31588 18176 32413 18204
rect 28368 18108 31156 18136
rect 28368 18068 28396 18108
rect 25424 18040 28396 18068
rect 28442 18028 28448 18080
rect 28500 18068 28506 18080
rect 31588 18068 31616 18176
rect 32401 18173 32413 18176
rect 32447 18173 32459 18207
rect 32401 18167 32459 18173
rect 32858 18164 32864 18216
rect 32916 18204 32922 18216
rect 34992 18204 35020 18235
rect 35820 18204 35848 18235
rect 36354 18232 36360 18284
rect 36412 18272 36418 18284
rect 36725 18275 36783 18281
rect 36725 18272 36737 18275
rect 36412 18244 36737 18272
rect 36412 18232 36418 18244
rect 36725 18241 36737 18244
rect 36771 18272 36783 18275
rect 37182 18272 37188 18284
rect 36771 18244 37188 18272
rect 36771 18241 36783 18244
rect 36725 18235 36783 18241
rect 37182 18232 37188 18244
rect 37240 18232 37246 18284
rect 37826 18272 37832 18284
rect 37787 18244 37832 18272
rect 37826 18232 37832 18244
rect 37884 18232 37890 18284
rect 32916 18176 35020 18204
rect 35084 18176 35848 18204
rect 32916 18164 32922 18176
rect 31662 18096 31668 18148
rect 31720 18136 31726 18148
rect 32953 18139 33011 18145
rect 32953 18136 32965 18139
rect 31720 18108 32965 18136
rect 31720 18096 31726 18108
rect 32953 18105 32965 18108
rect 32999 18136 33011 18139
rect 33042 18136 33048 18148
rect 32999 18108 33048 18136
rect 32999 18105 33011 18108
rect 32953 18099 33011 18105
rect 33042 18096 33048 18108
rect 33100 18096 33106 18148
rect 28500 18040 31616 18068
rect 34425 18071 34483 18077
rect 28500 18028 28506 18040
rect 34425 18037 34437 18071
rect 34471 18068 34483 18071
rect 35084 18068 35112 18176
rect 36446 18164 36452 18216
rect 36504 18204 36510 18216
rect 38470 18204 38476 18216
rect 36504 18176 38476 18204
rect 36504 18164 36510 18176
rect 38470 18164 38476 18176
rect 38528 18164 38534 18216
rect 35621 18139 35679 18145
rect 35621 18105 35633 18139
rect 35667 18136 35679 18139
rect 38010 18136 38016 18148
rect 35667 18108 38016 18136
rect 35667 18105 35679 18108
rect 35621 18099 35679 18105
rect 38010 18096 38016 18108
rect 38068 18096 38074 18148
rect 34471 18040 35112 18068
rect 34471 18037 34483 18040
rect 34425 18031 34483 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 11514 17824 11520 17876
rect 11572 17864 11578 17876
rect 12342 17864 12348 17876
rect 11572 17836 12348 17864
rect 11572 17824 11578 17836
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 20070 17824 20076 17876
rect 20128 17864 20134 17876
rect 24578 17864 24584 17876
rect 20128 17836 24584 17864
rect 20128 17824 20134 17836
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 25222 17824 25228 17876
rect 25280 17864 25286 17876
rect 25777 17867 25835 17873
rect 25777 17864 25789 17867
rect 25280 17836 25789 17864
rect 25280 17824 25286 17836
rect 25777 17833 25789 17836
rect 25823 17833 25835 17867
rect 25777 17827 25835 17833
rect 27985 17867 28043 17873
rect 27985 17833 27997 17867
rect 28031 17864 28043 17867
rect 28074 17864 28080 17876
rect 28031 17836 28080 17864
rect 28031 17833 28043 17836
rect 27985 17827 28043 17833
rect 28074 17824 28080 17836
rect 28132 17824 28138 17876
rect 28626 17864 28632 17876
rect 28587 17836 28632 17864
rect 28626 17824 28632 17836
rect 28684 17824 28690 17876
rect 30466 17824 30472 17876
rect 30524 17864 30530 17876
rect 34146 17864 34152 17876
rect 30524 17836 34152 17864
rect 30524 17824 30530 17836
rect 34146 17824 34152 17836
rect 34204 17824 34210 17876
rect 37921 17867 37979 17873
rect 37921 17833 37933 17867
rect 37967 17864 37979 17867
rect 38562 17864 38568 17876
rect 37967 17836 38568 17864
rect 37967 17833 37979 17836
rect 37921 17827 37979 17833
rect 38562 17824 38568 17836
rect 38620 17824 38626 17876
rect 21358 17756 21364 17808
rect 21416 17796 21422 17808
rect 30558 17796 30564 17808
rect 21416 17768 30564 17796
rect 21416 17756 21422 17768
rect 30558 17756 30564 17768
rect 30616 17756 30622 17808
rect 31018 17756 31024 17808
rect 31076 17796 31082 17808
rect 37277 17799 37335 17805
rect 31076 17768 36032 17796
rect 31076 17756 31082 17768
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 7926 17728 7932 17740
rect 7340 17700 7932 17728
rect 7340 17688 7346 17700
rect 7926 17688 7932 17700
rect 7984 17728 7990 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 7984 17700 9689 17728
rect 7984 17688 7990 17700
rect 9677 17697 9689 17700
rect 9723 17697 9735 17731
rect 9677 17691 9735 17697
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 11057 17731 11115 17737
rect 11057 17728 11069 17731
rect 9916 17700 11069 17728
rect 9916 17688 9922 17700
rect 11057 17697 11069 17700
rect 11103 17697 11115 17731
rect 13078 17728 13084 17740
rect 13039 17700 13084 17728
rect 11057 17691 11115 17697
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 20622 17688 20628 17740
rect 20680 17728 20686 17740
rect 23753 17731 23811 17737
rect 23753 17728 23765 17731
rect 20680 17700 23765 17728
rect 20680 17688 20686 17700
rect 23753 17697 23765 17700
rect 23799 17697 23811 17731
rect 30374 17728 30380 17740
rect 23753 17691 23811 17697
rect 26252 17700 27476 17728
rect 30335 17700 30380 17728
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 14274 17660 14280 17672
rect 8343 17632 9076 17660
rect 14235 17632 14280 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 8846 17524 8852 17536
rect 8435 17496 8852 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 8846 17484 8852 17496
rect 8904 17484 8910 17536
rect 9048 17524 9076 17632
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 15712 17632 18705 17660
rect 15712 17620 15718 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 19610 17660 19616 17672
rect 19571 17632 19616 17660
rect 18693 17623 18751 17629
rect 19610 17620 19616 17632
rect 19668 17620 19674 17672
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 23014 17660 23020 17672
rect 22612 17632 23020 17660
rect 22612 17620 22618 17632
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17660 23719 17663
rect 23934 17660 23940 17672
rect 23707 17632 23940 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 23934 17620 23940 17632
rect 23992 17620 23998 17672
rect 25130 17620 25136 17672
rect 25188 17660 25194 17672
rect 25682 17660 25688 17672
rect 25188 17632 25688 17660
rect 25188 17620 25194 17632
rect 25682 17620 25688 17632
rect 25740 17620 25746 17672
rect 9214 17592 9220 17604
rect 9175 17564 9220 17592
rect 9214 17552 9220 17564
rect 9272 17552 9278 17604
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 9364 17564 9409 17592
rect 9364 17552 9370 17564
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 12066 17592 12072 17604
rect 11204 17564 11249 17592
rect 12027 17564 12072 17592
rect 11204 17552 11210 17564
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 13173 17595 13231 17601
rect 13173 17561 13185 17595
rect 13219 17561 13231 17595
rect 13173 17555 13231 17561
rect 13725 17595 13783 17601
rect 13725 17561 13737 17595
rect 13771 17592 13783 17595
rect 15102 17592 15108 17604
rect 13771 17564 15108 17592
rect 13771 17561 13783 17564
rect 13725 17555 13783 17561
rect 10778 17524 10784 17536
rect 9048 17496 10784 17524
rect 10778 17484 10784 17496
rect 10836 17484 10842 17536
rect 13188 17524 13216 17555
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 16666 17552 16672 17604
rect 16724 17592 16730 17604
rect 26252 17592 26280 17700
rect 26421 17595 26479 17601
rect 26421 17592 26433 17595
rect 16724 17564 26280 17592
rect 26344 17564 26433 17592
rect 16724 17552 16730 17564
rect 26344 17536 26372 17564
rect 26421 17561 26433 17564
rect 26467 17561 26479 17595
rect 26421 17555 26479 17561
rect 26513 17595 26571 17601
rect 26513 17561 26525 17595
rect 26559 17592 26571 17595
rect 27246 17592 27252 17604
rect 26559 17564 27252 17592
rect 26559 17561 26571 17564
rect 26513 17555 26571 17561
rect 27246 17552 27252 17564
rect 27304 17552 27310 17604
rect 27448 17601 27476 17700
rect 30374 17688 30380 17700
rect 30432 17688 30438 17740
rect 31386 17688 31392 17740
rect 31444 17728 31450 17740
rect 31662 17728 31668 17740
rect 31444 17700 31668 17728
rect 31444 17688 31450 17700
rect 31662 17688 31668 17700
rect 31720 17688 31726 17740
rect 35342 17728 35348 17740
rect 32876 17700 35348 17728
rect 27890 17660 27896 17672
rect 27851 17632 27896 17660
rect 27890 17620 27896 17632
rect 27948 17620 27954 17672
rect 28166 17620 28172 17672
rect 28224 17660 28230 17672
rect 32876 17669 32904 17700
rect 35342 17688 35348 17700
rect 35400 17688 35406 17740
rect 35894 17728 35900 17740
rect 35855 17700 35900 17728
rect 35894 17688 35900 17700
rect 35952 17688 35958 17740
rect 36004 17728 36032 17768
rect 37277 17765 37289 17799
rect 37323 17796 37335 17799
rect 39574 17796 39580 17808
rect 37323 17768 39580 17796
rect 37323 17765 37335 17768
rect 37277 17759 37335 17765
rect 39574 17756 39580 17768
rect 39632 17756 39638 17808
rect 37734 17728 37740 17740
rect 36004 17700 37740 17728
rect 37734 17688 37740 17700
rect 37792 17688 37798 17740
rect 28537 17663 28595 17669
rect 28537 17660 28549 17663
rect 28224 17632 28549 17660
rect 28224 17620 28230 17632
rect 28537 17629 28549 17632
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17660 31355 17663
rect 32861 17663 32919 17669
rect 31343 17632 31754 17660
rect 31343 17629 31355 17632
rect 31297 17623 31355 17629
rect 27433 17595 27491 17601
rect 27433 17561 27445 17595
rect 27479 17592 27491 17595
rect 28994 17592 29000 17604
rect 27479 17564 29000 17592
rect 27479 17561 27491 17564
rect 27433 17555 27491 17561
rect 28994 17552 29000 17564
rect 29052 17552 29058 17604
rect 29822 17592 29828 17604
rect 29783 17564 29828 17592
rect 29822 17552 29828 17564
rect 29880 17552 29886 17604
rect 29917 17595 29975 17601
rect 29917 17561 29929 17595
rect 29963 17561 29975 17595
rect 31726 17592 31754 17632
rect 32861 17629 32873 17663
rect 32907 17629 32919 17663
rect 33502 17660 33508 17672
rect 33463 17632 33508 17660
rect 32861 17623 32919 17629
rect 33502 17620 33508 17632
rect 33560 17620 33566 17672
rect 34146 17620 34152 17672
rect 34204 17660 34210 17672
rect 34204 17632 34249 17660
rect 34204 17620 34210 17632
rect 34790 17620 34796 17672
rect 34848 17660 34854 17672
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 34848 17632 34897 17660
rect 34848 17620 34854 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 37182 17660 37188 17672
rect 37143 17632 37188 17660
rect 34885 17623 34943 17629
rect 37182 17620 37188 17632
rect 37240 17620 37246 17672
rect 37826 17660 37832 17672
rect 37787 17632 37832 17660
rect 37826 17620 37832 17632
rect 37884 17620 37890 17672
rect 33410 17592 33416 17604
rect 31726 17564 33416 17592
rect 29917 17555 29975 17561
rect 14090 17524 14096 17536
rect 13188 17496 14096 17524
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14366 17524 14372 17536
rect 14327 17496 14372 17524
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 18785 17527 18843 17533
rect 18785 17524 18797 17527
rect 18564 17496 18797 17524
rect 18564 17484 18570 17496
rect 18785 17493 18797 17496
rect 18831 17493 18843 17527
rect 18785 17487 18843 17493
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 20070 17524 20076 17536
rect 19475 17496 20076 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 22922 17484 22928 17536
rect 22980 17524 22986 17536
rect 23109 17527 23167 17533
rect 23109 17524 23121 17527
rect 22980 17496 23121 17524
rect 22980 17484 22986 17496
rect 23109 17493 23121 17496
rect 23155 17493 23167 17527
rect 23109 17487 23167 17493
rect 26326 17484 26332 17536
rect 26384 17484 26390 17536
rect 27522 17484 27528 17536
rect 27580 17524 27586 17536
rect 29932 17524 29960 17555
rect 33410 17552 33416 17564
rect 33468 17552 33474 17604
rect 34241 17595 34299 17601
rect 34241 17561 34253 17595
rect 34287 17592 34299 17595
rect 35069 17595 35127 17601
rect 35069 17592 35081 17595
rect 34287 17564 35081 17592
rect 34287 17561 34299 17564
rect 34241 17555 34299 17561
rect 35069 17561 35081 17564
rect 35115 17561 35127 17595
rect 35069 17555 35127 17561
rect 27580 17496 29960 17524
rect 31389 17527 31447 17533
rect 27580 17484 27586 17496
rect 31389 17493 31401 17527
rect 31435 17524 31447 17527
rect 32858 17524 32864 17536
rect 31435 17496 32864 17524
rect 31435 17493 31447 17496
rect 31389 17487 31447 17493
rect 32858 17484 32864 17496
rect 32916 17484 32922 17536
rect 32953 17527 33011 17533
rect 32953 17493 32965 17527
rect 32999 17524 33011 17527
rect 33502 17524 33508 17536
rect 32999 17496 33508 17524
rect 32999 17493 33011 17496
rect 32953 17487 33011 17493
rect 33502 17484 33508 17496
rect 33560 17484 33566 17536
rect 33597 17527 33655 17533
rect 33597 17493 33609 17527
rect 33643 17524 33655 17527
rect 35342 17524 35348 17536
rect 33643 17496 35348 17524
rect 33643 17493 33655 17496
rect 33597 17487 33655 17493
rect 35342 17484 35348 17496
rect 35400 17484 35406 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 11204 17292 17785 17320
rect 11204 17280 11210 17292
rect 17773 17289 17785 17292
rect 17819 17289 17831 17323
rect 17773 17283 17831 17289
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 19300 17292 19349 17320
rect 19300 17280 19306 17292
rect 19337 17289 19349 17292
rect 19383 17289 19395 17323
rect 19337 17283 19395 17289
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 20496 17292 23980 17320
rect 20496 17280 20502 17292
rect 8846 17252 8852 17264
rect 8807 17224 8852 17252
rect 8846 17212 8852 17224
rect 8904 17212 8910 17264
rect 20070 17252 20076 17264
rect 20031 17224 20076 17252
rect 20070 17212 20076 17224
rect 20128 17212 20134 17264
rect 20625 17255 20683 17261
rect 20625 17221 20637 17255
rect 20671 17252 20683 17255
rect 21358 17252 21364 17264
rect 20671 17224 21364 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 21358 17212 21364 17224
rect 21416 17212 21422 17264
rect 22462 17212 22468 17264
rect 22520 17252 22526 17264
rect 22922 17252 22928 17264
rect 22520 17224 22928 17252
rect 22520 17212 22526 17224
rect 22922 17212 22928 17224
rect 22980 17212 22986 17264
rect 23017 17255 23075 17261
rect 23017 17221 23029 17255
rect 23063 17252 23075 17255
rect 23842 17252 23848 17264
rect 23063 17224 23848 17252
rect 23063 17221 23075 17224
rect 23017 17215 23075 17221
rect 23842 17212 23848 17224
rect 23900 17212 23906 17264
rect 23952 17261 23980 17292
rect 26142 17280 26148 17332
rect 26200 17320 26206 17332
rect 27249 17323 27307 17329
rect 27249 17320 27261 17323
rect 26200 17292 27261 17320
rect 26200 17280 26206 17292
rect 27249 17289 27261 17292
rect 27295 17289 27307 17323
rect 29178 17320 29184 17332
rect 29139 17292 29184 17320
rect 27249 17283 27307 17289
rect 29178 17280 29184 17292
rect 29236 17280 29242 17332
rect 32309 17323 32367 17329
rect 29840 17292 31754 17320
rect 23937 17255 23995 17261
rect 23937 17221 23949 17255
rect 23983 17221 23995 17255
rect 23937 17215 23995 17221
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17153 17739 17187
rect 19242 17184 19248 17196
rect 19203 17156 19248 17184
rect 17681 17147 17739 17153
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 8628 17088 8769 17116
rect 8628 17076 8634 17088
rect 8757 17085 8769 17088
rect 8803 17116 8815 17119
rect 9030 17116 9036 17128
rect 8803 17088 9036 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 9122 17076 9128 17128
rect 9180 17116 9186 17128
rect 9180 17088 9225 17116
rect 9180 17076 9186 17088
rect 17696 17048 17724 17147
rect 19242 17144 19248 17156
rect 19300 17144 19306 17196
rect 22002 17184 22008 17196
rect 21963 17156 22008 17184
rect 22002 17144 22008 17156
rect 22060 17144 22066 17196
rect 25682 17144 25688 17196
rect 25740 17184 25746 17196
rect 29840 17193 29868 17292
rect 30190 17212 30196 17264
rect 30248 17252 30254 17264
rect 30653 17255 30711 17261
rect 30653 17252 30665 17255
rect 30248 17224 30665 17252
rect 30248 17212 30254 17224
rect 30653 17221 30665 17224
rect 30699 17221 30711 17255
rect 30653 17215 30711 17221
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 25740 17156 27169 17184
rect 25740 17144 25746 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 29089 17187 29147 17193
rect 29089 17153 29101 17187
rect 29135 17153 29147 17187
rect 29089 17147 29147 17153
rect 29825 17187 29883 17193
rect 29825 17153 29837 17187
rect 29871 17153 29883 17187
rect 31726 17184 31754 17292
rect 32309 17289 32321 17323
rect 32355 17320 32367 17323
rect 32355 17292 38056 17320
rect 32355 17289 32367 17292
rect 32309 17283 32367 17289
rect 33502 17252 33508 17264
rect 33463 17224 33508 17252
rect 33502 17212 33508 17224
rect 33560 17212 33566 17264
rect 35342 17252 35348 17264
rect 35303 17224 35348 17252
rect 35342 17212 35348 17224
rect 35400 17212 35406 17264
rect 36817 17255 36875 17261
rect 36817 17221 36829 17255
rect 36863 17252 36875 17255
rect 37458 17252 37464 17264
rect 36863 17224 37464 17252
rect 36863 17221 36875 17224
rect 36817 17215 36875 17221
rect 37458 17212 37464 17224
rect 37516 17212 37522 17264
rect 32030 17184 32036 17196
rect 31726 17156 32036 17184
rect 29825 17147 29883 17153
rect 19978 17116 19984 17128
rect 19939 17088 19984 17116
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 21450 17048 21456 17060
rect 17696 17020 21456 17048
rect 21450 17008 21456 17020
rect 21508 17048 21514 17060
rect 24302 17048 24308 17060
rect 21508 17020 24308 17048
rect 21508 17008 21514 17020
rect 24302 17008 24308 17020
rect 24360 17008 24366 17060
rect 27172 17048 27200 17147
rect 29104 17116 29132 17147
rect 32030 17144 32036 17156
rect 32088 17184 32094 17196
rect 38028 17193 38056 17292
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 32088 17156 32505 17184
rect 32088 17144 32094 17156
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 32493 17147 32551 17153
rect 36725 17187 36783 17193
rect 36725 17153 36737 17187
rect 36771 17153 36783 17187
rect 36725 17147 36783 17153
rect 38013 17187 38071 17193
rect 38013 17153 38025 17187
rect 38059 17153 38071 17187
rect 38013 17147 38071 17153
rect 30282 17116 30288 17128
rect 29104 17088 30288 17116
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 30558 17116 30564 17128
rect 30519 17088 30564 17116
rect 30558 17076 30564 17088
rect 30616 17076 30622 17128
rect 31205 17119 31263 17125
rect 31205 17085 31217 17119
rect 31251 17116 31263 17119
rect 32122 17116 32128 17128
rect 31251 17088 32128 17116
rect 31251 17085 31263 17088
rect 31205 17079 31263 17085
rect 32122 17076 32128 17088
rect 32180 17076 32186 17128
rect 33413 17119 33471 17125
rect 33413 17085 33425 17119
rect 33459 17085 33471 17119
rect 33413 17079 33471 17085
rect 34057 17119 34115 17125
rect 34057 17085 34069 17119
rect 34103 17116 34115 17119
rect 34606 17116 34612 17128
rect 34103 17088 34612 17116
rect 34103 17085 34115 17088
rect 34057 17079 34115 17085
rect 27172 17020 30328 17048
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16980 1639 16983
rect 9766 16980 9772 16992
rect 1627 16952 9772 16980
rect 1627 16949 1639 16952
rect 1581 16943 1639 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 20990 16940 20996 16992
rect 21048 16980 21054 16992
rect 22097 16983 22155 16989
rect 22097 16980 22109 16983
rect 21048 16952 22109 16980
rect 21048 16940 21054 16952
rect 22097 16949 22109 16952
rect 22143 16949 22155 16983
rect 29914 16980 29920 16992
rect 29875 16952 29920 16980
rect 22097 16943 22155 16949
rect 29914 16940 29920 16952
rect 29972 16940 29978 16992
rect 30300 16980 30328 17020
rect 30374 17008 30380 17060
rect 30432 17048 30438 17060
rect 33428 17048 33456 17079
rect 34606 17076 34612 17088
rect 34664 17076 34670 17128
rect 35253 17119 35311 17125
rect 35253 17085 35265 17119
rect 35299 17116 35311 17119
rect 35342 17116 35348 17128
rect 35299 17088 35348 17116
rect 35299 17085 35311 17088
rect 35253 17079 35311 17085
rect 35342 17076 35348 17088
rect 35400 17076 35406 17128
rect 36078 17116 36084 17128
rect 36039 17088 36084 17116
rect 36078 17076 36084 17088
rect 36136 17116 36142 17128
rect 36354 17116 36360 17128
rect 36136 17088 36360 17116
rect 36136 17076 36142 17088
rect 36354 17076 36360 17088
rect 36412 17076 36418 17128
rect 30432 17020 33456 17048
rect 30432 17008 30438 17020
rect 31110 16980 31116 16992
rect 30300 16952 31116 16980
rect 31110 16940 31116 16952
rect 31168 16940 31174 16992
rect 33042 16940 33048 16992
rect 33100 16980 33106 16992
rect 36740 16980 36768 17147
rect 38194 17048 38200 17060
rect 38155 17020 38200 17048
rect 38194 17008 38200 17020
rect 38252 17008 38258 17060
rect 33100 16952 36768 16980
rect 33100 16940 33106 16952
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 27430 16776 27436 16788
rect 19300 16748 27436 16776
rect 19300 16736 19306 16748
rect 27430 16736 27436 16748
rect 27488 16736 27494 16788
rect 28258 16776 28264 16788
rect 28171 16748 28264 16776
rect 28258 16736 28264 16748
rect 28316 16776 28322 16788
rect 31018 16776 31024 16788
rect 28316 16748 31024 16776
rect 28316 16736 28322 16748
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 35253 16779 35311 16785
rect 35253 16776 35265 16779
rect 34848 16748 35265 16776
rect 34848 16736 34854 16748
rect 35253 16745 35265 16748
rect 35299 16745 35311 16779
rect 39390 16776 39396 16788
rect 35253 16739 35311 16745
rect 36372 16748 39396 16776
rect 23658 16668 23664 16720
rect 23716 16708 23722 16720
rect 28276 16708 28304 16736
rect 23716 16680 28304 16708
rect 23716 16668 23722 16680
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 14458 16640 14464 16652
rect 13596 16612 14464 16640
rect 13596 16600 13602 16612
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20220 16612 20576 16640
rect 20220 16600 20226 16612
rect 20548 16581 20576 16612
rect 22738 16600 22744 16652
rect 22796 16640 22802 16652
rect 23474 16640 23480 16652
rect 22796 16612 23480 16640
rect 22796 16600 22802 16612
rect 23474 16600 23480 16612
rect 23532 16640 23538 16652
rect 25961 16643 26019 16649
rect 23532 16612 25360 16640
rect 23532 16600 23538 16612
rect 21169 16585 21227 16591
rect 21169 16584 21181 16585
rect 21215 16584 21227 16585
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 21169 16545 21180 16584
rect 20533 16535 20591 16541
rect 21174 16532 21180 16545
rect 21232 16532 21238 16584
rect 21542 16532 21548 16584
rect 21600 16572 21606 16584
rect 21600 16544 23152 16572
rect 21600 16532 21606 16544
rect 20625 16507 20683 16513
rect 20625 16473 20637 16507
rect 20671 16504 20683 16507
rect 22186 16504 22192 16516
rect 20671 16476 22192 16504
rect 20671 16473 20683 16476
rect 20625 16467 20683 16473
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 23124 16504 23152 16544
rect 23198 16532 23204 16584
rect 23256 16572 23262 16584
rect 25332 16581 25360 16612
rect 25961 16609 25973 16643
rect 26007 16640 26019 16643
rect 26326 16640 26332 16652
rect 26007 16612 26332 16640
rect 26007 16609 26019 16612
rect 25961 16603 26019 16609
rect 26326 16600 26332 16612
rect 26384 16600 26390 16652
rect 26436 16649 26464 16680
rect 28350 16668 28356 16720
rect 28408 16708 28414 16720
rect 34882 16708 34888 16720
rect 28408 16680 30236 16708
rect 28408 16668 28414 16680
rect 26421 16643 26479 16649
rect 26421 16609 26433 16643
rect 26467 16609 26479 16643
rect 26421 16603 26479 16609
rect 27338 16600 27344 16652
rect 27396 16640 27402 16652
rect 29086 16640 29092 16652
rect 27396 16612 28304 16640
rect 27396 16600 27402 16612
rect 28276 16581 28304 16612
rect 28920 16612 29092 16640
rect 28920 16581 28948 16612
rect 29086 16600 29092 16612
rect 29144 16600 29150 16652
rect 30208 16649 30236 16680
rect 31772 16680 34888 16708
rect 30193 16643 30251 16649
rect 30193 16609 30205 16643
rect 30239 16609 30251 16643
rect 30193 16603 30251 16609
rect 30837 16643 30895 16649
rect 30837 16609 30849 16643
rect 30883 16640 30895 16643
rect 31386 16640 31392 16652
rect 30883 16612 31392 16640
rect 30883 16609 30895 16612
rect 30837 16603 30895 16609
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 31772 16649 31800 16680
rect 34882 16668 34888 16680
rect 34940 16708 34946 16720
rect 35710 16708 35716 16720
rect 34940 16680 35716 16708
rect 34940 16668 34946 16680
rect 35710 16668 35716 16680
rect 35768 16668 35774 16720
rect 31757 16643 31815 16649
rect 31757 16609 31769 16643
rect 31803 16609 31815 16643
rect 31757 16603 31815 16609
rect 33321 16643 33379 16649
rect 33321 16609 33333 16643
rect 33367 16640 33379 16643
rect 35342 16640 35348 16652
rect 33367 16612 35348 16640
rect 33367 16609 33379 16612
rect 33321 16603 33379 16609
rect 35342 16600 35348 16612
rect 35400 16600 35406 16652
rect 36372 16640 36400 16748
rect 39390 16736 39396 16748
rect 39448 16736 39454 16788
rect 38102 16708 38108 16720
rect 35452 16612 36400 16640
rect 36464 16680 38108 16708
rect 25317 16575 25375 16581
rect 23256 16544 23301 16572
rect 23256 16532 23262 16544
rect 25317 16541 25329 16575
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 28261 16575 28319 16581
rect 28261 16541 28273 16575
rect 28307 16541 28319 16575
rect 28261 16535 28319 16541
rect 28905 16575 28963 16581
rect 28905 16541 28917 16575
rect 28951 16541 28963 16575
rect 28905 16535 28963 16541
rect 35161 16575 35219 16581
rect 35161 16541 35173 16575
rect 35207 16572 35219 16575
rect 35452 16572 35480 16612
rect 35986 16572 35992 16584
rect 35207 16544 35480 16572
rect 35947 16544 35992 16572
rect 35207 16541 35219 16544
rect 35161 16535 35219 16541
rect 35986 16532 35992 16544
rect 36044 16532 36050 16584
rect 36464 16581 36492 16680
rect 38102 16668 38108 16680
rect 38160 16668 38166 16720
rect 39298 16640 39304 16652
rect 37752 16612 39304 16640
rect 36449 16575 36507 16581
rect 36449 16541 36461 16575
rect 36495 16541 36507 16575
rect 36449 16535 36507 16541
rect 36998 16532 37004 16584
rect 37056 16572 37062 16584
rect 37752 16581 37780 16612
rect 39298 16600 39304 16612
rect 39356 16600 39362 16652
rect 37285 16575 37343 16581
rect 37285 16572 37297 16575
rect 37056 16544 37297 16572
rect 37056 16532 37062 16544
rect 37285 16541 37297 16544
rect 37331 16572 37343 16575
rect 37737 16575 37795 16581
rect 37331 16544 37596 16572
rect 37331 16541 37343 16544
rect 37285 16535 37343 16541
rect 25409 16507 25467 16513
rect 23124 16476 23704 16504
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 20162 16436 20168 16448
rect 11940 16408 20168 16436
rect 11940 16396 11946 16408
rect 20162 16396 20168 16408
rect 20220 16396 20226 16448
rect 21269 16439 21327 16445
rect 21269 16405 21281 16439
rect 21315 16436 21327 16439
rect 22646 16436 22652 16448
rect 21315 16408 22652 16436
rect 21315 16405 21327 16408
rect 21269 16399 21327 16405
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 23293 16439 23351 16445
rect 23293 16405 23305 16439
rect 23339 16436 23351 16439
rect 23566 16436 23572 16448
rect 23339 16408 23572 16436
rect 23339 16405 23351 16408
rect 23293 16399 23351 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 23676 16436 23704 16476
rect 25409 16473 25421 16507
rect 25455 16504 25467 16507
rect 26145 16507 26203 16513
rect 26145 16504 26157 16507
rect 25455 16476 26157 16504
rect 25455 16473 25467 16476
rect 25409 16467 25467 16473
rect 26145 16473 26157 16476
rect 26191 16473 26203 16507
rect 26145 16467 26203 16473
rect 30282 16464 30288 16516
rect 30340 16504 30346 16516
rect 30340 16476 30385 16504
rect 30340 16464 30346 16476
rect 31846 16464 31852 16516
rect 31904 16504 31910 16516
rect 32766 16504 32772 16516
rect 31904 16476 31949 16504
rect 32727 16476 32772 16504
rect 31904 16464 31910 16476
rect 32766 16464 32772 16476
rect 32824 16464 32830 16516
rect 32858 16464 32864 16516
rect 32916 16504 32922 16516
rect 33413 16507 33471 16513
rect 33413 16504 33425 16507
rect 32916 16476 33425 16504
rect 32916 16464 32922 16476
rect 33413 16473 33425 16476
rect 33459 16473 33471 16507
rect 34330 16504 34336 16516
rect 34291 16476 34336 16504
rect 33413 16467 33471 16473
rect 34330 16464 34336 16476
rect 34388 16464 34394 16516
rect 36541 16507 36599 16513
rect 36541 16504 36553 16507
rect 34440 16476 36553 16504
rect 27246 16436 27252 16448
rect 23676 16408 27252 16436
rect 27246 16396 27252 16408
rect 27304 16396 27310 16448
rect 27614 16396 27620 16448
rect 27672 16436 27678 16448
rect 28353 16439 28411 16445
rect 28353 16436 28365 16439
rect 27672 16408 28365 16436
rect 27672 16396 27678 16408
rect 28353 16405 28365 16408
rect 28399 16405 28411 16439
rect 28353 16399 28411 16405
rect 28997 16439 29055 16445
rect 28997 16405 29009 16439
rect 29043 16436 29055 16439
rect 29454 16436 29460 16448
rect 29043 16408 29460 16436
rect 29043 16405 29055 16408
rect 28997 16399 29055 16405
rect 29454 16396 29460 16408
rect 29512 16396 29518 16448
rect 29822 16396 29828 16448
rect 29880 16436 29886 16448
rect 34440 16436 34468 16476
rect 36541 16473 36553 16476
rect 36587 16473 36599 16507
rect 37568 16504 37596 16544
rect 37737 16541 37749 16575
rect 37783 16541 37795 16575
rect 37737 16535 37795 16541
rect 37829 16575 37887 16581
rect 37829 16541 37841 16575
rect 37875 16572 37887 16575
rect 37918 16572 37924 16584
rect 37875 16544 37924 16572
rect 37875 16541 37887 16544
rect 37829 16535 37887 16541
rect 37918 16532 37924 16544
rect 37976 16532 37982 16584
rect 38746 16504 38752 16516
rect 37568 16476 38752 16504
rect 36541 16467 36599 16473
rect 38746 16464 38752 16476
rect 38804 16464 38810 16516
rect 29880 16408 34468 16436
rect 29880 16396 29886 16408
rect 35526 16396 35532 16448
rect 35584 16436 35590 16448
rect 35805 16439 35863 16445
rect 35805 16436 35817 16439
rect 35584 16408 35817 16436
rect 35584 16396 35590 16408
rect 35805 16405 35817 16408
rect 35851 16405 35863 16439
rect 35805 16399 35863 16405
rect 37093 16439 37151 16445
rect 37093 16405 37105 16439
rect 37139 16436 37151 16439
rect 37642 16436 37648 16448
rect 37139 16408 37648 16436
rect 37139 16405 37151 16408
rect 37093 16399 37151 16405
rect 37642 16396 37648 16408
rect 37700 16396 37706 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 15010 16232 15016 16244
rect 13780 16204 15016 16232
rect 13780 16192 13786 16204
rect 15010 16192 15016 16204
rect 15068 16232 15074 16244
rect 15068 16204 18644 16232
rect 15068 16192 15074 16204
rect 17034 16164 17040 16176
rect 16995 16136 17040 16164
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 18506 16164 18512 16176
rect 18467 16136 18512 16164
rect 18506 16124 18512 16136
rect 18564 16124 18570 16176
rect 18616 16164 18644 16204
rect 18966 16192 18972 16244
rect 19024 16232 19030 16244
rect 22094 16232 22100 16244
rect 19024 16204 22100 16232
rect 19024 16192 19030 16204
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 25590 16232 25596 16244
rect 23768 16204 25596 16232
rect 19061 16167 19119 16173
rect 19061 16164 19073 16167
rect 18616 16136 19073 16164
rect 19061 16133 19073 16136
rect 19107 16133 19119 16167
rect 22112 16164 22140 16192
rect 22112 16136 23152 16164
rect 19061 16127 19119 16133
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 6733 16099 6791 16105
rect 1627 16068 2774 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 2746 15960 2774 16068
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 7926 16096 7932 16108
rect 7887 16068 7932 16096
rect 6733 16059 6791 16065
rect 6748 16028 6776 16059
rect 7926 16056 7932 16068
rect 7984 16056 7990 16108
rect 22370 16096 22376 16108
rect 20732 16068 22376 16096
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 6748 16000 8033 16028
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 12250 15988 12256 16040
rect 12308 16028 12314 16040
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 12308 16000 16957 16028
rect 12308 15988 12314 16000
rect 16945 15997 16957 16000
rect 16991 16028 17003 16031
rect 17770 16028 17776 16040
rect 16991 16000 17776 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 18417 16031 18475 16037
rect 18417 15997 18429 16031
rect 18463 16028 18475 16031
rect 20732 16028 20760 16068
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 23124 16105 23152 16136
rect 23768 16105 23796 16204
rect 25590 16192 25596 16204
rect 25648 16192 25654 16244
rect 29822 16232 29828 16244
rect 26160 16204 29828 16232
rect 25314 16164 25320 16176
rect 25275 16136 25320 16164
rect 25314 16124 25320 16136
rect 25372 16124 25378 16176
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 18463 16000 20760 16028
rect 20809 16031 20867 16037
rect 18463 15997 18475 16000
rect 18417 15991 18475 15997
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20990 16028 20996 16040
rect 20951 16000 20996 16028
rect 20809 15991 20867 15997
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 2746 15932 6561 15960
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 6549 15923 6607 15929
rect 15102 15920 15108 15972
rect 15160 15960 15166 15972
rect 17494 15960 17500 15972
rect 15160 15932 17500 15960
rect 15160 15920 15166 15932
rect 17494 15920 17500 15932
rect 17552 15920 17558 15972
rect 1762 15892 1768 15904
rect 1723 15864 1768 15892
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 20824 15892 20852 15991
rect 20990 15988 20996 16000
rect 21048 15988 21054 16040
rect 22278 15988 22284 16040
rect 22336 16028 22342 16040
rect 25225 16031 25283 16037
rect 22336 16000 23980 16028
rect 22336 15988 22342 16000
rect 23952 15972 23980 16000
rect 25225 15997 25237 16031
rect 25271 16028 25283 16031
rect 26160 16028 26188 16204
rect 29822 16192 29828 16204
rect 29880 16192 29886 16244
rect 30282 16192 30288 16244
rect 30340 16232 30346 16244
rect 30929 16235 30987 16241
rect 30929 16232 30941 16235
rect 30340 16204 30941 16232
rect 30340 16192 30346 16204
rect 30929 16201 30941 16204
rect 30975 16201 30987 16235
rect 30929 16195 30987 16201
rect 31481 16235 31539 16241
rect 31481 16201 31493 16235
rect 31527 16232 31539 16235
rect 31527 16204 31754 16232
rect 31527 16201 31539 16204
rect 31481 16195 31539 16201
rect 27798 16164 27804 16176
rect 27759 16136 27804 16164
rect 27798 16124 27804 16136
rect 27856 16124 27862 16176
rect 27982 16124 27988 16176
rect 28040 16164 28046 16176
rect 28353 16167 28411 16173
rect 28353 16164 28365 16167
rect 28040 16136 28365 16164
rect 28040 16124 28046 16136
rect 28353 16133 28365 16136
rect 28399 16164 28411 16167
rect 28442 16164 28448 16176
rect 28399 16136 28448 16164
rect 28399 16133 28411 16136
rect 28353 16127 28411 16133
rect 28442 16124 28448 16136
rect 28500 16124 28506 16176
rect 29454 16164 29460 16176
rect 29415 16136 29460 16164
rect 29454 16124 29460 16136
rect 29512 16124 29518 16176
rect 31570 16164 31576 16176
rect 30852 16136 31576 16164
rect 30852 16105 30880 16136
rect 31570 16124 31576 16136
rect 31628 16124 31634 16176
rect 31726 16164 31754 16204
rect 35986 16192 35992 16244
rect 36044 16232 36050 16244
rect 36817 16235 36875 16241
rect 36817 16232 36829 16235
rect 36044 16204 36829 16232
rect 36044 16192 36050 16204
rect 36817 16201 36829 16204
rect 36863 16201 36875 16235
rect 36817 16195 36875 16201
rect 32493 16167 32551 16173
rect 32493 16164 32505 16167
rect 31726 16136 32505 16164
rect 32493 16133 32505 16136
rect 32539 16133 32551 16167
rect 32493 16127 32551 16133
rect 32674 16124 32680 16176
rect 32732 16164 32738 16176
rect 34422 16164 34428 16176
rect 32732 16136 33548 16164
rect 34383 16136 34428 16164
rect 32732 16124 32738 16136
rect 30837 16099 30895 16105
rect 30837 16065 30849 16099
rect 30883 16065 30895 16099
rect 30837 16059 30895 16065
rect 31018 16056 31024 16108
rect 31076 16096 31082 16108
rect 33520 16105 33548 16136
rect 34422 16124 34428 16136
rect 34480 16124 34486 16176
rect 34514 16124 34520 16176
rect 34572 16164 34578 16176
rect 36173 16167 36231 16173
rect 34572 16136 36124 16164
rect 34572 16124 34578 16136
rect 31665 16099 31723 16105
rect 31665 16096 31677 16099
rect 31076 16068 31677 16096
rect 31076 16056 31082 16068
rect 31665 16065 31677 16068
rect 31711 16065 31723 16099
rect 31665 16059 31723 16065
rect 33505 16099 33563 16105
rect 33505 16065 33517 16099
rect 33551 16065 33563 16099
rect 33505 16059 33563 16065
rect 35437 16099 35495 16105
rect 35437 16065 35449 16099
rect 35483 16096 35495 16099
rect 35618 16096 35624 16108
rect 35483 16068 35624 16096
rect 35483 16065 35495 16068
rect 35437 16059 35495 16065
rect 35618 16056 35624 16068
rect 35676 16056 35682 16108
rect 36096 16105 36124 16136
rect 36173 16133 36185 16167
rect 36219 16164 36231 16167
rect 37366 16164 37372 16176
rect 36219 16136 37372 16164
rect 36219 16133 36231 16136
rect 36173 16127 36231 16133
rect 37366 16124 37372 16136
rect 37424 16124 37430 16176
rect 36081 16099 36139 16105
rect 36081 16065 36093 16099
rect 36127 16065 36139 16099
rect 36722 16096 36728 16108
rect 36683 16068 36728 16096
rect 36081 16059 36139 16065
rect 36722 16056 36728 16068
rect 36780 16056 36786 16108
rect 38010 16096 38016 16108
rect 37971 16068 38016 16096
rect 38010 16056 38016 16068
rect 38068 16056 38074 16108
rect 25271 16000 26188 16028
rect 26237 16031 26295 16037
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 26237 15997 26249 16031
rect 26283 15997 26295 16031
rect 26237 15991 26295 15997
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 16028 27767 16031
rect 29365 16031 29423 16037
rect 27755 16000 29316 16028
rect 27755 15997 27767 16000
rect 27709 15991 27767 15997
rect 21266 15920 21272 15972
rect 21324 15960 21330 15972
rect 23845 15963 23903 15969
rect 23845 15960 23857 15963
rect 21324 15932 23857 15960
rect 21324 15920 21330 15932
rect 23845 15929 23857 15932
rect 23891 15929 23903 15963
rect 23845 15923 23903 15929
rect 23934 15920 23940 15972
rect 23992 15960 23998 15972
rect 26252 15960 26280 15991
rect 23992 15932 26280 15960
rect 29288 15960 29316 16000
rect 29365 15997 29377 16031
rect 29411 16028 29423 16031
rect 29454 16028 29460 16040
rect 29411 16000 29460 16028
rect 29411 15997 29423 16000
rect 29365 15991 29423 15997
rect 29454 15988 29460 16000
rect 29512 16028 29518 16040
rect 29914 16028 29920 16040
rect 29512 16000 29920 16028
rect 29512 15988 29518 16000
rect 29914 15988 29920 16000
rect 29972 15988 29978 16040
rect 30285 16031 30343 16037
rect 30285 15997 30297 16031
rect 30331 16028 30343 16031
rect 30374 16028 30380 16040
rect 30331 16000 30380 16028
rect 30331 15997 30343 16000
rect 30285 15991 30343 15997
rect 30374 15988 30380 16000
rect 30432 15988 30438 16040
rect 32401 16031 32459 16037
rect 32401 16028 32413 16031
rect 31726 16000 32413 16028
rect 31726 15960 31754 16000
rect 32401 15997 32413 16000
rect 32447 15997 32459 16031
rect 33042 16028 33048 16040
rect 32955 16000 33048 16028
rect 32401 15991 32459 15997
rect 29288 15932 31754 15960
rect 32416 15960 32444 15991
rect 33042 15988 33048 16000
rect 33100 16028 33106 16040
rect 34333 16031 34391 16037
rect 34333 16028 34345 16031
rect 33100 16000 34345 16028
rect 33100 15988 33106 16000
rect 34333 15997 34345 16000
rect 34379 15997 34391 16031
rect 34333 15991 34391 15997
rect 34977 16031 35035 16037
rect 34977 15997 34989 16031
rect 35023 16028 35035 16031
rect 36740 16028 36768 16056
rect 35023 16000 36768 16028
rect 35023 15997 35035 16000
rect 34977 15991 35035 15997
rect 34514 15960 34520 15972
rect 32416 15932 34520 15960
rect 23992 15920 23998 15932
rect 34514 15920 34520 15932
rect 34572 15920 34578 15972
rect 35529 15963 35587 15969
rect 35529 15929 35541 15963
rect 35575 15960 35587 15963
rect 37642 15960 37648 15972
rect 35575 15932 37648 15960
rect 35575 15929 35587 15932
rect 35529 15923 35587 15929
rect 37642 15920 37648 15932
rect 37700 15920 37706 15972
rect 21174 15892 21180 15904
rect 12492 15864 20852 15892
rect 21135 15864 21180 15892
rect 12492 15852 12498 15864
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 23201 15895 23259 15901
rect 23201 15861 23213 15895
rect 23247 15892 23259 15895
rect 24670 15892 24676 15904
rect 23247 15864 24676 15892
rect 23247 15861 23259 15864
rect 23201 15855 23259 15861
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 25958 15852 25964 15904
rect 26016 15892 26022 15904
rect 26786 15892 26792 15904
rect 26016 15864 26792 15892
rect 26016 15852 26022 15864
rect 26786 15852 26792 15864
rect 26844 15852 26850 15904
rect 27430 15852 27436 15904
rect 27488 15892 27494 15904
rect 30926 15892 30932 15904
rect 27488 15864 30932 15892
rect 27488 15852 27494 15864
rect 30926 15852 30932 15864
rect 30984 15852 30990 15904
rect 33597 15895 33655 15901
rect 33597 15861 33609 15895
rect 33643 15892 33655 15895
rect 37090 15892 37096 15904
rect 33643 15864 37096 15892
rect 33643 15861 33655 15864
rect 33597 15855 33655 15861
rect 37090 15852 37096 15864
rect 37148 15852 37154 15904
rect 38194 15892 38200 15904
rect 38155 15864 38200 15892
rect 38194 15852 38200 15864
rect 38252 15852 38258 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 11756 15660 19334 15688
rect 11756 15648 11762 15660
rect 19306 15620 19334 15660
rect 23400 15660 23980 15688
rect 23400 15620 23428 15660
rect 23952 15620 23980 15660
rect 24026 15648 24032 15700
rect 24084 15688 24090 15700
rect 25222 15688 25228 15700
rect 24084 15660 25228 15688
rect 24084 15648 24090 15660
rect 25222 15648 25228 15660
rect 25280 15688 25286 15700
rect 26142 15688 26148 15700
rect 25280 15660 26148 15688
rect 25280 15648 25286 15660
rect 26142 15648 26148 15660
rect 26200 15648 26206 15700
rect 26237 15691 26295 15697
rect 26237 15657 26249 15691
rect 26283 15688 26295 15691
rect 27798 15688 27804 15700
rect 26283 15660 27804 15688
rect 26283 15657 26295 15660
rect 26237 15651 26295 15657
rect 27798 15648 27804 15660
rect 27856 15648 27862 15700
rect 27893 15691 27951 15697
rect 27893 15657 27905 15691
rect 27939 15688 27951 15691
rect 29270 15688 29276 15700
rect 27939 15660 29276 15688
rect 27939 15657 27951 15660
rect 27893 15651 27951 15657
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 31018 15688 31024 15700
rect 30979 15660 31024 15688
rect 31018 15648 31024 15660
rect 31076 15648 31082 15700
rect 34514 15648 34520 15700
rect 34572 15688 34578 15700
rect 35618 15688 35624 15700
rect 34572 15660 35624 15688
rect 34572 15648 34578 15660
rect 35618 15648 35624 15660
rect 35676 15648 35682 15700
rect 33042 15620 33048 15632
rect 19306 15592 23428 15620
rect 23492 15592 23704 15620
rect 23952 15592 33048 15620
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15552 11391 15555
rect 13170 15552 13176 15564
rect 11379 15524 13176 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 23492 15552 23520 15592
rect 16592 15524 23520 15552
rect 23676 15552 23704 15592
rect 33042 15580 33048 15592
rect 33100 15580 33106 15632
rect 23676 15524 31800 15552
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15484 6883 15487
rect 8754 15484 8760 15496
rect 6871 15456 8760 15484
rect 6871 15453 6883 15456
rect 6825 15447 6883 15453
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 15909 15487 15967 15493
rect 15909 15484 15921 15487
rect 14608 15456 15921 15484
rect 14608 15444 14614 15456
rect 15909 15453 15921 15456
rect 15955 15484 15967 15487
rect 16592 15484 16620 15524
rect 23593 15497 23651 15503
rect 15955 15456 16620 15484
rect 15955 15453 15967 15456
rect 15909 15447 15967 15453
rect 16758 15444 16764 15496
rect 16816 15484 16822 15496
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 16816 15456 20545 15484
rect 16816 15444 16822 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20622 15444 20628 15496
rect 20680 15484 20686 15496
rect 22278 15484 22284 15496
rect 20680 15456 22284 15484
rect 20680 15444 20686 15456
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 22462 15484 22468 15496
rect 22423 15456 22468 15484
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 22646 15484 22652 15496
rect 22607 15456 22652 15484
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23593 15463 23605 15497
rect 23639 15494 23651 15497
rect 23639 15484 23796 15494
rect 24210 15484 24216 15496
rect 23639 15466 24216 15484
rect 23639 15463 23651 15466
rect 23593 15457 23651 15463
rect 23768 15456 24216 15466
rect 24210 15444 24216 15456
rect 24268 15444 24274 15496
rect 24578 15484 24584 15496
rect 24539 15456 24584 15484
rect 24578 15444 24584 15456
rect 24636 15444 24642 15496
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15484 25559 15487
rect 25958 15484 25964 15496
rect 25547 15456 25964 15484
rect 25547 15453 25559 15456
rect 25501 15447 25559 15453
rect 25958 15444 25964 15456
rect 26016 15444 26022 15496
rect 26142 15444 26148 15496
rect 26200 15484 26206 15496
rect 27246 15484 27252 15496
rect 26200 15456 26245 15484
rect 27207 15456 27252 15484
rect 26200 15444 26206 15456
rect 27246 15444 27252 15456
rect 27304 15444 27310 15496
rect 27433 15487 27491 15493
rect 27433 15453 27445 15487
rect 27479 15484 27491 15487
rect 28166 15484 28172 15496
rect 27479 15456 28172 15484
rect 27479 15453 27491 15456
rect 27433 15447 27491 15453
rect 28166 15444 28172 15456
rect 28224 15444 28230 15496
rect 29178 15444 29184 15496
rect 29236 15484 29242 15496
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29236 15456 29929 15484
rect 29236 15444 29242 15456
rect 29917 15453 29929 15456
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 30377 15487 30435 15493
rect 30377 15453 30389 15487
rect 30423 15484 30435 15487
rect 30926 15484 30932 15496
rect 30423 15456 30932 15484
rect 30423 15453 30435 15456
rect 30377 15447 30435 15453
rect 30926 15444 30932 15456
rect 30984 15444 30990 15496
rect 31202 15484 31208 15496
rect 31163 15456 31208 15484
rect 31202 15444 31208 15456
rect 31260 15444 31266 15496
rect 31662 15484 31668 15496
rect 31623 15456 31668 15484
rect 31662 15444 31668 15456
rect 31720 15444 31726 15496
rect 31772 15484 31800 15524
rect 31846 15512 31852 15564
rect 31904 15552 31910 15564
rect 33965 15555 34023 15561
rect 33965 15552 33977 15555
rect 31904 15524 33088 15552
rect 31904 15512 31910 15524
rect 31938 15484 31944 15496
rect 31772 15456 31944 15484
rect 31938 15444 31944 15456
rect 31996 15484 32002 15496
rect 32309 15487 32367 15493
rect 32309 15484 32321 15487
rect 31996 15456 32321 15484
rect 31996 15444 32002 15456
rect 32309 15453 32321 15456
rect 32355 15484 32367 15487
rect 32766 15484 32772 15496
rect 32355 15456 32772 15484
rect 32355 15453 32367 15456
rect 32309 15447 32367 15453
rect 32766 15444 32772 15456
rect 32824 15444 32830 15496
rect 32950 15484 32956 15496
rect 32911 15456 32956 15484
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 33060 15493 33088 15524
rect 33428 15524 33977 15552
rect 33045 15487 33103 15493
rect 33045 15453 33057 15487
rect 33091 15453 33103 15487
rect 33045 15447 33103 15453
rect 10318 15416 10324 15428
rect 10279 15388 10324 15416
rect 10318 15376 10324 15388
rect 10376 15376 10382 15428
rect 10410 15376 10416 15428
rect 10468 15416 10474 15428
rect 10468 15388 10513 15416
rect 10468 15376 10474 15388
rect 12710 15376 12716 15428
rect 12768 15416 12774 15428
rect 17218 15416 17224 15428
rect 12768 15388 17224 15416
rect 12768 15376 12774 15388
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 17494 15376 17500 15428
rect 17552 15416 17558 15428
rect 23290 15416 23296 15428
rect 17552 15388 23296 15416
rect 17552 15376 17558 15388
rect 23290 15376 23296 15388
rect 23348 15376 23354 15428
rect 28442 15416 28448 15428
rect 28403 15388 28448 15416
rect 28442 15376 28448 15388
rect 28500 15376 28506 15428
rect 28537 15419 28595 15425
rect 28537 15385 28549 15419
rect 28583 15416 28595 15419
rect 28902 15416 28908 15428
rect 28583 15388 28908 15416
rect 28583 15385 28595 15388
rect 28537 15379 28595 15385
rect 28902 15376 28908 15388
rect 28960 15376 28966 15428
rect 29089 15419 29147 15425
rect 29089 15385 29101 15419
rect 29135 15416 29147 15419
rect 33428 15416 33456 15524
rect 33965 15521 33977 15524
rect 34011 15552 34023 15555
rect 34146 15552 34152 15564
rect 34011 15524 34152 15552
rect 34011 15521 34023 15524
rect 33965 15515 34023 15521
rect 34146 15512 34152 15524
rect 34204 15512 34210 15564
rect 36630 15552 36636 15564
rect 34900 15524 36636 15552
rect 34900 15493 34928 15524
rect 36630 15512 36636 15524
rect 36688 15512 36694 15564
rect 37001 15555 37059 15561
rect 37001 15521 37013 15555
rect 37047 15552 37059 15555
rect 37550 15552 37556 15564
rect 37047 15524 37556 15552
rect 37047 15521 37059 15524
rect 37001 15515 37059 15521
rect 37550 15512 37556 15524
rect 37608 15552 37614 15564
rect 37829 15555 37887 15561
rect 37829 15552 37841 15555
rect 37608 15524 37841 15552
rect 37608 15512 37614 15524
rect 37829 15521 37841 15524
rect 37875 15521 37887 15555
rect 37829 15515 37887 15521
rect 34885 15487 34943 15493
rect 34885 15453 34897 15487
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15484 35771 15487
rect 35894 15484 35900 15496
rect 35759 15456 35900 15484
rect 35759 15453 35771 15456
rect 35713 15447 35771 15453
rect 35894 15444 35900 15456
rect 35952 15444 35958 15496
rect 33686 15416 33692 15428
rect 29135 15388 33456 15416
rect 33647 15388 33692 15416
rect 29135 15385 29147 15388
rect 29089 15379 29147 15385
rect 33686 15376 33692 15388
rect 33744 15376 33750 15428
rect 33781 15419 33839 15425
rect 33781 15385 33793 15419
rect 33827 15385 33839 15419
rect 33781 15379 33839 15385
rect 34977 15419 35035 15425
rect 34977 15385 34989 15419
rect 35023 15416 35035 15419
rect 36354 15416 36360 15428
rect 35023 15388 36124 15416
rect 36315 15388 36360 15416
rect 35023 15385 35035 15388
rect 34977 15379 35035 15385
rect 1762 15308 1768 15360
rect 1820 15348 1826 15360
rect 6641 15351 6699 15357
rect 6641 15348 6653 15351
rect 1820 15320 6653 15348
rect 1820 15308 1826 15320
rect 6641 15317 6653 15320
rect 6687 15317 6699 15351
rect 6641 15311 6699 15317
rect 15749 15351 15807 15357
rect 15749 15317 15761 15351
rect 15795 15348 15807 15351
rect 16298 15348 16304 15360
rect 15795 15320 16304 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 17236 15348 17264 15376
rect 20530 15348 20536 15360
rect 17236 15320 20536 15348
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 20625 15351 20683 15357
rect 20625 15317 20637 15351
rect 20671 15348 20683 15351
rect 21634 15348 21640 15360
rect 20671 15320 21640 15348
rect 20671 15317 20683 15320
rect 20625 15311 20683 15317
rect 21634 15308 21640 15320
rect 21692 15308 21698 15360
rect 23106 15348 23112 15360
rect 23067 15320 23112 15348
rect 23106 15308 23112 15320
rect 23164 15308 23170 15360
rect 23198 15308 23204 15360
rect 23256 15348 23262 15360
rect 23661 15351 23719 15357
rect 23661 15348 23673 15351
rect 23256 15320 23673 15348
rect 23256 15308 23262 15320
rect 23661 15317 23673 15320
rect 23707 15317 23719 15351
rect 23661 15311 23719 15317
rect 24673 15351 24731 15357
rect 24673 15317 24685 15351
rect 24719 15348 24731 15351
rect 25406 15348 25412 15360
rect 24719 15320 25412 15348
rect 24719 15317 24731 15320
rect 24673 15311 24731 15317
rect 25406 15308 25412 15320
rect 25464 15308 25470 15360
rect 25593 15351 25651 15357
rect 25593 15317 25605 15351
rect 25639 15348 25651 15351
rect 27798 15348 27804 15360
rect 25639 15320 27804 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 27798 15308 27804 15320
rect 27856 15308 27862 15360
rect 28166 15308 28172 15360
rect 28224 15348 28230 15360
rect 29733 15351 29791 15357
rect 29733 15348 29745 15351
rect 28224 15320 29745 15348
rect 28224 15308 28230 15320
rect 29733 15317 29745 15320
rect 29779 15317 29791 15351
rect 30466 15348 30472 15360
rect 30427 15320 30472 15348
rect 29733 15311 29791 15317
rect 30466 15308 30472 15320
rect 30524 15308 30530 15360
rect 31110 15308 31116 15360
rect 31168 15348 31174 15360
rect 31757 15351 31815 15357
rect 31757 15348 31769 15351
rect 31168 15320 31769 15348
rect 31168 15308 31174 15320
rect 31757 15317 31769 15320
rect 31803 15317 31815 15351
rect 32398 15348 32404 15360
rect 32359 15320 32404 15348
rect 31757 15311 31815 15317
rect 32398 15308 32404 15320
rect 32456 15308 32462 15360
rect 33796 15348 33824 15379
rect 35529 15351 35587 15357
rect 35529 15348 35541 15351
rect 33796 15320 35541 15348
rect 35529 15317 35541 15320
rect 35575 15317 35587 15351
rect 36096 15348 36124 15388
rect 36354 15376 36360 15388
rect 36412 15376 36418 15428
rect 36449 15419 36507 15425
rect 36449 15385 36461 15419
rect 36495 15385 36507 15419
rect 36449 15379 36507 15385
rect 37553 15419 37611 15425
rect 37553 15385 37565 15419
rect 37599 15385 37611 15419
rect 37553 15379 37611 15385
rect 36464 15348 36492 15379
rect 36096 15320 36492 15348
rect 37568 15348 37596 15379
rect 37642 15376 37648 15428
rect 37700 15416 37706 15428
rect 37700 15388 37745 15416
rect 37700 15376 37706 15388
rect 37734 15348 37740 15360
rect 37568 15320 37740 15348
rect 35529 15311 35587 15317
rect 37734 15308 37740 15320
rect 37792 15308 37798 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 8110 15144 8116 15156
rect 8071 15116 8116 15144
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 13630 15144 13636 15156
rect 13044 15116 13636 15144
rect 13044 15104 13050 15116
rect 13630 15104 13636 15116
rect 13688 15104 13694 15156
rect 16117 15147 16175 15153
rect 16117 15113 16129 15147
rect 16163 15144 16175 15147
rect 17034 15144 17040 15156
rect 16163 15116 17040 15144
rect 16163 15113 16175 15116
rect 16117 15107 16175 15113
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 20165 15147 20223 15153
rect 20165 15144 20177 15147
rect 20036 15116 20177 15144
rect 20036 15104 20042 15116
rect 20165 15113 20177 15116
rect 20211 15113 20223 15147
rect 20165 15107 20223 15113
rect 23106 15104 23112 15156
rect 23164 15144 23170 15156
rect 23382 15144 23388 15156
rect 23164 15116 23388 15144
rect 23164 15104 23170 15116
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 26421 15147 26479 15153
rect 26421 15113 26433 15147
rect 26467 15144 26479 15147
rect 28810 15144 28816 15156
rect 26467 15116 28816 15144
rect 26467 15113 26479 15116
rect 26421 15107 26479 15113
rect 28810 15104 28816 15116
rect 28868 15104 28874 15156
rect 28994 15104 29000 15156
rect 29052 15144 29058 15156
rect 29549 15147 29607 15153
rect 29549 15144 29561 15147
rect 29052 15116 29561 15144
rect 29052 15104 29058 15116
rect 29549 15113 29561 15116
rect 29595 15113 29607 15147
rect 35894 15144 35900 15156
rect 29549 15107 29607 15113
rect 29656 15116 35020 15144
rect 35855 15116 35900 15144
rect 2038 15036 2044 15088
rect 2096 15076 2102 15088
rect 7558 15076 7564 15088
rect 2096 15048 7564 15076
rect 2096 15036 2102 15048
rect 7558 15036 7564 15048
rect 7616 15036 7622 15088
rect 14366 15076 14372 15088
rect 14327 15048 14372 15076
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 14921 15079 14979 15085
rect 14921 15045 14933 15079
rect 14967 15076 14979 15079
rect 15010 15076 15016 15088
rect 14967 15048 15016 15076
rect 14967 15045 14979 15048
rect 14921 15039 14979 15045
rect 15010 15036 15016 15048
rect 15068 15036 15074 15088
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 16942 15076 16948 15088
rect 16724 15048 16948 15076
rect 16724 15036 16730 15048
rect 16942 15036 16948 15048
rect 17000 15036 17006 15088
rect 29656 15076 29684 15116
rect 22066 15048 29684 15076
rect 8018 15008 8024 15020
rect 7979 14980 8024 15008
rect 8018 14968 8024 14980
rect 8076 14968 8082 15020
rect 9766 15008 9772 15020
rect 9727 14980 9772 15008
rect 9766 14968 9772 14980
rect 9824 14968 9830 15020
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 16298 15008 16304 15020
rect 16259 14980 16304 15008
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 17586 14968 17592 15020
rect 17644 15008 17650 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 17644 14980 20085 15008
rect 17644 14968 17650 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20162 14968 20168 15020
rect 20220 15008 20226 15020
rect 22066 15008 22094 15048
rect 30466 15036 30472 15088
rect 30524 15076 30530 15088
rect 30837 15079 30895 15085
rect 30837 15076 30849 15079
rect 30524 15048 30849 15076
rect 30524 15036 30530 15048
rect 30837 15045 30849 15048
rect 30883 15045 30895 15079
rect 30837 15039 30895 15045
rect 32214 15036 32220 15088
rect 32272 15076 32278 15088
rect 32272 15048 32996 15076
rect 32272 15036 32278 15048
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 20220 14980 22201 15008
rect 20220 14968 20226 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 23566 15008 23572 15020
rect 23527 14980 23572 15008
rect 22189 14971 22247 14977
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 25038 15008 25044 15020
rect 24999 14980 25044 15008
rect 25038 14968 25044 14980
rect 25096 14968 25102 15020
rect 26602 15008 26608 15020
rect 26563 14980 26608 15008
rect 26602 14968 26608 14980
rect 26660 14968 26666 15020
rect 26878 14968 26884 15020
rect 26936 15008 26942 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26936 14980 27169 15008
rect 26936 14968 26942 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27249 15011 27307 15017
rect 27249 14977 27261 15011
rect 27295 15008 27307 15011
rect 27522 15008 27528 15020
rect 27295 14980 27528 15008
rect 27295 14977 27307 14980
rect 27249 14971 27307 14977
rect 27522 14968 27528 14980
rect 27580 14968 27586 15020
rect 27706 14968 27712 15020
rect 27764 15008 27770 15020
rect 28997 15011 29055 15017
rect 27764 14980 28948 15008
rect 27764 14968 27770 14980
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14940 14335 14943
rect 15194 14940 15200 14952
rect 14323 14912 15200 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 21542 14900 21548 14952
rect 21600 14940 21606 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 21600 14912 22293 14940
rect 21600 14900 21606 14912
rect 22281 14909 22293 14912
rect 22327 14940 22339 14943
rect 23385 14943 23443 14949
rect 23385 14940 23397 14943
rect 22327 14912 23397 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 23385 14909 23397 14912
rect 23431 14909 23443 14943
rect 23385 14903 23443 14909
rect 28353 14943 28411 14949
rect 28353 14909 28365 14943
rect 28399 14909 28411 14943
rect 28534 14940 28540 14952
rect 28495 14912 28540 14940
rect 28353 14903 28411 14909
rect 17129 14875 17187 14881
rect 17129 14841 17141 14875
rect 17175 14872 17187 14875
rect 26878 14872 26884 14884
rect 17175 14844 26884 14872
rect 17175 14841 17187 14844
rect 17129 14835 17187 14841
rect 26878 14832 26884 14844
rect 26936 14832 26942 14884
rect 28368 14872 28396 14903
rect 28534 14900 28540 14912
rect 28592 14900 28598 14952
rect 28920 14940 28948 14980
rect 28997 14977 29009 15011
rect 29043 15008 29055 15011
rect 29270 15008 29276 15020
rect 29043 14980 29276 15008
rect 29043 14977 29055 14980
rect 28997 14971 29055 14977
rect 29270 14968 29276 14980
rect 29328 14968 29334 15020
rect 29457 15011 29515 15017
rect 29457 14977 29469 15011
rect 29503 15008 29515 15011
rect 30282 15008 30288 15020
rect 29503 14980 30288 15008
rect 29503 14977 29515 14980
rect 29457 14971 29515 14977
rect 30282 14968 30288 14980
rect 30340 14968 30346 15020
rect 32306 15008 32312 15020
rect 32267 14980 32312 15008
rect 32306 14968 32312 14980
rect 32364 14968 32370 15020
rect 32968 15017 32996 15048
rect 34606 15036 34612 15088
rect 34664 15076 34670 15088
rect 34882 15076 34888 15088
rect 34664 15048 34888 15076
rect 34664 15036 34670 15048
rect 34882 15036 34888 15048
rect 34940 15036 34946 15088
rect 34992 15076 35020 15116
rect 35894 15104 35900 15116
rect 35952 15104 35958 15156
rect 38289 15079 38347 15085
rect 38289 15076 38301 15079
rect 34992 15048 38301 15076
rect 38289 15045 38301 15048
rect 38335 15045 38347 15079
rect 38289 15039 38347 15045
rect 32953 15011 33011 15017
rect 32953 14977 32965 15011
rect 32999 14977 33011 15011
rect 32953 14971 33011 14977
rect 34149 15011 34207 15017
rect 34149 14977 34161 15011
rect 34195 15008 34207 15011
rect 35253 15011 35311 15017
rect 35253 15008 35265 15011
rect 34195 14980 35265 15008
rect 34195 14977 34207 14980
rect 34149 14971 34207 14977
rect 35253 14977 35265 14980
rect 35299 14977 35311 15011
rect 36081 15011 36139 15017
rect 36081 15008 36093 15011
rect 35253 14971 35311 14977
rect 35360 14980 36093 15008
rect 30745 14943 30803 14949
rect 30745 14940 30757 14943
rect 28920 14912 30757 14940
rect 30745 14909 30757 14912
rect 30791 14940 30803 14943
rect 30834 14940 30840 14952
rect 30791 14912 30840 14940
rect 30791 14909 30803 14912
rect 30745 14903 30803 14909
rect 30834 14900 30840 14912
rect 30892 14900 30898 14952
rect 31018 14940 31024 14952
rect 30979 14912 31024 14940
rect 31018 14900 31024 14912
rect 31076 14900 31082 14952
rect 33962 14940 33968 14952
rect 31128 14912 33968 14940
rect 28368 14844 29132 14872
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10778 14804 10784 14816
rect 9907 14776 10784 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 24029 14807 24087 14813
rect 24029 14773 24041 14807
rect 24075 14804 24087 14807
rect 24946 14804 24952 14816
rect 24075 14776 24952 14804
rect 24075 14773 24087 14776
rect 24029 14767 24087 14773
rect 24946 14764 24952 14776
rect 25004 14764 25010 14816
rect 25038 14764 25044 14816
rect 25096 14804 25102 14816
rect 25133 14807 25191 14813
rect 25133 14804 25145 14807
rect 25096 14776 25145 14804
rect 25096 14764 25102 14776
rect 25133 14773 25145 14776
rect 25179 14773 25191 14807
rect 29104 14804 29132 14844
rect 30282 14832 30288 14884
rect 30340 14872 30346 14884
rect 31128 14872 31156 14912
rect 33962 14900 33968 14912
rect 34020 14940 34026 14952
rect 34333 14943 34391 14949
rect 34020 14912 34284 14940
rect 34020 14900 34026 14912
rect 33045 14875 33103 14881
rect 33045 14872 33057 14875
rect 30340 14844 31156 14872
rect 31220 14844 33057 14872
rect 30340 14832 30346 14844
rect 29454 14804 29460 14816
rect 29104 14776 29460 14804
rect 25133 14767 25191 14773
rect 29454 14764 29460 14776
rect 29512 14764 29518 14816
rect 30558 14764 30564 14816
rect 30616 14804 30622 14816
rect 31220 14804 31248 14844
rect 33045 14841 33057 14844
rect 33091 14841 33103 14875
rect 34256 14872 34284 14912
rect 34333 14909 34345 14943
rect 34379 14940 34391 14943
rect 34514 14940 34520 14952
rect 34379 14912 34520 14940
rect 34379 14909 34391 14912
rect 34333 14903 34391 14909
rect 34514 14900 34520 14912
rect 34572 14900 34578 14952
rect 35360 14872 35388 14980
rect 36081 14977 36093 14980
rect 36127 14977 36139 15011
rect 36081 14971 36139 14977
rect 36725 15011 36783 15017
rect 36725 14977 36737 15011
rect 36771 15008 36783 15011
rect 36998 15008 37004 15020
rect 36771 14980 37004 15008
rect 36771 14977 36783 14980
rect 36725 14971 36783 14977
rect 36998 14968 37004 14980
rect 37056 14968 37062 15020
rect 38102 15008 38108 15020
rect 38063 14980 38108 15008
rect 38102 14968 38108 14980
rect 38160 14968 38166 15020
rect 36817 14943 36875 14949
rect 36817 14909 36829 14943
rect 36863 14909 36875 14943
rect 36817 14903 36875 14909
rect 34256 14844 35388 14872
rect 33045 14835 33103 14841
rect 35618 14832 35624 14884
rect 35676 14872 35682 14884
rect 36832 14872 36860 14903
rect 35676 14844 36860 14872
rect 35676 14832 35682 14844
rect 30616 14776 31248 14804
rect 30616 14764 30622 14776
rect 31294 14764 31300 14816
rect 31352 14804 31358 14816
rect 32401 14807 32459 14813
rect 32401 14804 32413 14807
rect 31352 14776 32413 14804
rect 31352 14764 31358 14776
rect 32401 14773 32413 14776
rect 32447 14773 32459 14807
rect 32401 14767 32459 14773
rect 33686 14764 33692 14816
rect 33744 14804 33750 14816
rect 34517 14807 34575 14813
rect 34517 14804 34529 14807
rect 33744 14776 34529 14804
rect 33744 14764 33750 14776
rect 34517 14773 34529 14776
rect 34563 14773 34575 14807
rect 34517 14767 34575 14773
rect 34882 14764 34888 14816
rect 34940 14804 34946 14816
rect 35802 14804 35808 14816
rect 34940 14776 35808 14804
rect 34940 14764 34946 14776
rect 35802 14764 35808 14776
rect 35860 14764 35866 14816
rect 35894 14764 35900 14816
rect 35952 14804 35958 14816
rect 36906 14804 36912 14816
rect 35952 14776 36912 14804
rect 35952 14764 35958 14776
rect 36906 14764 36912 14776
rect 36964 14764 36970 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 1854 14600 1860 14612
rect 1627 14572 1860 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 7616 14572 17693 14600
rect 7616 14560 7622 14572
rect 17681 14569 17693 14572
rect 17727 14569 17739 14603
rect 20806 14600 20812 14612
rect 17681 14563 17739 14569
rect 17788 14572 20812 14600
rect 12066 14492 12072 14544
rect 12124 14532 12130 14544
rect 17788 14532 17816 14572
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 20901 14603 20959 14609
rect 20901 14569 20913 14603
rect 20947 14600 20959 14603
rect 22738 14600 22744 14612
rect 20947 14572 22744 14600
rect 20947 14569 20959 14572
rect 20901 14563 20959 14569
rect 22738 14560 22744 14572
rect 22796 14560 22802 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 28442 14600 28448 14612
rect 25188 14572 28448 14600
rect 25188 14560 25194 14572
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 28534 14560 28540 14612
rect 28592 14600 28598 14612
rect 29825 14603 29883 14609
rect 29825 14600 29837 14603
rect 28592 14572 29837 14600
rect 28592 14560 28598 14572
rect 29825 14569 29837 14572
rect 29871 14569 29883 14603
rect 29825 14563 29883 14569
rect 30282 14560 30288 14612
rect 30340 14600 30346 14612
rect 31294 14600 31300 14612
rect 30340 14572 31300 14600
rect 30340 14560 30346 14572
rect 31294 14560 31300 14572
rect 31352 14560 31358 14612
rect 33321 14603 33379 14609
rect 33321 14569 33333 14603
rect 33367 14600 33379 14603
rect 33686 14600 33692 14612
rect 33367 14572 33692 14600
rect 33367 14569 33379 14572
rect 33321 14563 33379 14569
rect 33686 14560 33692 14572
rect 33744 14560 33750 14612
rect 34241 14603 34299 14609
rect 34241 14569 34253 14603
rect 34287 14600 34299 14603
rect 36906 14600 36912 14612
rect 34287 14572 36912 14600
rect 34287 14569 34299 14572
rect 34241 14563 34299 14569
rect 36906 14560 36912 14572
rect 36964 14560 36970 14612
rect 12124 14504 17816 14532
rect 12124 14492 12130 14504
rect 17862 14492 17868 14544
rect 17920 14532 17926 14544
rect 21266 14532 21272 14544
rect 17920 14504 21272 14532
rect 17920 14492 17926 14504
rect 21266 14492 21272 14504
rect 21324 14492 21330 14544
rect 23290 14532 23296 14544
rect 21376 14504 23296 14532
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16942 14464 16948 14476
rect 16071 14436 16948 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17037 14467 17095 14473
rect 17037 14433 17049 14467
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9030 14396 9036 14408
rect 8720 14368 9036 14396
rect 8720 14356 8726 14368
rect 9030 14356 9036 14368
rect 9088 14396 9094 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 9088 14368 9137 14396
rect 9088 14356 9094 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 14918 14396 14924 14408
rect 12299 14368 12434 14396
rect 14879 14368 14924 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 12406 14328 12434 14368
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15194 14396 15200 14408
rect 15059 14368 15200 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 17052 14396 17080 14427
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19484 14436 20668 14464
rect 19484 14424 19490 14436
rect 20640 14405 20668 14436
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 21376 14464 21404 14504
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 26602 14492 26608 14544
rect 26660 14532 26666 14544
rect 29730 14532 29736 14544
rect 26660 14504 29736 14532
rect 26660 14492 26666 14504
rect 29730 14492 29736 14504
rect 29788 14492 29794 14544
rect 30374 14492 30380 14544
rect 30432 14532 30438 14544
rect 31018 14532 31024 14544
rect 30432 14504 31024 14532
rect 30432 14492 30438 14504
rect 31018 14492 31024 14504
rect 31076 14492 31082 14544
rect 34977 14535 35035 14541
rect 31588 14504 32996 14532
rect 21542 14464 21548 14476
rect 20772 14436 21404 14464
rect 21503 14436 21548 14464
rect 20772 14424 20778 14436
rect 21542 14424 21548 14436
rect 21600 14424 21606 14476
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 21876 14436 23060 14464
rect 21876 14424 21882 14436
rect 23032 14405 23060 14436
rect 23106 14424 23112 14476
rect 23164 14464 23170 14476
rect 26694 14464 26700 14476
rect 23164 14436 26700 14464
rect 23164 14424 23170 14436
rect 26694 14424 26700 14436
rect 26752 14424 26758 14476
rect 26878 14424 26884 14476
rect 26936 14464 26942 14476
rect 26936 14436 31524 14464
rect 26936 14424 26942 14436
rect 20625 14399 20683 14405
rect 17052 14368 19564 14396
rect 12406 14300 15240 14328
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 9217 14263 9275 14269
rect 9217 14260 9229 14263
rect 8904 14232 9229 14260
rect 8904 14220 8910 14232
rect 9217 14229 9229 14232
rect 9263 14229 9275 14263
rect 9217 14223 9275 14229
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12345 14263 12403 14269
rect 12345 14260 12357 14263
rect 11940 14232 12357 14260
rect 11940 14220 11946 14232
rect 12345 14229 12357 14232
rect 12391 14229 12403 14263
rect 15212 14260 15240 14300
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 16117 14331 16175 14337
rect 16117 14328 16129 14331
rect 15344 14300 16129 14328
rect 15344 14288 15350 14300
rect 16117 14297 16129 14300
rect 16163 14297 16175 14331
rect 16117 14291 16175 14297
rect 17126 14288 17132 14340
rect 17184 14328 17190 14340
rect 17586 14328 17592 14340
rect 17184 14300 17592 14328
rect 17184 14288 17190 14300
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 16850 14260 16856 14272
rect 15212 14232 16856 14260
rect 12345 14223 12403 14229
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 19536 14260 19564 14368
rect 20625 14365 20637 14399
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14365 23075 14399
rect 23658 14396 23664 14408
rect 23619 14368 23664 14396
rect 23017 14359 23075 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14396 24639 14399
rect 26786 14396 26792 14408
rect 24627 14368 26792 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 26786 14356 26792 14368
rect 26844 14356 26850 14408
rect 28442 14356 28448 14408
rect 28500 14396 28506 14408
rect 28997 14399 29055 14405
rect 28997 14396 29009 14399
rect 28500 14368 29009 14396
rect 28500 14356 28506 14368
rect 28997 14365 29009 14368
rect 29043 14365 29055 14399
rect 29730 14396 29736 14408
rect 29691 14368 29736 14396
rect 28997 14359 29055 14365
rect 29730 14356 29736 14368
rect 29788 14356 29794 14408
rect 21634 14288 21640 14340
rect 21692 14328 21698 14340
rect 21692 14300 21737 14328
rect 21692 14288 21698 14300
rect 21818 14288 21824 14340
rect 21876 14328 21882 14340
rect 22370 14328 22376 14340
rect 21876 14300 22376 14328
rect 21876 14288 21882 14300
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 22557 14331 22615 14337
rect 22557 14297 22569 14331
rect 22603 14328 22615 14331
rect 22830 14328 22836 14340
rect 22603 14300 22836 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 22830 14288 22836 14300
rect 22888 14288 22894 14340
rect 24854 14288 24860 14340
rect 24912 14328 24918 14340
rect 27525 14331 27583 14337
rect 27525 14328 27537 14331
rect 24912 14300 27537 14328
rect 24912 14288 24918 14300
rect 27525 14297 27537 14300
rect 27571 14297 27583 14331
rect 27525 14291 27583 14297
rect 27614 14288 27620 14340
rect 27672 14328 27678 14340
rect 28534 14328 28540 14340
rect 27672 14300 27717 14328
rect 28495 14300 28540 14328
rect 27672 14288 27678 14300
rect 28534 14288 28540 14300
rect 28592 14288 28598 14340
rect 30466 14328 30472 14340
rect 28644 14300 30472 14328
rect 22922 14260 22928 14272
rect 19536 14232 22928 14260
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 23106 14260 23112 14272
rect 23067 14232 23112 14260
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 23566 14220 23572 14272
rect 23624 14260 23630 14272
rect 23753 14263 23811 14269
rect 23753 14260 23765 14263
rect 23624 14232 23765 14260
rect 23624 14220 23630 14232
rect 23753 14229 23765 14232
rect 23799 14229 23811 14263
rect 23753 14223 23811 14229
rect 24673 14263 24731 14269
rect 24673 14229 24685 14263
rect 24719 14260 24731 14263
rect 24762 14260 24768 14272
rect 24719 14232 24768 14260
rect 24719 14229 24731 14232
rect 24673 14223 24731 14229
rect 24762 14220 24768 14232
rect 24820 14220 24826 14272
rect 24946 14220 24952 14272
rect 25004 14260 25010 14272
rect 28644 14260 28672 14300
rect 30466 14288 30472 14300
rect 30524 14288 30530 14340
rect 30558 14288 30564 14340
rect 30616 14328 30622 14340
rect 31113 14331 31171 14337
rect 31113 14328 31125 14331
rect 30616 14300 30661 14328
rect 30760 14300 31125 14328
rect 30616 14288 30622 14300
rect 25004 14232 28672 14260
rect 29089 14263 29147 14269
rect 25004 14220 25010 14232
rect 29089 14229 29101 14263
rect 29135 14260 29147 14263
rect 29454 14260 29460 14272
rect 29135 14232 29460 14260
rect 29135 14229 29147 14232
rect 29089 14223 29147 14229
rect 29454 14220 29460 14232
rect 29512 14220 29518 14272
rect 30006 14220 30012 14272
rect 30064 14260 30070 14272
rect 30760 14260 30788 14300
rect 31113 14297 31125 14300
rect 31159 14297 31171 14331
rect 31496 14328 31524 14436
rect 31588 14405 31616 14504
rect 32398 14424 32404 14476
rect 32456 14464 32462 14476
rect 32861 14467 32919 14473
rect 32861 14464 32873 14467
rect 32456 14436 32873 14464
rect 32456 14424 32462 14436
rect 32861 14433 32873 14436
rect 32907 14433 32919 14467
rect 32968 14464 32996 14504
rect 34977 14501 34989 14535
rect 35023 14532 35035 14535
rect 37642 14532 37648 14544
rect 35023 14504 37648 14532
rect 35023 14501 35035 14504
rect 34977 14495 35035 14501
rect 37642 14492 37648 14504
rect 37700 14492 37706 14544
rect 32968 14436 35020 14464
rect 32861 14427 32919 14433
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14365 31631 14399
rect 31573 14359 31631 14365
rect 32677 14399 32735 14405
rect 32677 14365 32689 14399
rect 32723 14365 32735 14399
rect 34146 14396 34152 14408
rect 34107 14368 34152 14396
rect 32677 14359 32735 14365
rect 32692 14328 32720 14359
rect 34146 14356 34152 14368
rect 34204 14356 34210 14408
rect 34238 14356 34244 14408
rect 34296 14396 34302 14408
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34296 14368 34897 14396
rect 34296 14356 34302 14368
rect 34885 14365 34897 14368
rect 34931 14365 34943 14399
rect 34992 14396 35020 14436
rect 35342 14424 35348 14476
rect 35400 14464 35406 14476
rect 36541 14467 36599 14473
rect 36541 14464 36553 14467
rect 35400 14436 36553 14464
rect 35400 14424 35406 14436
rect 36541 14433 36553 14436
rect 36587 14433 36599 14467
rect 36541 14427 36599 14433
rect 36722 14424 36728 14476
rect 36780 14464 36786 14476
rect 37461 14467 37519 14473
rect 37461 14464 37473 14467
rect 36780 14436 37473 14464
rect 36780 14424 36786 14436
rect 37461 14433 37473 14436
rect 37507 14433 37519 14467
rect 37461 14427 37519 14433
rect 35894 14396 35900 14408
rect 34992 14368 35900 14396
rect 34885 14359 34943 14365
rect 35894 14356 35900 14368
rect 35952 14356 35958 14408
rect 36446 14396 36452 14408
rect 36407 14368 36452 14396
rect 36446 14356 36452 14368
rect 36504 14356 36510 14408
rect 35618 14328 35624 14340
rect 31496 14300 31800 14328
rect 32692 14300 35624 14328
rect 31113 14291 31171 14297
rect 30064 14232 30788 14260
rect 30064 14220 30070 14232
rect 30834 14220 30840 14272
rect 30892 14260 30898 14272
rect 31665 14263 31723 14269
rect 31665 14260 31677 14263
rect 30892 14232 31677 14260
rect 30892 14220 30898 14232
rect 31665 14229 31677 14232
rect 31711 14229 31723 14263
rect 31772 14260 31800 14300
rect 35618 14288 35624 14300
rect 35676 14288 35682 14340
rect 35805 14331 35863 14337
rect 35805 14297 35817 14331
rect 35851 14328 35863 14331
rect 37185 14331 37243 14337
rect 37185 14328 37197 14331
rect 35851 14300 37197 14328
rect 35851 14297 35863 14300
rect 35805 14291 35863 14297
rect 37185 14297 37197 14300
rect 37231 14297 37243 14331
rect 37185 14291 37243 14297
rect 37274 14288 37280 14340
rect 37332 14328 37338 14340
rect 37332 14300 37377 14328
rect 37332 14288 37338 14300
rect 38010 14260 38016 14272
rect 31772 14232 38016 14260
rect 31665 14223 31723 14229
rect 38010 14220 38016 14232
rect 38068 14220 38074 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9214 14016 9220 14068
rect 9272 14056 9278 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 9272 14028 9321 14056
rect 9272 14016 9278 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 9309 14019 9367 14025
rect 14921 14059 14979 14065
rect 14921 14025 14933 14059
rect 14967 14056 14979 14059
rect 23014 14056 23020 14068
rect 14967 14028 18828 14056
rect 14967 14025 14979 14028
rect 14921 14019 14979 14025
rect 11882 13988 11888 14000
rect 11843 13960 11888 13988
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 17862 13988 17868 14000
rect 17823 13960 17868 13988
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 11054 13920 11060 13932
rect 10560 13892 11060 13920
rect 10560 13880 10566 13892
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13688 13892 14289 13920
rect 13688 13880 13694 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 10318 13852 10324 13864
rect 8711 13824 10324 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 10836 13824 11805 13852
rect 10836 13812 10842 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 12066 13852 12072 13864
rect 12027 13824 12072 13852
rect 11793 13815 11851 13821
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 14458 13852 14464 13864
rect 14419 13824 14464 13852
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 17770 13852 17776 13864
rect 17731 13824 17776 13852
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 18414 13852 18420 13864
rect 18375 13824 18420 13852
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 18800 13852 18828 14028
rect 18892 14028 23020 14056
rect 18892 13929 18920 14028
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 30190 14056 30196 14068
rect 30151 14028 30196 14056
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 32401 14059 32459 14065
rect 32401 14056 32413 14059
rect 31726 14028 32413 14056
rect 20625 13991 20683 13997
rect 20625 13957 20637 13991
rect 20671 13988 20683 13991
rect 21174 13988 21180 14000
rect 20671 13960 21180 13988
rect 20671 13957 20683 13960
rect 20625 13951 20683 13957
rect 21174 13948 21180 13960
rect 21232 13948 21238 14000
rect 22186 13988 22192 14000
rect 22147 13960 22192 13988
rect 22186 13948 22192 13960
rect 22244 13948 22250 14000
rect 22922 13948 22928 14000
rect 22980 13988 22986 14000
rect 24762 13988 24768 14000
rect 22980 13960 24532 13988
rect 24723 13960 24768 13988
rect 22980 13948 22986 13960
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13889 18935 13923
rect 21818 13920 21824 13932
rect 18877 13883 18935 13889
rect 19812 13892 21824 13920
rect 19812 13852 19840 13892
rect 21818 13880 21824 13892
rect 21876 13880 21882 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23569 13923 23627 13929
rect 23569 13920 23581 13923
rect 23532 13892 23581 13920
rect 23532 13880 23538 13892
rect 23569 13889 23581 13892
rect 23615 13889 23627 13923
rect 23569 13883 23627 13889
rect 19978 13852 19984 13864
rect 18800 13824 19840 13852
rect 19939 13824 19984 13852
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 20162 13852 20168 13864
rect 20123 13824 20168 13852
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 21315 13824 22109 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 23290 13852 23296 13864
rect 23155 13824 23296 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 15838 13744 15844 13796
rect 15896 13784 15902 13796
rect 21910 13784 21916 13796
rect 15896 13756 21916 13784
rect 15896 13744 15902 13756
rect 21910 13744 21916 13756
rect 21968 13744 21974 13796
rect 24504 13784 24532 13960
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 28261 13991 28319 13997
rect 28261 13988 28273 13991
rect 27856 13960 28273 13988
rect 27856 13948 27862 13960
rect 28261 13957 28273 13960
rect 28307 13957 28319 13991
rect 28261 13951 28319 13957
rect 28813 13991 28871 13997
rect 28813 13957 28825 13991
rect 28859 13988 28871 13991
rect 30006 13988 30012 14000
rect 28859 13960 30012 13988
rect 28859 13957 28871 13960
rect 28813 13951 28871 13957
rect 30006 13948 30012 13960
rect 30064 13988 30070 14000
rect 30558 13988 30564 14000
rect 30064 13960 30564 13988
rect 30064 13948 30070 13960
rect 30558 13948 30564 13960
rect 30616 13948 30622 14000
rect 29086 13880 29092 13932
rect 29144 13920 29150 13932
rect 29457 13923 29515 13929
rect 29457 13920 29469 13923
rect 29144 13892 29469 13920
rect 29144 13880 29150 13892
rect 29457 13889 29469 13892
rect 29503 13889 29515 13923
rect 30098 13920 30104 13932
rect 30059 13892 30104 13920
rect 29457 13883 29515 13889
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 31205 13923 31263 13929
rect 31205 13889 31217 13923
rect 31251 13920 31263 13923
rect 31726 13920 31754 14028
rect 32401 14025 32413 14028
rect 32447 14025 32459 14059
rect 32401 14019 32459 14025
rect 33781 14059 33839 14065
rect 33781 14025 33793 14059
rect 33827 14025 33839 14059
rect 34514 14056 34520 14068
rect 34475 14028 34520 14056
rect 33781 14019 33839 14025
rect 33796 13988 33824 14019
rect 34514 14016 34520 14028
rect 34572 14016 34578 14068
rect 35802 13988 35808 14000
rect 33796 13960 34744 13988
rect 35763 13960 35808 13988
rect 32582 13920 32588 13932
rect 31251 13892 31754 13920
rect 32543 13892 32588 13920
rect 31251 13889 31263 13892
rect 31205 13883 31263 13889
rect 32582 13880 32588 13892
rect 32640 13880 32646 13932
rect 32766 13880 32772 13932
rect 32824 13920 32830 13932
rect 34716 13929 34744 13960
rect 35802 13948 35808 13960
rect 35860 13948 35866 14000
rect 33965 13923 34023 13929
rect 33965 13920 33977 13923
rect 32824 13892 33977 13920
rect 32824 13880 32830 13892
rect 33965 13889 33977 13892
rect 34011 13889 34023 13923
rect 33965 13883 34023 13889
rect 34701 13923 34759 13929
rect 34701 13889 34713 13923
rect 34747 13889 34759 13923
rect 34701 13883 34759 13889
rect 36354 13880 36360 13932
rect 36412 13920 36418 13932
rect 38013 13923 38071 13929
rect 38013 13920 38025 13923
rect 36412 13892 38025 13920
rect 36412 13880 36418 13892
rect 38013 13889 38025 13892
rect 38059 13889 38071 13923
rect 38013 13883 38071 13889
rect 24670 13852 24676 13864
rect 24631 13824 24676 13852
rect 24670 13812 24676 13824
rect 24728 13812 24734 13864
rect 24949 13855 25007 13861
rect 24949 13852 24961 13855
rect 24780 13824 24961 13852
rect 24780 13784 24808 13824
rect 24949 13821 24961 13824
rect 24995 13852 25007 13855
rect 24995 13824 27568 13852
rect 24995 13821 25007 13824
rect 24949 13815 25007 13821
rect 24504 13756 24808 13784
rect 27540 13784 27568 13824
rect 27614 13812 27620 13864
rect 27672 13852 27678 13864
rect 28169 13855 28227 13861
rect 28169 13852 28181 13855
rect 27672 13824 28181 13852
rect 27672 13812 27678 13824
rect 28169 13821 28181 13824
rect 28215 13821 28227 13855
rect 30374 13852 30380 13864
rect 28169 13815 28227 13821
rect 28276 13824 30380 13852
rect 28276 13784 28304 13824
rect 30374 13812 30380 13824
rect 30432 13812 30438 13864
rect 31018 13852 31024 13864
rect 30979 13824 31024 13852
rect 31018 13812 31024 13824
rect 31076 13812 31082 13864
rect 35710 13852 35716 13864
rect 35671 13824 35716 13852
rect 35710 13812 35716 13824
rect 35768 13812 35774 13864
rect 35894 13812 35900 13864
rect 35952 13852 35958 13864
rect 35989 13855 36047 13861
rect 35989 13852 36001 13855
rect 35952 13824 36001 13852
rect 35952 13812 35958 13824
rect 35989 13821 36001 13824
rect 36035 13821 36047 13855
rect 35989 13815 36047 13821
rect 27540 13756 28304 13784
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 18966 13716 18972 13728
rect 18927 13688 18972 13716
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 21174 13676 21180 13728
rect 21232 13716 21238 13728
rect 26326 13716 26332 13728
rect 21232 13688 26332 13716
rect 21232 13676 21238 13688
rect 26326 13676 26332 13688
rect 26384 13676 26390 13728
rect 29270 13716 29276 13728
rect 29231 13688 29276 13716
rect 29270 13676 29276 13688
rect 29328 13676 29334 13728
rect 31294 13676 31300 13728
rect 31352 13716 31358 13728
rect 31389 13719 31447 13725
rect 31389 13716 31401 13719
rect 31352 13688 31401 13716
rect 31352 13676 31358 13688
rect 31389 13685 31401 13688
rect 31435 13685 31447 13719
rect 38194 13716 38200 13728
rect 38155 13688 38200 13716
rect 31389 13679 31447 13685
rect 38194 13676 38200 13688
rect 38252 13676 38258 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14516 13484 14749 13512
rect 14516 13472 14522 13484
rect 14737 13481 14749 13484
rect 14783 13481 14795 13515
rect 14737 13475 14795 13481
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 28258 13512 28264 13524
rect 21140 13484 28264 13512
rect 21140 13472 21146 13484
rect 28258 13472 28264 13484
rect 28316 13472 28322 13524
rect 28442 13472 28448 13524
rect 28500 13512 28506 13524
rect 28626 13512 28632 13524
rect 28500 13484 28632 13512
rect 28500 13472 28506 13484
rect 28626 13472 28632 13484
rect 28684 13512 28690 13524
rect 30377 13515 30435 13521
rect 28684 13484 29040 13512
rect 28684 13472 28690 13484
rect 18598 13444 18604 13456
rect 12406 13416 18604 13444
rect 10778 13376 10784 13388
rect 10739 13348 10784 13376
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 11054 13376 11060 13388
rect 11015 13348 11060 13376
rect 11054 13336 11060 13348
rect 11112 13376 11118 13388
rect 12406 13376 12434 13416
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 23293 13447 23351 13453
rect 23293 13413 23305 13447
rect 23339 13413 23351 13447
rect 23293 13407 23351 13413
rect 24581 13447 24639 13453
rect 24581 13413 24593 13447
rect 24627 13444 24639 13447
rect 24627 13416 26556 13444
rect 24627 13413 24639 13416
rect 24581 13407 24639 13413
rect 16942 13376 16948 13388
rect 11112 13348 12434 13376
rect 16903 13348 16948 13376
rect 11112 13336 11118 13348
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17218 13376 17224 13388
rect 17179 13348 17224 13376
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 19978 13376 19984 13388
rect 19939 13348 19984 13376
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 23308 13376 23336 13407
rect 26326 13376 26332 13388
rect 23308 13348 24808 13376
rect 26287 13348 26332 13376
rect 14826 13268 14832 13320
rect 14884 13308 14890 13320
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14884 13280 14933 13308
rect 14884 13268 14890 13280
rect 14921 13277 14933 13280
rect 14967 13277 14979 13311
rect 14921 13271 14979 13277
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 22094 13308 22100 13320
rect 21591 13280 22100 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 24780 13317 24808 13348
rect 26326 13336 26332 13348
rect 26384 13336 26390 13388
rect 26528 13385 26556 13416
rect 26694 13404 26700 13456
rect 26752 13444 26758 13456
rect 28905 13447 28963 13453
rect 28905 13444 28917 13447
rect 26752 13416 28917 13444
rect 26752 13404 26758 13416
rect 28905 13413 28917 13416
rect 28951 13413 28963 13447
rect 29012 13444 29040 13484
rect 30377 13481 30389 13515
rect 30423 13512 30435 13515
rect 30466 13512 30472 13524
rect 30423 13484 30472 13512
rect 30423 13481 30435 13484
rect 30377 13475 30435 13481
rect 30466 13472 30472 13484
rect 30524 13472 30530 13524
rect 34149 13515 34207 13521
rect 34149 13481 34161 13515
rect 34195 13512 34207 13515
rect 35802 13512 35808 13524
rect 34195 13484 35808 13512
rect 34195 13481 34207 13484
rect 34149 13475 34207 13481
rect 35802 13472 35808 13484
rect 35860 13472 35866 13524
rect 38197 13515 38255 13521
rect 38197 13481 38209 13515
rect 38243 13512 38255 13515
rect 38654 13512 38660 13524
rect 38243 13484 38660 13512
rect 38243 13481 38255 13484
rect 38197 13475 38255 13481
rect 38654 13472 38660 13484
rect 38712 13472 38718 13524
rect 37550 13444 37556 13456
rect 29012 13416 31340 13444
rect 37511 13416 37556 13444
rect 28905 13407 28963 13413
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13345 26571 13379
rect 26513 13339 26571 13345
rect 28721 13379 28779 13385
rect 28721 13345 28733 13379
rect 28767 13376 28779 13379
rect 29270 13376 29276 13388
rect 28767 13348 29276 13376
rect 28767 13345 28779 13348
rect 28721 13339 28779 13345
rect 29270 13336 29276 13348
rect 29328 13336 29334 13388
rect 29454 13336 29460 13388
rect 29512 13376 29518 13388
rect 29917 13379 29975 13385
rect 29917 13376 29929 13379
rect 29512 13348 29929 13376
rect 29512 13336 29518 13348
rect 29917 13345 29929 13348
rect 29963 13345 29975 13379
rect 31202 13376 31208 13388
rect 31163 13348 31208 13376
rect 29917 13339 29975 13345
rect 31202 13336 31208 13348
rect 31260 13336 31266 13388
rect 22649 13311 22707 13317
rect 22649 13277 22661 13311
rect 22695 13277 22707 13311
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 22649 13271 22707 13277
rect 23308 13280 23489 13308
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 10928 13212 10973 13240
rect 10928 13200 10934 13212
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17092 13212 17137 13240
rect 17092 13200 17098 13212
rect 18138 13200 18144 13252
rect 18196 13240 18202 13252
rect 22664 13240 22692 13271
rect 18196 13212 22692 13240
rect 18196 13200 18202 13212
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 18156 13172 18184 13200
rect 21634 13172 21640 13184
rect 13136 13144 18184 13172
rect 21595 13144 21640 13172
rect 13136 13132 13142 13144
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 22738 13172 22744 13184
rect 22699 13144 22744 13172
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 23308 13172 23336 13280
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 27154 13308 27160 13320
rect 24765 13271 24823 13277
rect 26712 13280 27160 13308
rect 26712 13172 26740 13280
rect 27154 13268 27160 13280
rect 27212 13308 27218 13320
rect 27893 13311 27951 13317
rect 27893 13308 27905 13311
rect 27212 13280 27905 13308
rect 27212 13268 27218 13280
rect 27893 13277 27905 13280
rect 27939 13277 27951 13311
rect 27893 13271 27951 13277
rect 28537 13311 28595 13317
rect 28537 13277 28549 13311
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13308 29791 13311
rect 31018 13308 31024 13320
rect 29779 13280 31024 13308
rect 29779 13277 29791 13280
rect 29733 13271 29791 13277
rect 28552 13240 28580 13271
rect 31018 13268 31024 13280
rect 31076 13268 31082 13320
rect 31312 13308 31340 13416
rect 37550 13404 37556 13416
rect 37608 13404 37614 13456
rect 31389 13379 31447 13385
rect 31389 13345 31401 13379
rect 31435 13376 31447 13379
rect 32401 13379 32459 13385
rect 32401 13376 32413 13379
rect 31435 13348 32413 13376
rect 31435 13345 31447 13348
rect 31389 13339 31447 13345
rect 32401 13345 32413 13348
rect 32447 13345 32459 13379
rect 32401 13339 32459 13345
rect 35342 13336 35348 13388
rect 35400 13376 35406 13388
rect 35400 13348 38148 13376
rect 35400 13336 35406 13348
rect 32306 13308 32312 13320
rect 31312 13280 32312 13308
rect 32306 13268 32312 13280
rect 32364 13268 32370 13320
rect 32950 13308 32956 13320
rect 32911 13280 32956 13308
rect 32950 13268 32956 13280
rect 33008 13268 33014 13320
rect 33318 13268 33324 13320
rect 33376 13308 33382 13320
rect 34057 13311 34115 13317
rect 34057 13308 34069 13311
rect 33376 13280 34069 13308
rect 33376 13268 33382 13280
rect 34057 13277 34069 13280
rect 34103 13277 34115 13311
rect 34057 13271 34115 13277
rect 34514 13268 34520 13320
rect 34572 13308 34578 13320
rect 38120 13317 38148 13348
rect 35069 13311 35127 13317
rect 35069 13308 35081 13311
rect 34572 13280 35081 13308
rect 34572 13268 34578 13280
rect 35069 13277 35081 13280
rect 35115 13277 35127 13311
rect 35069 13271 35127 13277
rect 38105 13311 38163 13317
rect 38105 13277 38117 13311
rect 38151 13277 38163 13311
rect 38105 13271 38163 13277
rect 30466 13240 30472 13252
rect 28552 13212 30472 13240
rect 30466 13200 30472 13212
rect 30524 13200 30530 13252
rect 33045 13243 33103 13249
rect 33045 13209 33057 13243
rect 33091 13240 33103 13243
rect 34790 13240 34796 13252
rect 33091 13212 34796 13240
rect 33091 13209 33103 13212
rect 33045 13203 33103 13209
rect 34790 13200 34796 13212
rect 34848 13200 34854 13252
rect 35618 13200 35624 13252
rect 35676 13240 35682 13252
rect 36998 13240 37004 13252
rect 35676 13212 37004 13240
rect 35676 13200 35682 13212
rect 36998 13200 37004 13212
rect 37056 13200 37062 13252
rect 37090 13200 37096 13252
rect 37148 13240 37154 13252
rect 37148 13212 37193 13240
rect 37148 13200 37154 13212
rect 26970 13172 26976 13184
rect 23308 13144 26740 13172
rect 26931 13144 26976 13172
rect 26970 13132 26976 13144
rect 27028 13132 27034 13184
rect 27985 13175 28043 13181
rect 27985 13141 27997 13175
rect 28031 13172 28043 13175
rect 28994 13172 29000 13184
rect 28031 13144 29000 13172
rect 28031 13141 28043 13144
rect 27985 13135 28043 13141
rect 28994 13132 29000 13144
rect 29052 13132 29058 13184
rect 31294 13132 31300 13184
rect 31352 13172 31358 13184
rect 31849 13175 31907 13181
rect 31849 13172 31861 13175
rect 31352 13144 31861 13172
rect 31352 13132 31358 13144
rect 31849 13141 31861 13144
rect 31895 13141 31907 13175
rect 34882 13172 34888 13184
rect 34843 13144 34888 13172
rect 31849 13135 31907 13141
rect 34882 13132 34888 13144
rect 34940 13132 34946 13184
rect 35526 13172 35532 13184
rect 35487 13144 35532 13172
rect 35526 13132 35532 13144
rect 35584 13132 35590 13184
rect 36170 13172 36176 13184
rect 36131 13144 36176 13172
rect 36170 13132 36176 13144
rect 36228 13132 36234 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 28077 12971 28135 12977
rect 1636 12940 26832 12968
rect 1636 12928 1642 12940
rect 5442 12900 5448 12912
rect 1596 12872 5448 12900
rect 1596 12841 1624 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 10597 12903 10655 12909
rect 10597 12869 10609 12903
rect 10643 12900 10655 12903
rect 10870 12900 10876 12912
rect 10643 12872 10876 12900
rect 10643 12869 10655 12872
rect 10597 12863 10655 12869
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 12250 12900 12256 12912
rect 12211 12872 12256 12900
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 18325 12903 18383 12909
rect 18325 12869 18337 12903
rect 18371 12900 18383 12903
rect 18966 12900 18972 12912
rect 18371 12872 18972 12900
rect 18371 12869 18383 12872
rect 18325 12863 18383 12869
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 22738 12860 22744 12912
rect 22796 12900 22802 12912
rect 23661 12903 23719 12909
rect 23661 12900 23673 12903
rect 22796 12872 23673 12900
rect 22796 12860 22802 12872
rect 23661 12869 23673 12872
rect 23707 12869 23719 12903
rect 23661 12863 23719 12869
rect 24213 12903 24271 12909
rect 24213 12869 24225 12903
rect 24259 12900 24271 12903
rect 24762 12900 24768 12912
rect 24259 12872 24768 12900
rect 24259 12869 24271 12872
rect 24213 12863 24271 12869
rect 24762 12860 24768 12872
rect 24820 12860 24826 12912
rect 25038 12900 25044 12912
rect 24999 12872 25044 12900
rect 25038 12860 25044 12872
rect 25096 12860 25102 12912
rect 26804 12900 26832 12940
rect 28077 12937 28089 12971
rect 28123 12968 28135 12971
rect 29086 12968 29092 12980
rect 28123 12940 29092 12968
rect 28123 12937 28135 12940
rect 28077 12931 28135 12937
rect 29086 12928 29092 12940
rect 29144 12928 29150 12980
rect 32582 12968 32588 12980
rect 32543 12940 32588 12968
rect 32582 12928 32588 12940
rect 32640 12928 32646 12980
rect 33321 12971 33379 12977
rect 33321 12937 33333 12971
rect 33367 12968 33379 12971
rect 33367 12940 36308 12968
rect 33367 12937 33379 12940
rect 33321 12931 33379 12937
rect 31573 12903 31631 12909
rect 31573 12900 31585 12903
rect 26804 12872 31585 12900
rect 31573 12869 31585 12872
rect 31619 12869 31631 12903
rect 31573 12863 31631 12869
rect 32122 12860 32128 12912
rect 32180 12900 32186 12912
rect 34882 12900 34888 12912
rect 32180 12872 34100 12900
rect 34843 12872 34888 12900
rect 32180 12860 32186 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12832 4307 12835
rect 4706 12832 4712 12844
rect 4295 12804 4712 12832
rect 4295 12801 4307 12804
rect 4249 12795 4307 12801
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 12158 12832 12164 12844
rect 12119 12804 12164 12832
rect 10505 12795 10563 12801
rect 10520 12764 10548 12795
rect 12158 12792 12164 12804
rect 12216 12792 12222 12844
rect 15013 12835 15071 12841
rect 15013 12801 15025 12835
rect 15059 12832 15071 12835
rect 15838 12832 15844 12844
rect 15059 12804 15844 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 19886 12832 19892 12844
rect 19847 12804 19892 12832
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 23106 12832 23112 12844
rect 22235 12804 23112 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 23106 12792 23112 12804
rect 23164 12792 23170 12844
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12832 25651 12835
rect 27614 12832 27620 12844
rect 25639 12804 27620 12832
rect 25639 12801 25651 12804
rect 25593 12795 25651 12801
rect 13078 12764 13084 12776
rect 10520 12736 13084 12764
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 17460 12736 18245 12764
rect 17460 12724 17466 12736
rect 18233 12733 18245 12736
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18414 12724 18420 12776
rect 18472 12764 18478 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18472 12736 18889 12764
rect 18472 12724 18478 12736
rect 18877 12733 18889 12736
rect 18923 12764 18935 12767
rect 22005 12767 22063 12773
rect 18923 12736 20300 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 14826 12696 14832 12708
rect 14787 12668 14832 12696
rect 14826 12656 14832 12668
rect 14884 12656 14890 12708
rect 19705 12699 19763 12705
rect 19705 12665 19717 12699
rect 19751 12696 19763 12699
rect 20162 12696 20168 12708
rect 19751 12668 20168 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 20162 12656 20168 12668
rect 20220 12656 20226 12708
rect 20272 12696 20300 12736
rect 22005 12733 22017 12767
rect 22051 12764 22063 12767
rect 23566 12764 23572 12776
rect 22051 12736 23572 12764
rect 22051 12733 22063 12736
rect 22005 12727 22063 12733
rect 23566 12724 23572 12736
rect 23624 12724 23630 12776
rect 24670 12724 24676 12776
rect 24728 12764 24734 12776
rect 24949 12767 25007 12773
rect 24949 12764 24961 12767
rect 24728 12736 24961 12764
rect 24728 12724 24734 12736
rect 24949 12733 24961 12736
rect 24995 12733 25007 12767
rect 24949 12727 25007 12733
rect 22370 12696 22376 12708
rect 20272 12668 22094 12696
rect 22331 12668 22376 12696
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 4062 12628 4068 12640
rect 4023 12600 4068 12628
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 22066 12628 22094 12668
rect 22370 12656 22376 12668
rect 22428 12656 22434 12708
rect 25608 12628 25636 12795
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 28258 12832 28264 12844
rect 28219 12804 28264 12832
rect 28258 12792 28264 12804
rect 28316 12792 28322 12844
rect 28994 12792 29000 12844
rect 29052 12832 29058 12844
rect 29273 12835 29331 12841
rect 29273 12832 29285 12835
rect 29052 12804 29285 12832
rect 29052 12792 29058 12804
rect 29273 12801 29285 12804
rect 29319 12801 29331 12835
rect 31294 12832 31300 12844
rect 29273 12795 29331 12801
rect 30116 12804 31300 12832
rect 29089 12767 29147 12773
rect 29089 12733 29101 12767
rect 29135 12764 29147 12767
rect 30116 12764 30144 12804
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 31389 12835 31447 12841
rect 31389 12801 31401 12835
rect 31435 12832 31447 12835
rect 31478 12832 31484 12844
rect 31435 12804 31484 12832
rect 31435 12801 31447 12804
rect 31389 12795 31447 12801
rect 29135 12736 30144 12764
rect 30193 12767 30251 12773
rect 29135 12733 29147 12736
rect 29089 12727 29147 12733
rect 30193 12733 30205 12767
rect 30239 12733 30251 12767
rect 30374 12764 30380 12776
rect 30335 12736 30380 12764
rect 30193 12727 30251 12733
rect 29178 12656 29184 12708
rect 29236 12696 29242 12708
rect 30208 12696 30236 12727
rect 30374 12724 30380 12736
rect 30432 12724 30438 12776
rect 31202 12724 31208 12776
rect 31260 12764 31266 12776
rect 31404 12764 31432 12795
rect 31478 12792 31484 12804
rect 31536 12792 31542 12844
rect 32306 12792 32312 12844
rect 32364 12832 32370 12844
rect 32769 12835 32827 12841
rect 32769 12832 32781 12835
rect 32364 12804 32781 12832
rect 32364 12792 32370 12804
rect 32769 12801 32781 12804
rect 32815 12801 32827 12835
rect 32769 12795 32827 12801
rect 33229 12835 33287 12841
rect 33229 12801 33241 12835
rect 33275 12832 33287 12835
rect 33594 12832 33600 12844
rect 33275 12804 33600 12832
rect 33275 12801 33287 12804
rect 33229 12795 33287 12801
rect 33594 12792 33600 12804
rect 33652 12792 33658 12844
rect 34072 12841 34100 12872
rect 34882 12860 34888 12872
rect 34940 12860 34946 12912
rect 34974 12860 34980 12912
rect 35032 12900 35038 12912
rect 35618 12900 35624 12912
rect 35032 12872 35624 12900
rect 35032 12860 35038 12872
rect 35618 12860 35624 12872
rect 35676 12860 35682 12912
rect 36170 12900 36176 12912
rect 36131 12872 36176 12900
rect 36170 12860 36176 12872
rect 36228 12860 36234 12912
rect 36280 12909 36308 12940
rect 36265 12903 36323 12909
rect 36265 12869 36277 12903
rect 36311 12869 36323 12903
rect 36265 12863 36323 12869
rect 34057 12835 34115 12841
rect 34057 12801 34069 12835
rect 34103 12801 34115 12835
rect 34057 12795 34115 12801
rect 31260 12736 31432 12764
rect 31260 12724 31266 12736
rect 29236 12668 30236 12696
rect 30837 12699 30895 12705
rect 29236 12656 29242 12668
rect 30837 12665 30849 12699
rect 30883 12696 30895 12699
rect 34072 12696 34100 12795
rect 37366 12792 37372 12844
rect 37424 12832 37430 12844
rect 38013 12835 38071 12841
rect 38013 12832 38025 12835
rect 37424 12804 38025 12832
rect 37424 12792 37430 12804
rect 38013 12801 38025 12804
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 34793 12767 34851 12773
rect 34793 12733 34805 12767
rect 34839 12764 34851 12767
rect 35526 12764 35532 12776
rect 34839 12736 35532 12764
rect 34839 12733 34851 12736
rect 34793 12727 34851 12733
rect 35526 12724 35532 12736
rect 35584 12724 35590 12776
rect 35802 12724 35808 12776
rect 35860 12764 35866 12776
rect 36449 12767 36507 12773
rect 36449 12764 36461 12767
rect 35860 12736 36461 12764
rect 35860 12724 35866 12736
rect 36449 12733 36461 12736
rect 36495 12733 36507 12767
rect 36449 12727 36507 12733
rect 35345 12699 35403 12705
rect 35345 12696 35357 12699
rect 30883 12668 31754 12696
rect 34072 12668 35357 12696
rect 30883 12665 30895 12668
rect 30837 12659 30895 12665
rect 22066 12600 25636 12628
rect 26970 12588 26976 12640
rect 27028 12628 27034 12640
rect 29457 12631 29515 12637
rect 29457 12628 29469 12631
rect 27028 12600 29469 12628
rect 27028 12588 27034 12600
rect 29457 12597 29469 12600
rect 29503 12628 29515 12631
rect 31570 12628 31576 12640
rect 29503 12600 31576 12628
rect 29503 12597 29515 12600
rect 29457 12591 29515 12597
rect 31570 12588 31576 12600
rect 31628 12588 31634 12640
rect 31726 12628 31754 12668
rect 35345 12665 35357 12668
rect 35391 12665 35403 12699
rect 35345 12659 35403 12665
rect 33042 12628 33048 12640
rect 31726 12600 33048 12628
rect 33042 12588 33048 12600
rect 33100 12588 33106 12640
rect 34149 12631 34207 12637
rect 34149 12597 34161 12631
rect 34195 12628 34207 12631
rect 36170 12628 36176 12640
rect 34195 12600 36176 12628
rect 34195 12597 34207 12600
rect 34149 12591 34207 12597
rect 36170 12588 36176 12600
rect 36228 12588 36234 12640
rect 38194 12628 38200 12640
rect 38155 12600 38200 12628
rect 38194 12588 38200 12600
rect 38252 12588 38258 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 4890 12424 4896 12436
rect 4851 12396 4896 12424
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 16942 12424 16948 12436
rect 14415 12396 16948 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 19705 12427 19763 12433
rect 19705 12393 19717 12427
rect 19751 12424 19763 12427
rect 19886 12424 19892 12436
rect 19751 12396 19892 12424
rect 19751 12393 19763 12396
rect 19705 12387 19763 12393
rect 19886 12384 19892 12396
rect 19944 12384 19950 12436
rect 31018 12384 31024 12436
rect 31076 12424 31082 12436
rect 33873 12427 33931 12433
rect 31076 12396 31800 12424
rect 31076 12384 31082 12396
rect 18598 12316 18604 12368
rect 18656 12356 18662 12368
rect 24486 12356 24492 12368
rect 18656 12328 24492 12356
rect 18656 12316 18662 12328
rect 24486 12316 24492 12328
rect 24544 12316 24550 12368
rect 30650 12316 30656 12368
rect 30708 12356 30714 12368
rect 31386 12356 31392 12368
rect 30708 12328 31392 12356
rect 30708 12316 30714 12328
rect 31386 12316 31392 12328
rect 31444 12316 31450 12368
rect 31772 12356 31800 12396
rect 33873 12393 33885 12427
rect 33919 12424 33931 12427
rect 34514 12424 34520 12436
rect 33919 12396 34520 12424
rect 33919 12393 33931 12396
rect 33873 12387 33931 12393
rect 34514 12384 34520 12396
rect 34572 12384 34578 12436
rect 34698 12384 34704 12436
rect 34756 12424 34762 12436
rect 35342 12424 35348 12436
rect 34756 12396 35348 12424
rect 34756 12384 34762 12396
rect 35342 12384 35348 12396
rect 35400 12384 35406 12436
rect 36998 12384 37004 12436
rect 37056 12424 37062 12436
rect 37737 12427 37795 12433
rect 37737 12424 37749 12427
rect 37056 12396 37749 12424
rect 37056 12384 37062 12396
rect 37737 12393 37749 12396
rect 37783 12393 37795 12427
rect 37737 12387 37795 12393
rect 31772 12328 35894 12356
rect 22002 12288 22008 12300
rect 19904 12260 22008 12288
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 1544 12192 4813 12220
rect 1544 12180 1550 12192
rect 4801 12189 4813 12192
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 19904 12229 19932 12260
rect 22002 12248 22008 12260
rect 22060 12248 22066 12300
rect 23934 12288 23940 12300
rect 22756 12260 23796 12288
rect 23895 12260 23940 12288
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13228 12192 14289 12220
rect 13228 12180 13234 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12220 20407 12223
rect 22756 12220 22784 12260
rect 20395 12192 22784 12220
rect 23768 12220 23796 12260
rect 23934 12248 23940 12260
rect 23992 12248 23998 12300
rect 25222 12288 25228 12300
rect 24044 12260 25228 12288
rect 24044 12220 24072 12260
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 29822 12288 29828 12300
rect 29783 12260 29828 12288
rect 29822 12248 29828 12260
rect 29880 12248 29886 12300
rect 30469 12291 30527 12297
rect 30469 12257 30481 12291
rect 30515 12288 30527 12291
rect 31297 12291 31355 12297
rect 31297 12288 31309 12291
rect 30515 12260 31309 12288
rect 30515 12257 30527 12260
rect 30469 12251 30527 12257
rect 31297 12257 31309 12260
rect 31343 12288 31355 12291
rect 34698 12288 34704 12300
rect 31343 12260 34704 12288
rect 31343 12257 31355 12260
rect 31297 12251 31355 12257
rect 34698 12248 34704 12260
rect 34756 12248 34762 12300
rect 34992 12297 35020 12328
rect 34977 12291 35035 12297
rect 34977 12257 34989 12291
rect 35023 12257 35035 12291
rect 35618 12288 35624 12300
rect 35579 12260 35624 12288
rect 34977 12251 35035 12257
rect 35618 12248 35624 12260
rect 35676 12248 35682 12300
rect 35866 12288 35894 12328
rect 37001 12291 37059 12297
rect 37001 12288 37013 12291
rect 35866 12260 37013 12288
rect 37001 12257 37013 12260
rect 37047 12257 37059 12291
rect 37001 12251 37059 12257
rect 23768 12192 24072 12220
rect 20395 12189 20407 12192
rect 20349 12183 20407 12189
rect 29638 12180 29644 12232
rect 29696 12180 29702 12232
rect 32309 12223 32367 12229
rect 32309 12189 32321 12223
rect 32355 12189 32367 12223
rect 32309 12183 32367 12189
rect 22278 12112 22284 12164
rect 22336 12152 22342 12164
rect 22925 12155 22983 12161
rect 22925 12152 22937 12155
rect 22336 12124 22937 12152
rect 22336 12112 22342 12124
rect 22925 12121 22937 12124
rect 22971 12121 22983 12155
rect 22925 12115 22983 12121
rect 23017 12155 23075 12161
rect 23017 12121 23029 12155
rect 23063 12152 23075 12155
rect 23198 12152 23204 12164
rect 23063 12124 23204 12152
rect 23063 12121 23075 12124
rect 23017 12115 23075 12121
rect 23198 12112 23204 12124
rect 23256 12112 23262 12164
rect 24670 12152 24676 12164
rect 24631 12124 24676 12152
rect 24670 12112 24676 12124
rect 24728 12112 24734 12164
rect 24765 12155 24823 12161
rect 24765 12121 24777 12155
rect 24811 12121 24823 12155
rect 25682 12152 25688 12164
rect 25643 12124 25688 12152
rect 24765 12115 24823 12121
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 20128 12056 20453 12084
rect 20128 12044 20134 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 23658 12044 23664 12096
rect 23716 12084 23722 12096
rect 24780 12084 24808 12115
rect 25682 12112 25688 12124
rect 25740 12112 25746 12164
rect 29656 12152 29684 12180
rect 29894 12155 29952 12161
rect 29894 12152 29906 12155
rect 29656 12124 29906 12152
rect 29894 12121 29906 12124
rect 29940 12121 29952 12155
rect 31021 12155 31079 12161
rect 31021 12152 31033 12155
rect 29894 12115 29952 12121
rect 30116 12124 31033 12152
rect 23716 12056 24808 12084
rect 23716 12044 23722 12056
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 30116 12084 30144 12124
rect 31021 12121 31033 12124
rect 31067 12121 31079 12155
rect 31021 12115 31079 12121
rect 31110 12112 31116 12164
rect 31168 12152 31174 12164
rect 31168 12124 31213 12152
rect 31168 12112 31174 12124
rect 31386 12112 31392 12164
rect 31444 12152 31450 12164
rect 32324 12152 32352 12183
rect 32950 12180 32956 12232
rect 33008 12220 33014 12232
rect 33413 12223 33471 12229
rect 33413 12220 33425 12223
rect 33008 12192 33425 12220
rect 33008 12180 33014 12192
rect 33413 12189 33425 12192
rect 33459 12189 33471 12223
rect 33413 12183 33471 12189
rect 34057 12223 34115 12229
rect 34057 12189 34069 12223
rect 34103 12189 34115 12223
rect 34057 12183 34115 12189
rect 36909 12223 36967 12229
rect 36909 12189 36921 12223
rect 36955 12189 36967 12223
rect 36909 12183 36967 12189
rect 37645 12223 37703 12229
rect 37645 12189 37657 12223
rect 37691 12220 37703 12223
rect 39022 12220 39028 12232
rect 37691 12192 39028 12220
rect 37691 12189 37703 12192
rect 37645 12183 37703 12189
rect 34072 12152 34100 12183
rect 31444 12124 32352 12152
rect 32416 12124 34100 12152
rect 31444 12112 31450 12124
rect 32122 12084 32128 12096
rect 26660 12056 30144 12084
rect 32083 12056 32128 12084
rect 26660 12044 26666 12056
rect 32122 12044 32128 12056
rect 32180 12044 32186 12096
rect 32214 12044 32220 12096
rect 32272 12084 32278 12096
rect 32416 12084 32444 12124
rect 35066 12112 35072 12164
rect 35124 12152 35130 12164
rect 36924 12152 36952 12183
rect 39022 12180 39028 12192
rect 39080 12180 39086 12232
rect 37734 12152 37740 12164
rect 35124 12124 35169 12152
rect 36924 12124 37740 12152
rect 35124 12112 35130 12124
rect 37734 12112 37740 12124
rect 37792 12112 37798 12164
rect 33226 12084 33232 12096
rect 32272 12056 32444 12084
rect 33187 12056 33232 12084
rect 32272 12044 32278 12056
rect 33226 12044 33232 12056
rect 33284 12044 33290 12096
rect 34606 12044 34612 12096
rect 34664 12084 34670 12096
rect 36081 12087 36139 12093
rect 36081 12084 36093 12087
rect 34664 12056 36093 12084
rect 34664 12044 34670 12056
rect 36081 12053 36093 12056
rect 36127 12053 36139 12087
rect 36081 12047 36139 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 12618 11880 12624 11892
rect 12579 11852 12624 11880
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 17034 11880 17040 11892
rect 16255 11852 17040 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 29641 11883 29699 11889
rect 21508 11852 26464 11880
rect 21508 11840 21514 11852
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16945 11815 17003 11821
rect 16080 11784 16896 11812
rect 16080 11772 16086 11784
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 9030 11744 9036 11756
rect 6963 11716 9036 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 12526 11744 12532 11756
rect 12487 11716 12532 11744
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11744 16175 11747
rect 16758 11744 16764 11756
rect 16163 11716 16764 11744
rect 16163 11713 16175 11716
rect 16117 11707 16175 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16868 11753 16896 11784
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 16991 11784 17693 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 17681 11781 17693 11784
rect 17727 11781 17739 11815
rect 18598 11812 18604 11824
rect 18559 11784 18604 11812
rect 17681 11775 17739 11781
rect 18598 11772 18604 11784
rect 18656 11772 18662 11824
rect 20070 11812 20076 11824
rect 20031 11784 20076 11812
rect 20070 11772 20076 11784
rect 20128 11772 20134 11824
rect 20898 11772 20904 11824
rect 20956 11812 20962 11824
rect 20993 11815 21051 11821
rect 20993 11812 21005 11815
rect 20956 11784 21005 11812
rect 20956 11772 20962 11784
rect 20993 11781 21005 11784
rect 21039 11781 21051 11815
rect 23750 11812 23756 11824
rect 20993 11775 21051 11781
rect 22020 11784 23756 11812
rect 22020 11753 22048 11784
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 25406 11812 25412 11824
rect 25367 11784 25412 11812
rect 25406 11772 25412 11784
rect 25464 11772 25470 11824
rect 26436 11753 26464 11852
rect 29641 11849 29653 11883
rect 29687 11880 29699 11883
rect 30374 11880 30380 11892
rect 29687 11852 30380 11880
rect 29687 11849 29699 11852
rect 29641 11843 29699 11849
rect 30374 11840 30380 11852
rect 30432 11840 30438 11892
rect 32950 11880 32956 11892
rect 32911 11852 32956 11880
rect 32950 11840 32956 11852
rect 33008 11840 33014 11892
rect 34514 11880 34520 11892
rect 33060 11852 34520 11880
rect 30742 11812 30748 11824
rect 29564 11784 30748 11812
rect 29564 11753 29592 11784
rect 30742 11772 30748 11784
rect 30800 11772 30806 11824
rect 30837 11815 30895 11821
rect 30837 11781 30849 11815
rect 30883 11812 30895 11815
rect 30926 11812 30932 11824
rect 30883 11784 30932 11812
rect 30883 11781 30895 11784
rect 30837 11775 30895 11781
rect 30926 11772 30932 11784
rect 30984 11772 30990 11824
rect 31570 11772 31576 11824
rect 31628 11772 31634 11824
rect 31662 11772 31668 11824
rect 31720 11812 31726 11824
rect 31757 11815 31815 11821
rect 31757 11812 31769 11815
rect 31720 11784 31769 11812
rect 31720 11772 31726 11784
rect 31757 11781 31769 11784
rect 31803 11812 31815 11815
rect 33060 11812 33088 11852
rect 34514 11840 34520 11852
rect 34572 11840 34578 11892
rect 35710 11840 35716 11892
rect 35768 11880 35774 11892
rect 36541 11883 36599 11889
rect 36541 11880 36553 11883
rect 35768 11852 36553 11880
rect 35768 11840 35774 11852
rect 36541 11849 36553 11852
rect 36587 11849 36599 11883
rect 36541 11843 36599 11849
rect 31803 11784 33088 11812
rect 31803 11781 31815 11784
rect 31757 11775 31815 11781
rect 34422 11772 34428 11824
rect 34480 11812 34486 11824
rect 34480 11784 35204 11812
rect 34480 11772 34486 11784
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 22005 11747 22063 11753
rect 16853 11707 16911 11713
rect 18524 11716 18828 11744
rect 16868 11608 16896 11707
rect 17589 11679 17647 11685
rect 17589 11645 17601 11679
rect 17635 11676 17647 11679
rect 18524 11676 18552 11716
rect 18800 11688 18828 11716
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11713 22707 11747
rect 22649 11707 22707 11713
rect 26421 11747 26479 11753
rect 26421 11713 26433 11747
rect 26467 11713 26479 11747
rect 26421 11707 26479 11713
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11713 29607 11747
rect 31588 11744 31616 11772
rect 32309 11747 32367 11753
rect 32309 11744 32321 11747
rect 31588 11716 32321 11744
rect 29549 11707 29607 11713
rect 32309 11713 32321 11716
rect 32355 11713 32367 11747
rect 33137 11747 33195 11753
rect 33137 11744 33149 11747
rect 32309 11707 32367 11713
rect 32416 11716 33149 11744
rect 17635 11648 18552 11676
rect 17635 11645 17647 11648
rect 17589 11639 17647 11645
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 18840 11648 19993 11676
rect 18840 11636 18846 11648
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 22020 11676 22048 11707
rect 20128 11648 22048 11676
rect 20128 11636 20134 11648
rect 22664 11608 22692 11707
rect 25317 11679 25375 11685
rect 25317 11645 25329 11679
rect 25363 11676 25375 11679
rect 27246 11676 27252 11688
rect 25363 11648 27252 11676
rect 25363 11645 25375 11648
rect 25317 11639 25375 11645
rect 27246 11636 27252 11648
rect 27304 11636 27310 11688
rect 30745 11679 30803 11685
rect 30745 11645 30757 11679
rect 30791 11676 30803 11679
rect 31294 11676 31300 11688
rect 30791 11648 31300 11676
rect 30791 11645 30803 11648
rect 30745 11639 30803 11645
rect 31294 11636 31300 11648
rect 31352 11636 31358 11688
rect 32214 11676 32220 11688
rect 31726 11648 32220 11676
rect 16868 11580 22692 11608
rect 24854 11568 24860 11620
rect 24912 11608 24918 11620
rect 25866 11608 25872 11620
rect 24912 11580 25872 11608
rect 24912 11568 24918 11580
rect 25866 11568 25872 11580
rect 25924 11568 25930 11620
rect 30190 11568 30196 11620
rect 30248 11608 30254 11620
rect 31726 11608 31754 11648
rect 32214 11636 32220 11648
rect 32272 11636 32278 11688
rect 32416 11608 32444 11716
rect 33137 11713 33149 11716
rect 33183 11713 33195 11747
rect 33137 11707 33195 11713
rect 33226 11704 33232 11756
rect 33284 11744 33290 11756
rect 34793 11747 34851 11753
rect 34793 11744 34805 11747
rect 33284 11716 34805 11744
rect 33284 11704 33290 11716
rect 34793 11713 34805 11716
rect 34839 11713 34851 11747
rect 34793 11707 34851 11713
rect 34606 11676 34612 11688
rect 34567 11648 34612 11676
rect 34606 11636 34612 11648
rect 34664 11636 34670 11688
rect 35176 11676 35204 11784
rect 35434 11704 35440 11756
rect 35492 11744 35498 11756
rect 35805 11747 35863 11753
rect 35805 11744 35817 11747
rect 35492 11716 35817 11744
rect 35492 11704 35498 11716
rect 35805 11713 35817 11716
rect 35851 11713 35863 11747
rect 36446 11744 36452 11756
rect 36407 11716 36452 11744
rect 35805 11707 35863 11713
rect 36446 11704 36452 11716
rect 36504 11704 36510 11756
rect 37550 11704 37556 11756
rect 37608 11744 37614 11756
rect 37737 11747 37795 11753
rect 37737 11744 37749 11747
rect 37608 11716 37749 11744
rect 37608 11704 37614 11716
rect 37737 11713 37749 11716
rect 37783 11713 37795 11747
rect 37737 11707 37795 11713
rect 35897 11679 35955 11685
rect 35897 11676 35909 11679
rect 35176 11648 35909 11676
rect 35897 11645 35909 11648
rect 35943 11645 35955 11679
rect 35897 11639 35955 11645
rect 30248 11580 31754 11608
rect 32232 11580 32444 11608
rect 30248 11568 30254 11580
rect 6733 11543 6791 11549
rect 6733 11509 6745 11543
rect 6779 11540 6791 11543
rect 7558 11540 7564 11552
rect 6779 11512 7564 11540
rect 6779 11509 6791 11512
rect 6733 11503 6791 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 13538 11540 13544 11552
rect 9088 11512 13544 11540
rect 9088 11500 9094 11512
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 22097 11543 22155 11549
rect 22097 11540 22109 11543
rect 21324 11512 22109 11540
rect 21324 11500 21330 11512
rect 22097 11509 22109 11512
rect 22143 11509 22155 11543
rect 22097 11503 22155 11509
rect 22741 11543 22799 11549
rect 22741 11509 22753 11543
rect 22787 11540 22799 11543
rect 23474 11540 23480 11552
rect 22787 11512 23480 11540
rect 22787 11509 22799 11512
rect 22741 11503 22799 11509
rect 23474 11500 23480 11512
rect 23532 11500 23538 11552
rect 26513 11543 26571 11549
rect 26513 11509 26525 11543
rect 26559 11540 26571 11543
rect 27338 11540 27344 11552
rect 26559 11512 27344 11540
rect 26559 11509 26571 11512
rect 26513 11503 26571 11509
rect 27338 11500 27344 11512
rect 27396 11500 27402 11552
rect 30742 11500 30748 11552
rect 30800 11540 30806 11552
rect 32232 11540 32260 11580
rect 33042 11568 33048 11620
rect 33100 11608 33106 11620
rect 34790 11608 34796 11620
rect 33100 11580 34796 11608
rect 33100 11568 33106 11580
rect 34790 11568 34796 11580
rect 34848 11608 34854 11620
rect 34977 11611 35035 11617
rect 34977 11608 34989 11611
rect 34848 11580 34989 11608
rect 34848 11568 34854 11580
rect 34977 11577 34989 11580
rect 35023 11577 35035 11611
rect 34977 11571 35035 11577
rect 32398 11540 32404 11552
rect 30800 11512 32260 11540
rect 32359 11512 32404 11540
rect 30800 11500 30806 11512
rect 32398 11500 32404 11512
rect 32456 11500 32462 11552
rect 37826 11540 37832 11552
rect 37787 11512 37832 11540
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 9030 11336 9036 11348
rect 1811 11308 9036 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9180 11308 9689 11336
rect 9180 11296 9186 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 10376 11308 10793 11336
rect 10376 11296 10382 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 19981 11339 20039 11345
rect 19981 11336 19993 11339
rect 10781 11299 10839 11305
rect 16546 11308 19993 11336
rect 7377 11271 7435 11277
rect 7377 11237 7389 11271
rect 7423 11268 7435 11271
rect 7423 11240 9352 11268
rect 7423 11237 7435 11240
rect 7377 11231 7435 11237
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 8570 11200 8576 11212
rect 6595 11172 8576 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 9324 11209 9352 11240
rect 9309 11203 9367 11209
rect 9309 11169 9321 11203
rect 9355 11169 9367 11203
rect 16546 11200 16574 11308
rect 19981 11305 19993 11308
rect 20027 11305 20039 11339
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 19981 11299 20039 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 29638 11296 29644 11348
rect 29696 11336 29702 11348
rect 29917 11339 29975 11345
rect 29917 11336 29929 11339
rect 29696 11308 29929 11336
rect 29696 11296 29702 11308
rect 29917 11305 29929 11308
rect 29963 11305 29975 11339
rect 29917 11299 29975 11305
rect 30745 11339 30803 11345
rect 30745 11305 30757 11339
rect 30791 11336 30803 11339
rect 31110 11336 31116 11348
rect 30791 11308 31116 11336
rect 30791 11305 30803 11308
rect 30745 11299 30803 11305
rect 31110 11296 31116 11308
rect 31168 11296 31174 11348
rect 35986 11336 35992 11348
rect 31726 11308 35992 11336
rect 18417 11271 18475 11277
rect 18417 11237 18429 11271
rect 18463 11268 18475 11271
rect 18782 11268 18788 11280
rect 18463 11240 18788 11268
rect 18463 11237 18475 11240
rect 18417 11231 18475 11237
rect 18782 11228 18788 11240
rect 18840 11228 18846 11280
rect 20990 11228 20996 11280
rect 21048 11268 21054 11280
rect 21453 11271 21511 11277
rect 21453 11268 21465 11271
rect 21048 11240 21465 11268
rect 21048 11228 21054 11240
rect 21453 11237 21465 11240
rect 21499 11237 21511 11271
rect 21453 11231 21511 11237
rect 25682 11228 25688 11280
rect 25740 11268 25746 11280
rect 31726 11268 31754 11308
rect 35986 11296 35992 11308
rect 36044 11296 36050 11348
rect 25740 11240 31754 11268
rect 35529 11271 35587 11277
rect 25740 11228 25746 11240
rect 35529 11237 35541 11271
rect 35575 11268 35587 11271
rect 38010 11268 38016 11280
rect 35575 11240 38016 11268
rect 35575 11237 35587 11240
rect 35529 11231 35587 11237
rect 38010 11228 38016 11240
rect 38068 11228 38074 11280
rect 21266 11200 21272 11212
rect 9309 11163 9367 11169
rect 10612 11172 16574 11200
rect 21227 11172 21272 11200
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 3476 11104 6469 11132
rect 3476 11092 3482 11104
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 7558 11132 7564 11144
rect 7519 11104 7564 11132
rect 6457 11095 6515 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 9122 11132 9128 11144
rect 9083 11104 9128 11132
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 1670 11064 1676 11076
rect 1631 11036 1676 11064
rect 1670 11024 1676 11036
rect 1728 11024 1734 11076
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 10612 11064 10640 11172
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 22370 11200 22376 11212
rect 21376 11172 22376 11200
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 12986 11132 12992 11144
rect 10735 11104 12992 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 14918 11132 14924 11144
rect 13311 11104 14924 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15838 11132 15844 11144
rect 15799 11104 15844 11132
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 18138 11092 18144 11144
rect 18196 11132 18202 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 18196 11104 18337 11132
rect 18196 11092 18202 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21376 11132 21404 11172
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 31294 11200 31300 11212
rect 31255 11172 31300 11200
rect 31294 11160 31300 11172
rect 31352 11160 31358 11212
rect 37550 11160 37556 11212
rect 37608 11200 37614 11212
rect 37829 11203 37887 11209
rect 37829 11200 37841 11203
rect 37608 11172 37841 11200
rect 37608 11160 37614 11172
rect 37829 11169 37841 11172
rect 37875 11169 37887 11203
rect 37829 11163 37887 11169
rect 21131 11104 21404 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22189 11135 22247 11141
rect 22189 11132 22201 11135
rect 22152 11104 22201 11132
rect 22152 11092 22158 11104
rect 22189 11101 22201 11104
rect 22235 11101 22247 11135
rect 22189 11095 22247 11101
rect 30101 11135 30159 11141
rect 30101 11101 30113 11135
rect 30147 11101 30159 11135
rect 30650 11132 30656 11144
rect 30611 11104 30656 11132
rect 30101 11095 30159 11101
rect 4028 11036 10640 11064
rect 4028 11024 4034 11036
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 13449 11067 13507 11073
rect 13449 11064 13461 11067
rect 13412 11036 13461 11064
rect 13412 11024 13418 11036
rect 13449 11033 13461 11036
rect 13495 11033 13507 11067
rect 13449 11027 13507 11033
rect 19889 11067 19947 11073
rect 19889 11033 19901 11067
rect 19935 11064 19947 11067
rect 22554 11064 22560 11076
rect 19935 11036 22560 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 30116 11064 30144 11095
rect 30650 11092 30656 11104
rect 30708 11092 30714 11144
rect 34790 11092 34796 11144
rect 34848 11132 34854 11144
rect 34885 11135 34943 11141
rect 34885 11132 34897 11135
rect 34848 11104 34897 11132
rect 34848 11092 34854 11104
rect 34885 11101 34897 11104
rect 34931 11101 34943 11135
rect 34885 11095 34943 11101
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11132 35035 11135
rect 35713 11135 35771 11141
rect 35713 11132 35725 11135
rect 35023 11104 35725 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 35713 11101 35725 11104
rect 35759 11101 35771 11135
rect 36814 11132 36820 11144
rect 36775 11104 36820 11132
rect 35713 11095 35771 11101
rect 36814 11092 36820 11104
rect 36872 11092 36878 11144
rect 32122 11064 32128 11076
rect 30116 11036 32128 11064
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 36722 11024 36728 11076
rect 36780 11064 36786 11076
rect 37001 11067 37059 11073
rect 37001 11064 37013 11067
rect 36780 11036 37013 11064
rect 36780 11024 36786 11036
rect 37001 11033 37013 11036
rect 37047 11033 37059 11067
rect 37550 11064 37556 11076
rect 37511 11036 37556 11064
rect 37001 11027 37059 11033
rect 37550 11024 37556 11036
rect 37608 11024 37614 11076
rect 37642 11024 37648 11076
rect 37700 11064 37706 11076
rect 37700 11036 37745 11064
rect 37700 11024 37706 11036
rect 15930 10996 15936 11008
rect 15891 10968 15936 10996
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 28902 10996 28908 11008
rect 28863 10968 28908 10996
rect 28902 10956 28908 10968
rect 28960 10956 28966 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 4614 10792 4620 10804
rect 1627 10764 4620 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 8996 10764 9137 10792
rect 8996 10752 9002 10764
rect 9125 10761 9137 10764
rect 9171 10761 9183 10795
rect 16022 10792 16028 10804
rect 9125 10755 9183 10761
rect 14844 10764 16028 10792
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10656 14611 10659
rect 14844 10656 14872 10764
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 24670 10792 24676 10804
rect 20119 10764 24676 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 29549 10795 29607 10801
rect 29549 10761 29561 10795
rect 29595 10792 29607 10795
rect 29822 10792 29828 10804
rect 29595 10764 29828 10792
rect 29595 10761 29607 10764
rect 29549 10755 29607 10761
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 35989 10795 36047 10801
rect 35989 10761 36001 10795
rect 36035 10792 36047 10795
rect 36354 10792 36360 10804
rect 36035 10764 36360 10792
rect 36035 10761 36047 10764
rect 35989 10755 36047 10761
rect 36354 10752 36360 10764
rect 36412 10752 36418 10804
rect 38194 10792 38200 10804
rect 38155 10764 38200 10792
rect 38194 10752 38200 10764
rect 38252 10752 38258 10804
rect 14918 10684 14924 10736
rect 14976 10724 14982 10736
rect 22554 10724 22560 10736
rect 14976 10696 22560 10724
rect 14976 10684 14982 10696
rect 22554 10684 22560 10696
rect 22612 10684 22618 10736
rect 27338 10724 27344 10736
rect 27299 10696 27344 10724
rect 27338 10684 27344 10696
rect 27396 10684 27402 10736
rect 27893 10727 27951 10733
rect 27893 10693 27905 10727
rect 27939 10724 27951 10727
rect 28350 10724 28356 10736
rect 27939 10696 28356 10724
rect 27939 10693 27951 10696
rect 27893 10687 27951 10693
rect 28350 10684 28356 10696
rect 28408 10684 28414 10736
rect 35434 10684 35440 10736
rect 35492 10724 35498 10736
rect 35492 10696 36952 10724
rect 35492 10684 35498 10696
rect 15194 10656 15200 10668
rect 14599 10628 14872 10656
rect 15155 10628 15200 10656
rect 14599 10625 14611 10628
rect 14553 10619 14611 10625
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 15930 10656 15936 10668
rect 15427 10628 15936 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 19981 10659 20039 10665
rect 19981 10656 19993 10659
rect 16546 10628 19993 10656
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 16546 10588 16574 10628
rect 19981 10625 19993 10628
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22278 10656 22284 10668
rect 22235 10628 22284 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 24121 10659 24179 10665
rect 24121 10625 24133 10659
rect 24167 10656 24179 10659
rect 25222 10656 25228 10668
rect 24167 10628 25228 10656
rect 24167 10625 24179 10628
rect 24121 10619 24179 10625
rect 25222 10616 25228 10628
rect 25280 10616 25286 10668
rect 28902 10656 28908 10668
rect 28863 10628 28908 10656
rect 28902 10616 28908 10628
rect 28960 10616 28966 10668
rect 30009 10659 30067 10665
rect 30009 10625 30021 10659
rect 30055 10656 30067 10659
rect 36170 10656 36176 10668
rect 30055 10628 35894 10656
rect 36131 10628 36176 10656
rect 30055 10625 30067 10628
rect 30009 10619 30067 10625
rect 27246 10588 27252 10600
rect 14332 10560 16574 10588
rect 27207 10560 27252 10588
rect 14332 10548 14338 10560
rect 27246 10548 27252 10560
rect 27304 10588 27310 10600
rect 29086 10588 29092 10600
rect 27304 10560 28304 10588
rect 29047 10560 29092 10588
rect 27304 10548 27310 10560
rect 16850 10480 16856 10532
rect 16908 10520 16914 10532
rect 17770 10520 17776 10532
rect 16908 10492 17776 10520
rect 16908 10480 16914 10492
rect 17770 10480 17776 10492
rect 17828 10520 17834 10532
rect 25498 10520 25504 10532
rect 17828 10492 25504 10520
rect 17828 10480 17834 10492
rect 25498 10480 25504 10492
rect 25556 10480 25562 10532
rect 28276 10520 28304 10560
rect 29086 10548 29092 10560
rect 29144 10548 29150 10600
rect 35866 10588 35894 10628
rect 36170 10616 36176 10628
rect 36228 10616 36234 10668
rect 36924 10665 36952 10696
rect 36909 10659 36967 10665
rect 36909 10625 36921 10659
rect 36955 10625 36967 10659
rect 38010 10656 38016 10668
rect 37971 10628 38016 10656
rect 36909 10619 36967 10625
rect 38010 10616 38016 10628
rect 38068 10616 38074 10668
rect 38102 10588 38108 10600
rect 35866 10560 38108 10588
rect 38102 10548 38108 10560
rect 38160 10548 38166 10600
rect 30101 10523 30159 10529
rect 30101 10520 30113 10523
rect 28276 10492 30113 10520
rect 30101 10489 30113 10492
rect 30147 10489 30159 10523
rect 30101 10483 30159 10489
rect 14642 10452 14648 10464
rect 14603 10424 14648 10452
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 15841 10455 15899 10461
rect 15841 10421 15853 10455
rect 15887 10452 15899 10455
rect 16114 10452 16120 10464
rect 15887 10424 16120 10452
rect 15887 10421 15899 10424
rect 15841 10415 15899 10421
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 22281 10455 22339 10461
rect 22281 10421 22293 10455
rect 22327 10452 22339 10455
rect 22646 10452 22652 10464
rect 22327 10424 22652 10452
rect 22327 10421 22339 10424
rect 22281 10415 22339 10421
rect 22646 10412 22652 10424
rect 22704 10412 22710 10464
rect 24213 10455 24271 10461
rect 24213 10421 24225 10455
rect 24259 10452 24271 10455
rect 24762 10452 24768 10464
rect 24259 10424 24768 10452
rect 24259 10421 24271 10424
rect 24213 10415 24271 10421
rect 24762 10412 24768 10424
rect 24820 10412 24826 10464
rect 36725 10455 36783 10461
rect 36725 10421 36737 10455
rect 36771 10452 36783 10455
rect 37918 10452 37924 10464
rect 36771 10424 37924 10452
rect 36771 10421 36783 10424
rect 36725 10415 36783 10421
rect 37918 10412 37924 10424
rect 37976 10412 37982 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 16114 10208 16120 10220
rect 16172 10248 16178 10260
rect 17862 10248 17868 10260
rect 16172 10220 17868 10248
rect 16172 10208 16178 10220
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 26234 10208 26240 10260
rect 26292 10248 26298 10260
rect 27341 10251 27399 10257
rect 27341 10248 27353 10251
rect 26292 10220 27353 10248
rect 26292 10208 26298 10220
rect 27341 10217 27353 10220
rect 27387 10217 27399 10251
rect 30466 10248 30472 10260
rect 30427 10220 30472 10248
rect 27341 10211 27399 10217
rect 30466 10208 30472 10220
rect 30524 10208 30530 10260
rect 36725 10251 36783 10257
rect 36725 10217 36737 10251
rect 36771 10248 36783 10251
rect 37366 10248 37372 10260
rect 36771 10220 37372 10248
rect 36771 10217 36783 10220
rect 36725 10211 36783 10217
rect 37366 10208 37372 10220
rect 37424 10208 37430 10260
rect 38194 10248 38200 10260
rect 38155 10220 38200 10248
rect 38194 10208 38200 10220
rect 38252 10208 38258 10260
rect 22462 10140 22468 10192
rect 22520 10180 22526 10192
rect 25225 10183 25283 10189
rect 22520 10152 24624 10180
rect 22520 10140 22526 10152
rect 22554 10112 22560 10124
rect 22515 10084 22560 10112
rect 22554 10072 22560 10084
rect 22612 10072 22618 10124
rect 24596 10121 24624 10152
rect 25225 10149 25237 10183
rect 25271 10180 25283 10183
rect 29822 10180 29828 10192
rect 25271 10152 29828 10180
rect 25271 10149 25283 10152
rect 25225 10143 25283 10149
rect 29822 10140 29828 10152
rect 29880 10140 29886 10192
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 2225 10047 2283 10053
rect 2225 10013 2237 10047
rect 2271 10044 2283 10047
rect 10134 10044 10140 10056
rect 2271 10016 10140 10044
rect 2271 10013 2283 10016
rect 2225 10007 2283 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 12434 10044 12440 10056
rect 12395 10016 12440 10044
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12618 10044 12624 10056
rect 12579 10016 12624 10044
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 17770 10044 17776 10056
rect 17731 10016 17776 10044
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 21450 10044 21456 10056
rect 21411 10016 21456 10044
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 24765 10047 24823 10053
rect 24765 10013 24777 10047
rect 24811 10044 24823 10047
rect 24946 10044 24952 10056
rect 24811 10016 24952 10044
rect 24811 10013 24823 10016
rect 24765 10007 24823 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 27249 10047 27307 10053
rect 27249 10013 27261 10047
rect 27295 10013 27307 10047
rect 30374 10044 30380 10056
rect 30335 10016 30380 10044
rect 27249 10007 27307 10013
rect 22646 9936 22652 9988
rect 22704 9976 22710 9988
rect 23569 9979 23627 9985
rect 22704 9948 22749 9976
rect 22704 9936 22710 9948
rect 23569 9945 23581 9979
rect 23615 9945 23627 9979
rect 23569 9939 23627 9945
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2225 9911 2283 9917
rect 2225 9908 2237 9911
rect 2096 9880 2237 9908
rect 2096 9868 2102 9880
rect 2225 9877 2237 9880
rect 2271 9877 2283 9911
rect 2225 9871 2283 9877
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 14918 9908 14924 9920
rect 13127 9880 14924 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 17034 9868 17040 9920
rect 17092 9908 17098 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17092 9880 17877 9908
rect 17092 9868 17098 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 21545 9911 21603 9917
rect 21545 9877 21557 9911
rect 21591 9908 21603 9911
rect 22186 9908 22192 9920
rect 21591 9880 22192 9908
rect 21591 9877 21603 9880
rect 21545 9871 21603 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 23584 9908 23612 9939
rect 24670 9936 24676 9988
rect 24728 9976 24734 9988
rect 27264 9976 27292 10007
rect 30374 10004 30380 10016
rect 30432 10004 30438 10056
rect 36906 10044 36912 10056
rect 36867 10016 36912 10044
rect 36906 10004 36912 10016
rect 36964 10004 36970 10056
rect 37553 10047 37611 10053
rect 37553 10013 37565 10047
rect 37599 10044 37611 10047
rect 37826 10044 37832 10056
rect 37599 10016 37832 10044
rect 37599 10013 37611 10016
rect 37553 10007 37611 10013
rect 37826 10004 37832 10016
rect 37884 10004 37890 10056
rect 38013 10047 38071 10053
rect 38013 10013 38025 10047
rect 38059 10013 38071 10047
rect 38013 10007 38071 10013
rect 38028 9976 38056 10007
rect 24728 9948 27292 9976
rect 37384 9948 38056 9976
rect 24728 9936 24734 9948
rect 27706 9908 27712 9920
rect 23584 9880 27712 9908
rect 27706 9868 27712 9880
rect 27764 9868 27770 9920
rect 37384 9917 37412 9948
rect 37369 9911 37427 9917
rect 37369 9877 37381 9911
rect 37415 9877 37427 9911
rect 37369 9871 37427 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 12434 9704 12440 9716
rect 12395 9676 12440 9704
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 12676 9676 13185 9704
rect 12676 9664 12682 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 15746 9704 15752 9716
rect 15707 9676 15752 9704
rect 13173 9667 13231 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 23308 9676 23612 9704
rect 15838 9636 15844 9648
rect 14660 9608 15844 9636
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 14660 9577 14688 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 17034 9636 17040 9648
rect 16995 9608 17040 9636
rect 17034 9596 17040 9608
rect 17092 9596 17098 9648
rect 20990 9636 20996 9648
rect 20951 9608 20996 9636
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 22738 9636 22744 9648
rect 22066 9608 22744 9636
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20070 9568 20076 9580
rect 19935 9540 20076 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 15304 9500 15332 9531
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 14476 9472 15332 9500
rect 16546 9472 16957 9500
rect 14476 9441 14504 9472
rect 14461 9435 14519 9441
rect 14461 9401 14473 9435
rect 14507 9401 14519 9435
rect 14461 9395 14519 9401
rect 15105 9435 15163 9441
rect 15105 9401 15117 9435
rect 15151 9432 15163 9435
rect 15930 9432 15936 9444
rect 15151 9404 15936 9432
rect 15151 9401 15163 9404
rect 15105 9395 15163 9401
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1636 9336 1869 9364
rect 1636 9324 1642 9336
rect 1857 9333 1869 9336
rect 1903 9333 1915 9367
rect 1857 9327 1915 9333
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 16546 9364 16574 9472
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 17920 9472 20361 9500
rect 17920 9460 17926 9472
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20530 9500 20536 9512
rect 20491 9472 20536 9500
rect 20349 9463 20407 9469
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 17497 9435 17555 9441
rect 17497 9401 17509 9435
rect 17543 9432 17555 9435
rect 22066 9432 22094 9608
rect 22738 9596 22744 9608
rect 22796 9636 22802 9648
rect 23308 9636 23336 9676
rect 23474 9636 23480 9648
rect 22796 9608 23336 9636
rect 23435 9608 23480 9636
rect 22796 9596 22802 9608
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 23584 9636 23612 9676
rect 24780 9676 25084 9704
rect 24780 9636 24808 9676
rect 24946 9636 24952 9648
rect 23584 9608 24808 9636
rect 24907 9608 24952 9636
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 25056 9636 25084 9676
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 29181 9707 29239 9713
rect 29181 9704 29193 9707
rect 29144 9676 29193 9704
rect 29144 9664 29150 9676
rect 29181 9673 29193 9676
rect 29227 9673 29239 9707
rect 29181 9667 29239 9673
rect 27982 9636 27988 9648
rect 25056 9608 27988 9636
rect 27982 9596 27988 9608
rect 28040 9596 28046 9648
rect 22646 9568 22652 9580
rect 22607 9540 22652 9568
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 24854 9568 24860 9580
rect 24815 9540 24860 9568
rect 24854 9528 24860 9540
rect 24912 9528 24918 9580
rect 28902 9528 28908 9580
rect 28960 9568 28966 9580
rect 29365 9571 29423 9577
rect 29365 9568 29377 9571
rect 28960 9540 29377 9568
rect 28960 9528 28966 9540
rect 29365 9537 29377 9540
rect 29411 9537 29423 9571
rect 37918 9568 37924 9580
rect 37879 9540 37924 9568
rect 29365 9531 29423 9537
rect 37918 9528 37924 9540
rect 37976 9528 37982 9580
rect 23385 9503 23443 9509
rect 23385 9469 23397 9503
rect 23431 9500 23443 9503
rect 25958 9500 25964 9512
rect 23431 9472 25964 9500
rect 23431 9469 23443 9472
rect 23385 9463 23443 9469
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 17543 9404 22094 9432
rect 23937 9435 23995 9441
rect 17543 9401 17555 9404
rect 17497 9395 17555 9401
rect 23937 9401 23949 9435
rect 23983 9432 23995 9435
rect 25866 9432 25872 9444
rect 23983 9404 25872 9432
rect 23983 9401 23995 9404
rect 23937 9395 23995 9401
rect 25866 9392 25872 9404
rect 25924 9392 25930 9444
rect 37274 9392 37280 9444
rect 37332 9432 37338 9444
rect 37737 9435 37795 9441
rect 37737 9432 37749 9435
rect 37332 9404 37749 9432
rect 37332 9392 37338 9404
rect 37737 9401 37749 9404
rect 37783 9401 37795 9435
rect 37737 9395 37795 9401
rect 9180 9336 16574 9364
rect 19705 9367 19763 9373
rect 9180 9324 9186 9336
rect 19705 9333 19717 9367
rect 19751 9364 19763 9367
rect 20346 9364 20352 9376
rect 19751 9336 20352 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 22741 9367 22799 9373
rect 22741 9333 22753 9367
rect 22787 9364 22799 9367
rect 26878 9364 26884 9376
rect 22787 9336 26884 9364
rect 22787 9333 22799 9336
rect 22741 9327 22799 9333
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 14918 9160 14924 9172
rect 14879 9132 14924 9160
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 20165 9163 20223 9169
rect 20165 9129 20177 9163
rect 20211 9160 20223 9163
rect 20530 9160 20536 9172
rect 20211 9132 20536 9160
rect 20211 9129 20223 9132
rect 20165 9123 20223 9129
rect 20530 9120 20536 9132
rect 20588 9120 20594 9172
rect 22373 9163 22431 9169
rect 22373 9129 22385 9163
rect 22419 9160 22431 9163
rect 22462 9160 22468 9172
rect 22419 9132 22468 9160
rect 22419 9129 22431 9132
rect 22373 9123 22431 9129
rect 22462 9120 22468 9132
rect 22520 9120 22526 9172
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 9024 14519 9027
rect 14642 9024 14648 9036
rect 14507 8996 14648 9024
rect 14507 8993 14519 8996
rect 14461 8987 14519 8993
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 25317 9027 25375 9033
rect 25317 8993 25329 9027
rect 25363 9024 25375 9027
rect 28350 9024 28356 9036
rect 25363 8996 28356 9024
rect 25363 8993 25375 8996
rect 25317 8987 25375 8993
rect 28350 8984 28356 8996
rect 28408 8984 28414 9036
rect 30558 9024 30564 9036
rect 30519 8996 30564 9024
rect 30558 8984 30564 8996
rect 30616 8984 30622 9036
rect 37550 9024 37556 9036
rect 37511 8996 37556 9024
rect 37550 8984 37556 8996
rect 37608 8984 37614 9036
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 12492 8928 14289 8956
rect 12492 8916 12498 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 20346 8956 20352 8968
rect 20307 8928 20352 8956
rect 14277 8919 14335 8925
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 22278 8956 22284 8968
rect 22239 8928 22284 8956
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22922 8956 22928 8968
rect 22883 8928 22928 8956
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 25498 8916 25504 8968
rect 25556 8956 25562 8968
rect 27157 8959 27215 8965
rect 27157 8956 27169 8959
rect 25556 8928 27169 8956
rect 25556 8916 25562 8928
rect 27157 8925 27169 8928
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 32398 8916 32404 8968
rect 32456 8956 32462 8968
rect 32953 8959 33011 8965
rect 32953 8956 32965 8959
rect 32456 8928 32965 8956
rect 32456 8916 32462 8928
rect 32953 8925 32965 8928
rect 32999 8925 33011 8959
rect 32953 8919 33011 8925
rect 23201 8891 23259 8897
rect 23201 8857 23213 8891
rect 23247 8888 23259 8891
rect 24673 8891 24731 8897
rect 24673 8888 24685 8891
rect 23247 8860 24685 8888
rect 23247 8857 23259 8860
rect 23201 8851 23259 8857
rect 24673 8857 24685 8860
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 24762 8848 24768 8900
rect 24820 8888 24826 8900
rect 30098 8888 30104 8900
rect 24820 8860 24865 8888
rect 30059 8860 30104 8888
rect 24820 8848 24826 8860
rect 30098 8848 30104 8860
rect 30156 8848 30162 8900
rect 30193 8891 30251 8897
rect 30193 8857 30205 8891
rect 30239 8888 30251 8891
rect 30282 8888 30288 8900
rect 30239 8860 30288 8888
rect 30239 8857 30251 8860
rect 30193 8851 30251 8857
rect 30282 8848 30288 8860
rect 30340 8848 30346 8900
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 27249 8823 27307 8829
rect 27249 8789 27261 8823
rect 27295 8820 27307 8823
rect 27706 8820 27712 8832
rect 27295 8792 27712 8820
rect 27295 8789 27307 8792
rect 27249 8783 27307 8789
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 32769 8823 32827 8829
rect 32769 8789 32781 8823
rect 32815 8820 32827 8823
rect 33594 8820 33600 8832
rect 32815 8792 33600 8820
rect 32815 8789 32827 8792
rect 32769 8783 32827 8789
rect 33594 8780 33600 8792
rect 33652 8780 33658 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 17402 8616 17408 8628
rect 10459 8588 17408 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 28902 8616 28908 8628
rect 28863 8588 28908 8616
rect 28902 8576 28908 8588
rect 28960 8576 28966 8628
rect 30098 8616 30104 8628
rect 30059 8588 30104 8616
rect 30098 8576 30104 8588
rect 30156 8576 30162 8628
rect 38102 8616 38108 8628
rect 38063 8588 38108 8616
rect 38102 8576 38108 8588
rect 38160 8576 38166 8628
rect 22186 8548 22192 8560
rect 22147 8520 22192 8548
rect 22186 8508 22192 8520
rect 22244 8508 22250 8560
rect 22738 8548 22744 8560
rect 22699 8520 22744 8548
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 27706 8548 27712 8560
rect 27667 8520 27712 8548
rect 27706 8508 27712 8520
rect 27764 8508 27770 8560
rect 28261 8551 28319 8557
rect 28261 8517 28273 8551
rect 28307 8548 28319 8551
rect 28350 8548 28356 8560
rect 28307 8520 28356 8548
rect 28307 8517 28319 8520
rect 28261 8511 28319 8517
rect 28350 8508 28356 8520
rect 28408 8508 28414 8560
rect 4614 8440 4620 8492
rect 4672 8480 4678 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 4672 8452 10333 8480
rect 4672 8440 4678 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 24854 8440 24860 8492
rect 24912 8480 24918 8492
rect 26421 8483 26479 8489
rect 26421 8480 26433 8483
rect 24912 8452 26433 8480
rect 24912 8440 24918 8452
rect 26421 8449 26433 8452
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8480 29147 8483
rect 29362 8480 29368 8492
rect 29135 8452 29368 8480
rect 29135 8449 29147 8452
rect 29089 8443 29147 8449
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 22097 8415 22155 8421
rect 22097 8412 22109 8415
rect 21315 8384 22109 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 22097 8381 22109 8384
rect 22143 8381 22155 8415
rect 22097 8375 22155 8381
rect 26436 8344 26464 8443
rect 27617 8415 27675 8421
rect 27617 8381 27629 8415
rect 27663 8412 27675 8415
rect 27706 8412 27712 8424
rect 27663 8384 27712 8412
rect 27663 8381 27675 8384
rect 27617 8375 27675 8381
rect 27706 8372 27712 8384
rect 27764 8372 27770 8424
rect 29104 8344 29132 8443
rect 29362 8440 29368 8452
rect 29420 8440 29426 8492
rect 38286 8480 38292 8492
rect 38247 8452 38292 8480
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 26436 8316 29132 8344
rect 26510 8276 26516 8288
rect 26471 8248 26516 8276
rect 26510 8236 26516 8248
rect 26568 8236 26574 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 8018 8072 8024 8084
rect 1627 8044 8024 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 9122 8072 9128 8084
rect 8343 8044 9128 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 31849 8075 31907 8081
rect 31849 8072 31861 8075
rect 11572 8044 31861 8072
rect 11572 8032 11578 8044
rect 31849 8041 31861 8044
rect 31895 8072 31907 8075
rect 32398 8072 32404 8084
rect 31895 8044 32404 8072
rect 31895 8041 31907 8044
rect 31849 8035 31907 8041
rect 32398 8032 32404 8044
rect 32456 8032 32462 8084
rect 27706 8004 27712 8016
rect 27667 7976 27712 8004
rect 27706 7964 27712 7976
rect 27764 7964 27770 8016
rect 31573 8007 31631 8013
rect 31573 7973 31585 8007
rect 31619 8004 31631 8007
rect 38378 8004 38384 8016
rect 31619 7976 38384 8004
rect 31619 7973 31631 7976
rect 31573 7967 31631 7973
rect 38378 7964 38384 7976
rect 38436 7964 38442 8016
rect 23198 7896 23204 7948
rect 23256 7936 23262 7948
rect 37737 7939 37795 7945
rect 37737 7936 37749 7939
rect 23256 7908 37749 7936
rect 23256 7896 23262 7908
rect 37737 7905 37749 7908
rect 37783 7905 37795 7939
rect 37737 7899 37795 7905
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21729 7871 21787 7877
rect 21729 7868 21741 7871
rect 21048 7840 21741 7868
rect 21048 7828 21054 7840
rect 21729 7837 21741 7840
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 21821 7871 21879 7877
rect 21821 7837 21833 7871
rect 21867 7868 21879 7871
rect 23385 7871 23443 7877
rect 23385 7868 23397 7871
rect 21867 7840 23397 7868
rect 21867 7837 21879 7840
rect 21821 7831 21879 7837
rect 23385 7837 23397 7840
rect 23431 7837 23443 7871
rect 23385 7831 23443 7837
rect 27154 7828 27160 7880
rect 27212 7868 27218 7880
rect 27709 7871 27767 7877
rect 27709 7868 27721 7871
rect 27212 7840 27721 7868
rect 27212 7828 27218 7840
rect 27709 7837 27721 7840
rect 27755 7837 27767 7871
rect 32398 7868 32404 7880
rect 32359 7840 32404 7868
rect 27709 7831 27767 7837
rect 32398 7828 32404 7840
rect 32456 7828 32462 7880
rect 37458 7868 37464 7880
rect 37419 7840 37464 7868
rect 37458 7828 37464 7840
rect 37516 7828 37522 7880
rect 31386 7800 31392 7812
rect 31347 7772 31392 7800
rect 31386 7760 31392 7772
rect 31444 7760 31450 7812
rect 23201 7735 23259 7741
rect 23201 7701 23213 7735
rect 23247 7732 23259 7735
rect 27798 7732 27804 7744
rect 23247 7704 27804 7732
rect 23247 7701 23259 7704
rect 23201 7695 23259 7701
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 32217 7735 32275 7741
rect 32217 7701 32229 7735
rect 32263 7732 32275 7735
rect 34330 7732 34336 7744
rect 32263 7704 34336 7732
rect 32263 7701 32275 7704
rect 32217 7695 32275 7701
rect 34330 7692 34336 7704
rect 34388 7692 34394 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 26602 7528 26608 7540
rect 26563 7500 26608 7528
rect 26602 7488 26608 7500
rect 26660 7488 26666 7540
rect 37734 7488 37740 7540
rect 37792 7528 37798 7540
rect 38105 7531 38163 7537
rect 38105 7528 38117 7531
rect 37792 7500 38117 7528
rect 37792 7488 37798 7500
rect 38105 7497 38117 7500
rect 38151 7497 38163 7531
rect 38105 7491 38163 7497
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 22278 7392 22284 7404
rect 20487 7364 22284 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 22278 7352 22284 7364
rect 22336 7392 22342 7404
rect 23198 7392 23204 7404
rect 22336 7364 23204 7392
rect 22336 7352 22342 7364
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7392 23811 7395
rect 24854 7392 24860 7404
rect 23799 7364 24860 7392
rect 23799 7361 23811 7364
rect 23753 7355 23811 7361
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 25958 7392 25964 7404
rect 25919 7364 25964 7392
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 26145 7395 26203 7401
rect 26145 7361 26157 7395
rect 26191 7392 26203 7395
rect 26510 7392 26516 7404
rect 26191 7364 26516 7392
rect 26191 7361 26203 7364
rect 26145 7355 26203 7361
rect 26510 7352 26516 7364
rect 26568 7352 26574 7404
rect 38286 7392 38292 7404
rect 38247 7364 38292 7392
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 6546 7216 6552 7268
rect 6604 7256 6610 7268
rect 6604 7228 16574 7256
rect 6604 7216 6610 7228
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 9122 7188 9128 7200
rect 1627 7160 9128 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 16546 7188 16574 7228
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 16546 7160 20269 7188
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 20257 7151 20315 7157
rect 23569 7191 23627 7197
rect 23569 7157 23581 7191
rect 23615 7188 23627 7191
rect 24762 7188 24768 7200
rect 23615 7160 24768 7188
rect 23615 7157 23627 7160
rect 23569 7151 23627 7157
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 12434 6848 12440 6860
rect 9263 6820 12440 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 24029 6851 24087 6857
rect 24029 6817 24041 6851
rect 24075 6848 24087 6851
rect 26602 6848 26608 6860
rect 24075 6820 26608 6848
rect 24075 6817 24087 6820
rect 24029 6811 24087 6817
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 30558 6848 30564 6860
rect 29748 6820 30564 6848
rect 9122 6780 9128 6792
rect 9083 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 23382 6780 23388 6792
rect 23343 6752 23388 6780
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6780 23627 6783
rect 24762 6780 24768 6792
rect 23615 6752 24624 6780
rect 24723 6752 24768 6780
rect 23615 6749 23627 6752
rect 23569 6743 23627 6749
rect 24596 6653 24624 6752
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 29748 6789 29776 6820
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 31481 6851 31539 6857
rect 31481 6817 31493 6851
rect 31527 6848 31539 6851
rect 31662 6848 31668 6860
rect 31527 6820 31668 6848
rect 31527 6817 31539 6820
rect 31481 6811 31539 6817
rect 31662 6808 31668 6820
rect 31720 6808 31726 6860
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 30466 6712 30472 6724
rect 30427 6684 30472 6712
rect 30466 6672 30472 6684
rect 30524 6672 30530 6724
rect 30561 6715 30619 6721
rect 30561 6681 30573 6715
rect 30607 6712 30619 6715
rect 30834 6712 30840 6724
rect 30607 6684 30840 6712
rect 30607 6681 30619 6684
rect 30561 6675 30619 6681
rect 30834 6672 30840 6684
rect 30892 6672 30898 6724
rect 24581 6647 24639 6653
rect 24581 6613 24593 6647
rect 24627 6613 24639 6647
rect 29822 6644 29828 6656
rect 29783 6616 29828 6644
rect 24581 6607 24639 6613
rect 29822 6604 29828 6616
rect 29880 6604 29886 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 12434 6264 12440 6316
rect 12492 6304 12498 6316
rect 14921 6307 14979 6313
rect 14921 6304 14933 6307
rect 12492 6276 14933 6304
rect 12492 6264 12498 6276
rect 14921 6273 14933 6276
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 24489 6307 24547 6313
rect 24489 6304 24501 6307
rect 23348 6276 24501 6304
rect 23348 6264 23354 6276
rect 24489 6273 24501 6276
rect 24535 6273 24547 6307
rect 24489 6267 24547 6273
rect 29822 6264 29828 6316
rect 29880 6304 29886 6316
rect 30469 6307 30527 6313
rect 30469 6304 30481 6307
rect 29880 6276 30481 6304
rect 29880 6264 29886 6276
rect 30469 6273 30481 6276
rect 30515 6273 30527 6307
rect 30469 6267 30527 6273
rect 15013 6103 15071 6109
rect 15013 6069 15025 6103
rect 15059 6100 15071 6103
rect 23382 6100 23388 6112
rect 15059 6072 23388 6100
rect 15059 6069 15071 6072
rect 15013 6063 15071 6069
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 24581 6103 24639 6109
rect 24581 6069 24593 6103
rect 24627 6100 24639 6103
rect 26326 6100 26332 6112
rect 24627 6072 26332 6100
rect 24627 6069 24639 6072
rect 24581 6063 24639 6069
rect 26326 6060 26332 6072
rect 26384 6060 26390 6112
rect 30285 6103 30343 6109
rect 30285 6069 30297 6103
rect 30331 6100 30343 6103
rect 31662 6100 31668 6112
rect 30331 6072 31668 6100
rect 30331 6069 30343 6072
rect 30285 6063 30343 6069
rect 31662 6060 31668 6072
rect 31720 6060 31726 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1544 5868 1593 5896
rect 1544 5856 1550 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 26326 5692 26332 5704
rect 26287 5664 26332 5692
rect 26326 5652 26332 5664
rect 26384 5652 26390 5704
rect 38013 5695 38071 5701
rect 38013 5661 38025 5695
rect 38059 5661 38071 5695
rect 38013 5655 38071 5661
rect 13998 5584 14004 5636
rect 14056 5624 14062 5636
rect 37645 5627 37703 5633
rect 37645 5624 37657 5627
rect 14056 5596 37657 5624
rect 14056 5584 14062 5596
rect 37645 5593 37657 5596
rect 37691 5624 37703 5627
rect 38028 5624 38056 5655
rect 37691 5596 38056 5624
rect 37691 5593 37703 5596
rect 37645 5587 37703 5593
rect 26145 5559 26203 5565
rect 26145 5525 26157 5559
rect 26191 5556 26203 5559
rect 28902 5556 28908 5568
rect 26191 5528 28908 5556
rect 26191 5525 26203 5528
rect 26145 5519 26203 5525
rect 28902 5516 28908 5528
rect 28960 5516 28966 5568
rect 38194 5556 38200 5568
rect 38155 5528 38200 5556
rect 38194 5516 38200 5528
rect 38252 5516 38258 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 22649 5355 22707 5361
rect 22649 5352 22661 5355
rect 18748 5324 22661 5352
rect 18748 5312 18754 5324
rect 22649 5321 22661 5324
rect 22695 5321 22707 5355
rect 22649 5315 22707 5321
rect 23937 5355 23995 5361
rect 23937 5321 23949 5355
rect 23983 5352 23995 5355
rect 25958 5352 25964 5364
rect 23983 5324 25964 5352
rect 23983 5321 23995 5324
rect 23937 5315 23995 5321
rect 25958 5312 25964 5324
rect 26016 5312 26022 5364
rect 29457 5355 29515 5361
rect 29457 5321 29469 5355
rect 29503 5352 29515 5355
rect 30466 5352 30472 5364
rect 29503 5324 30472 5352
rect 29503 5321 29515 5324
rect 29457 5315 29515 5321
rect 30466 5312 30472 5324
rect 30524 5312 30530 5364
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5216 22615 5219
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 22603 5188 23857 5216
rect 22603 5185 22615 5188
rect 22557 5179 22615 5185
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 23860 5148 23888 5179
rect 27614 5176 27620 5228
rect 27672 5216 27678 5228
rect 29365 5219 29423 5225
rect 29365 5216 29377 5219
rect 27672 5188 29377 5216
rect 27672 5176 27678 5188
rect 29365 5185 29377 5188
rect 29411 5185 29423 5219
rect 29365 5179 29423 5185
rect 37734 5148 37740 5160
rect 23860 5120 37740 5148
rect 37734 5108 37740 5120
rect 37792 5108 37798 5160
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 37734 4672 37740 4684
rect 37695 4644 37740 4672
rect 37734 4632 37740 4644
rect 37792 4632 37798 4684
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 2225 4607 2283 4613
rect 2225 4604 2237 4607
rect 1627 4576 2237 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 2225 4573 2237 4576
rect 2271 4604 2283 4607
rect 36722 4604 36728 4616
rect 2271 4576 36728 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 36722 4564 36728 4576
rect 36780 4564 36786 4616
rect 37458 4604 37464 4616
rect 37419 4576 37464 4604
rect 37458 4564 37464 4576
rect 37516 4564 37522 4616
rect 1762 4468 1768 4480
rect 1723 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 36722 4088 36728 4140
rect 36780 4128 36786 4140
rect 38013 4131 38071 4137
rect 38013 4128 38025 4131
rect 36780 4100 38025 4128
rect 36780 4088 36786 4100
rect 38013 4097 38025 4100
rect 38059 4097 38071 4131
rect 38013 4091 38071 4097
rect 35894 3884 35900 3936
rect 35952 3924 35958 3936
rect 37829 3927 37887 3933
rect 37829 3924 37841 3927
rect 35952 3896 37841 3924
rect 35952 3884 35958 3896
rect 37829 3893 37841 3896
rect 37875 3893 37887 3927
rect 37829 3887 37887 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 36722 3720 36728 3732
rect 36683 3692 36728 3720
rect 36722 3680 36728 3692
rect 36780 3680 36786 3732
rect 37734 3584 37740 3596
rect 36924 3556 37740 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1854 3516 1860 3528
rect 1627 3488 1860 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 36924 3525 36952 3556
rect 37734 3544 37740 3556
rect 37792 3544 37798 3596
rect 36909 3519 36967 3525
rect 36909 3485 36921 3519
rect 36955 3485 36967 3519
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 36909 3479 36967 3485
rect 37016 3488 37565 3516
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 37016 3448 37044 3488
rect 37553 3485 37565 3488
rect 37599 3485 37611 3519
rect 37553 3479 37611 3485
rect 38013 3519 38071 3525
rect 38013 3485 38025 3519
rect 38059 3485 38071 3519
rect 38013 3479 38071 3485
rect 38028 3448 38056 3479
rect 36044 3420 37044 3448
rect 37384 3420 38056 3448
rect 36044 3408 36050 3420
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 37384 3389 37412 3420
rect 37369 3383 37427 3389
rect 37369 3349 37381 3383
rect 37415 3349 37427 3383
rect 38194 3380 38200 3392
rect 38155 3352 38200 3380
rect 37369 3343 37427 3349
rect 38194 3340 38200 3352
rect 38252 3340 38258 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3418 3176 3424 3188
rect 2363 3148 3424 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 3973 3179 4031 3185
rect 3973 3145 3985 3179
rect 4019 3176 4031 3179
rect 4614 3176 4620 3188
rect 4019 3148 4620 3176
rect 4019 3145 4031 3148
rect 3973 3139 4031 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 22649 3179 22707 3185
rect 22649 3145 22661 3179
rect 22695 3176 22707 3179
rect 22922 3176 22928 3188
rect 22695 3148 22928 3176
rect 22695 3145 22707 3148
rect 22649 3139 22707 3145
rect 22922 3136 22928 3148
rect 22980 3136 22986 3188
rect 35253 3179 35311 3185
rect 35253 3145 35265 3179
rect 35299 3176 35311 3179
rect 36446 3176 36452 3188
rect 35299 3148 36452 3176
rect 35299 3145 35311 3148
rect 35253 3139 35311 3145
rect 36446 3136 36452 3148
rect 36504 3136 36510 3188
rect 21634 3068 21640 3120
rect 21692 3108 21698 3120
rect 21692 3080 38056 3108
rect 21692 3068 21698 3080
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2774 3040 2780 3052
rect 2547 3012 2780 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 1596 2972 1624 3003
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2924 3012 3157 3040
rect 2924 3000 2930 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3936 3012 4169 3040
rect 3936 3000 3942 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 8202 3040 8208 3052
rect 5583 3012 8208 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13265 3043 13323 3049
rect 13265 3040 13277 3043
rect 13044 3012 13277 3040
rect 13044 3000 13050 3012
rect 13265 3009 13277 3012
rect 13311 3009 13323 3043
rect 13265 3003 13323 3009
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16816 3012 17049 3040
rect 16816 3000 16822 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 22833 3043 22891 3049
rect 22833 3040 22845 3043
rect 22612 3012 22845 3040
rect 22612 3000 22618 3012
rect 22833 3009 22845 3012
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 30377 3043 30435 3049
rect 30377 3040 30389 3043
rect 28960 3012 30389 3040
rect 28960 3000 28966 3012
rect 30377 3009 30389 3012
rect 30423 3009 30435 3043
rect 35434 3040 35440 3052
rect 35395 3012 35440 3040
rect 30377 3003 30435 3009
rect 35434 3000 35440 3012
rect 35492 3000 35498 3052
rect 35897 3043 35955 3049
rect 35897 3009 35909 3043
rect 35943 3009 35955 3043
rect 35897 3003 35955 3009
rect 31386 2972 31392 2984
rect 1596 2944 13124 2972
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2904 3019 2907
rect 9030 2904 9036 2916
rect 3007 2876 9036 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 13096 2913 13124 2944
rect 22066 2944 31392 2972
rect 13081 2907 13139 2913
rect 13081 2873 13093 2907
rect 13127 2873 13139 2907
rect 13081 2867 13139 2873
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 22066 2904 22094 2944
rect 31386 2932 31392 2944
rect 31444 2932 31450 2984
rect 31570 2932 31576 2984
rect 31628 2972 31634 2984
rect 35912 2972 35940 3003
rect 35986 3000 35992 3052
rect 36044 3040 36050 3052
rect 36909 3043 36967 3049
rect 36044 3012 36089 3040
rect 36044 3000 36050 3012
rect 36909 3009 36921 3043
rect 36955 3040 36967 3043
rect 37366 3040 37372 3052
rect 36955 3012 37372 3040
rect 36955 3009 36967 3012
rect 36909 3003 36967 3009
rect 37366 3000 37372 3012
rect 37424 3000 37430 3052
rect 38028 3049 38056 3080
rect 38013 3043 38071 3049
rect 38013 3009 38025 3043
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 31628 2944 35940 2972
rect 31628 2932 31634 2944
rect 16899 2876 22094 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 30374 2864 30380 2916
rect 30432 2904 30438 2916
rect 36725 2907 36783 2913
rect 36725 2904 36737 2907
rect 30432 2876 36737 2904
rect 30432 2864 30438 2876
rect 36725 2873 36737 2876
rect 36771 2873 36783 2907
rect 36725 2867 36783 2873
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1765 2839 1823 2845
rect 1765 2836 1777 2839
rect 716 2808 1777 2836
rect 716 2796 722 2808
rect 1765 2805 1777 2808
rect 1811 2805 1823 2839
rect 5350 2836 5356 2848
rect 5311 2808 5356 2836
rect 1765 2799 1823 2805
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 30561 2839 30619 2845
rect 30561 2836 30573 2839
rect 30340 2808 30573 2836
rect 30340 2796 30346 2808
rect 30561 2805 30573 2808
rect 30607 2805 30619 2839
rect 30561 2799 30619 2805
rect 38197 2839 38255 2845
rect 38197 2805 38209 2839
rect 38243 2836 38255 2839
rect 38654 2836 38660 2848
rect 38243 2808 38660 2836
rect 38243 2805 38255 2808
rect 38197 2799 38255 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 8260 2604 10425 2632
rect 8260 2592 8266 2604
rect 10413 2601 10425 2604
rect 10459 2601 10471 2635
rect 10413 2595 10471 2601
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 12526 2632 12532 2644
rect 11747 2604 12532 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13170 2632 13176 2644
rect 12636 2604 13176 2632
rect 14 2524 20 2576
rect 72 2564 78 2576
rect 2961 2567 3019 2573
rect 2961 2564 2973 2567
rect 72 2536 2973 2564
rect 72 2524 78 2536
rect 2961 2533 2973 2536
rect 3007 2533 3019 2567
rect 2961 2527 3019 2533
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 9769 2567 9827 2573
rect 9769 2533 9781 2567
rect 9815 2564 9827 2567
rect 12636 2564 12664 2604
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 20254 2632 20260 2644
rect 19536 2604 20260 2632
rect 19536 2564 19564 2604
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22094 2632 22100 2644
rect 22051 2604 22100 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 24581 2635 24639 2641
rect 24581 2601 24593 2635
rect 24627 2632 24639 2635
rect 24670 2632 24676 2644
rect 24627 2604 24676 2632
rect 24627 2601 24639 2604
rect 24581 2595 24639 2601
rect 24670 2592 24676 2604
rect 24728 2592 24734 2644
rect 27154 2632 27160 2644
rect 27115 2604 27160 2632
rect 27154 2592 27160 2604
rect 27212 2592 27218 2644
rect 9815 2536 12664 2564
rect 13188 2536 19564 2564
rect 20073 2567 20131 2573
rect 9815 2533 9827 2536
rect 9769 2527 9827 2533
rect 5350 2496 5356 2508
rect 2792 2468 5356 2496
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2792 2437 2820 2468
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 7300 2496 7328 2527
rect 12158 2496 12164 2508
rect 7300 2468 12164 2496
rect 12158 2456 12164 2468
rect 12216 2456 12222 2508
rect 13188 2505 13216 2536
rect 20073 2533 20085 2567
rect 20119 2564 20131 2567
rect 22646 2564 22652 2576
rect 20119 2536 22652 2564
rect 20119 2533 20131 2536
rect 20073 2527 20131 2533
rect 22646 2524 22652 2536
rect 22704 2524 22710 2576
rect 26206 2536 37504 2564
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 15197 2499 15255 2505
rect 15197 2465 15209 2499
rect 15243 2496 15255 2499
rect 16666 2496 16672 2508
rect 15243 2468 16672 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 26206 2496 26234 2536
rect 31202 2496 31208 2508
rect 21192 2468 26234 2496
rect 31163 2468 31208 2496
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 2004 2400 2053 2428
rect 2004 2388 2010 2400
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2397 2835 2431
rect 3970 2428 3976 2440
rect 3931 2400 3976 2428
rect 2777 2391 2835 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4120 2400 5273 2428
rect 4120 2388 4126 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 6546 2428 6552 2440
rect 6507 2400 6552 2428
rect 5261 2391 5319 2397
rect 6546 2388 6552 2400
rect 6604 2388 6610 2440
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7156 2400 7481 2428
rect 7156 2388 7162 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 9309 2431 9367 2437
rect 9309 2428 9321 2431
rect 8444 2400 9321 2428
rect 8444 2388 8450 2400
rect 9309 2397 9321 2400
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11885 2431 11943 2437
rect 11885 2428 11897 2431
rect 11664 2400 11897 2428
rect 11664 2388 11670 2400
rect 11885 2397 11897 2400
rect 11931 2397 11943 2431
rect 12894 2428 12900 2440
rect 12855 2400 12900 2428
rect 11885 2391 11943 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 13596 2400 14473 2428
rect 13596 2388 13602 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 14884 2400 14933 2428
rect 14884 2388 14890 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16172 2400 16865 2428
rect 16172 2388 16178 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18104 2400 18337 2428
rect 18104 2388 18110 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20036 2400 20269 2428
rect 20036 2388 20042 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 13354 2320 13360 2372
rect 13412 2360 13418 2372
rect 21192 2360 21220 2468
rect 31202 2456 31208 2468
rect 31260 2456 31266 2508
rect 32030 2456 32036 2508
rect 32088 2496 32094 2508
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 32088 2468 32597 2496
rect 32088 2456 32094 2468
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 34330 2456 34336 2508
rect 34388 2496 34394 2508
rect 34388 2468 36676 2496
rect 34388 2456 34394 2468
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21324 2400 22201 2428
rect 21324 2388 21330 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 23198 2428 23204 2440
rect 23159 2400 23204 2428
rect 22189 2391 22247 2397
rect 23198 2388 23204 2400
rect 23256 2388 23262 2440
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 13412 2332 21220 2360
rect 13412 2320 13418 2332
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2225 2295 2283 2301
rect 2225 2292 2237 2295
rect 2004 2264 2237 2292
rect 2004 2252 2010 2264
rect 2225 2261 2237 2264
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 3234 2252 3240 2304
rect 3292 2292 3298 2304
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3292 2264 4169 2292
rect 3292 2252 3298 2264
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5224 2264 5457 2292
rect 5224 2252 5230 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5445 2255 5503 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 12434 2292 12440 2304
rect 9171 2264 12440 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12986 2252 12992 2304
rect 13044 2292 13050 2304
rect 23492 2292 23520 2391
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24765 2431 24823 2437
rect 24765 2428 24777 2431
rect 24544 2400 24777 2428
rect 24544 2388 24550 2400
rect 24765 2397 24777 2400
rect 24811 2397 24823 2431
rect 24765 2391 24823 2397
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25832 2400 26065 2428
rect 25832 2388 25838 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 26053 2391 26111 2397
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27798 2428 27804 2440
rect 27759 2400 27804 2428
rect 27341 2391 27399 2397
rect 27798 2388 27804 2400
rect 27856 2388 27862 2440
rect 29730 2428 29736 2440
rect 29691 2400 29736 2428
rect 29730 2388 29736 2400
rect 29788 2388 29794 2440
rect 30926 2428 30932 2440
rect 30887 2400 30932 2428
rect 30926 2388 30932 2400
rect 30984 2388 30990 2440
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 33594 2428 33600 2440
rect 33555 2400 33600 2428
rect 32309 2391 32367 2397
rect 33594 2388 33600 2400
rect 33652 2388 33658 2440
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 31662 2320 31668 2372
rect 31720 2360 31726 2372
rect 34900 2360 34928 2391
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36648 2437 36676 2468
rect 37476 2437 37504 2536
rect 36633 2431 36691 2437
rect 35952 2400 35997 2428
rect 35952 2388 35958 2400
rect 36633 2397 36645 2431
rect 36679 2397 36691 2431
rect 36633 2391 36691 2397
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2428 37519 2431
rect 38013 2431 38071 2437
rect 38013 2428 38025 2431
rect 37507 2400 38025 2428
rect 37507 2397 37519 2400
rect 37461 2391 37519 2397
rect 38013 2397 38025 2400
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 37182 2360 37188 2372
rect 31720 2332 34928 2360
rect 36096 2332 37188 2360
rect 31720 2320 31726 2332
rect 13044 2264 23520 2292
rect 25869 2295 25927 2301
rect 13044 2252 13050 2264
rect 25869 2261 25881 2295
rect 25915 2292 25927 2295
rect 27614 2292 27620 2304
rect 25915 2264 27620 2292
rect 25915 2261 25927 2264
rect 25869 2255 25927 2261
rect 27614 2252 27620 2264
rect 27672 2252 27678 2304
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 27985 2295 28043 2301
rect 27985 2292 27997 2295
rect 27764 2264 27997 2292
rect 27764 2252 27770 2264
rect 27985 2261 27997 2264
rect 28031 2261 28043 2295
rect 27985 2255 28043 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 29052 2264 29929 2292
rect 29052 2252 29058 2264
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33781 2295 33839 2301
rect 33781 2292 33793 2295
rect 33560 2264 33793 2292
rect 33560 2252 33566 2264
rect 33781 2261 33793 2264
rect 33827 2261 33839 2295
rect 33781 2255 33839 2261
rect 34146 2252 34152 2304
rect 34204 2292 34210 2304
rect 36096 2301 36124 2332
rect 37182 2320 37188 2332
rect 37240 2320 37246 2372
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34204 2264 35081 2292
rect 34204 2252 34210 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 36081 2295 36139 2301
rect 36081 2261 36093 2295
rect 36127 2261 36139 2295
rect 36814 2292 36820 2304
rect 36775 2264 36820 2292
rect 36081 2255 36139 2261
rect 36814 2252 36820 2264
rect 36872 2252 36878 2304
rect 37090 2252 37096 2304
rect 37148 2292 37154 2304
rect 37645 2295 37703 2301
rect 37645 2292 37657 2295
rect 37148 2264 37657 2292
rect 37148 2252 37154 2264
rect 37645 2261 37657 2264
rect 37691 2261 37703 2295
rect 37645 2255 37703 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 2872 38292 2924 38344
rect 4620 38292 4672 38344
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 14740 37408 14792 37460
rect 17776 37408 17828 37460
rect 30932 37408 30984 37460
rect 1952 37272 2004 37324
rect 4896 37272 4948 37324
rect 8392 37272 8444 37324
rect 17868 37340 17920 37392
rect 18144 37340 18196 37392
rect 18972 37340 19024 37392
rect 28172 37340 28224 37392
rect 2136 37204 2188 37256
rect 3424 37204 3476 37256
rect 5172 37204 5224 37256
rect 5816 37204 5868 37256
rect 7104 37204 7156 37256
rect 9036 37204 9088 37256
rect 9496 37204 9548 37256
rect 8116 37136 8168 37188
rect 10048 37136 10100 37188
rect 6368 37068 6420 37120
rect 6644 37068 6696 37120
rect 7196 37111 7248 37120
rect 7196 37077 7205 37111
rect 7205 37077 7239 37111
rect 7239 37077 7248 37111
rect 7196 37068 7248 37077
rect 9128 37068 9180 37120
rect 9772 37068 9824 37120
rect 11060 37136 11112 37188
rect 12256 37204 12308 37256
rect 13636 37204 13688 37256
rect 13820 37204 13872 37256
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 15292 37204 15344 37256
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 10324 37068 10376 37120
rect 11336 37068 11388 37120
rect 15936 37136 15988 37188
rect 18236 37204 18288 37256
rect 22744 37272 22796 37324
rect 25780 37315 25832 37324
rect 25780 37281 25789 37315
rect 25789 37281 25823 37315
rect 25823 37281 25832 37315
rect 25780 37272 25832 37281
rect 20536 37204 20588 37256
rect 22560 37204 22612 37256
rect 23480 37247 23532 37256
rect 23480 37213 23489 37247
rect 23489 37213 23523 37247
rect 23523 37213 23532 37247
rect 23480 37204 23532 37213
rect 24492 37204 24544 37256
rect 26056 37247 26108 37256
rect 26056 37213 26065 37247
rect 26065 37213 26099 37247
rect 26099 37213 26108 37247
rect 26056 37204 26108 37213
rect 18328 37136 18380 37188
rect 18880 37136 18932 37188
rect 14924 37068 14976 37120
rect 15016 37111 15068 37120
rect 15016 37077 15025 37111
rect 15025 37077 15059 37111
rect 15059 37077 15068 37111
rect 15016 37068 15068 37077
rect 16120 37068 16172 37120
rect 16764 37068 16816 37120
rect 19340 37068 19392 37120
rect 19984 37068 20036 37120
rect 21272 37068 21324 37120
rect 23204 37068 23256 37120
rect 26424 37068 26476 37120
rect 27712 37204 27764 37256
rect 28080 37247 28132 37256
rect 28080 37213 28089 37247
rect 28089 37213 28123 37247
rect 28123 37213 28132 37247
rect 29092 37272 29144 37324
rect 28080 37204 28132 37213
rect 27528 37136 27580 37188
rect 31300 37204 31352 37256
rect 31576 37204 31628 37256
rect 32956 37204 33008 37256
rect 30380 37136 30432 37188
rect 30472 37068 30524 37120
rect 30748 37136 30800 37188
rect 31668 37068 31720 37120
rect 33508 37136 33560 37188
rect 38660 37272 38712 37324
rect 33692 37204 33744 37256
rect 36176 37247 36228 37256
rect 36176 37213 36185 37247
rect 36185 37213 36219 37247
rect 36219 37213 36228 37247
rect 36176 37204 36228 37213
rect 33140 37068 33192 37120
rect 34520 37068 34572 37120
rect 36084 37068 36136 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 2228 36796 2280 36848
rect 9772 36796 9824 36848
rect 9864 36796 9916 36848
rect 2780 36728 2832 36780
rect 4160 36771 4212 36780
rect 4160 36737 4169 36771
rect 4169 36737 4203 36771
rect 4203 36737 4212 36771
rect 4160 36728 4212 36737
rect 7196 36728 7248 36780
rect 8116 36728 8168 36780
rect 8484 36728 8536 36780
rect 8668 36771 8720 36780
rect 8668 36737 8677 36771
rect 8677 36737 8711 36771
rect 8711 36737 8720 36771
rect 8668 36728 8720 36737
rect 9680 36728 9732 36780
rect 11612 36796 11664 36848
rect 10600 36771 10652 36780
rect 10600 36737 10609 36771
rect 10609 36737 10643 36771
rect 10643 36737 10652 36771
rect 10600 36728 10652 36737
rect 12624 36728 12676 36780
rect 11060 36660 11112 36712
rect 1584 36592 1636 36644
rect 8024 36635 8076 36644
rect 2780 36524 2832 36576
rect 8024 36601 8033 36635
rect 8033 36601 8067 36635
rect 8067 36601 8076 36635
rect 8024 36592 8076 36601
rect 11980 36592 12032 36644
rect 12164 36660 12216 36712
rect 13636 36660 13688 36712
rect 14924 36864 14976 36916
rect 17776 36864 17828 36916
rect 18052 36864 18104 36916
rect 15660 36796 15712 36848
rect 17868 36796 17920 36848
rect 18420 36796 18472 36848
rect 15752 36771 15804 36780
rect 15752 36737 15761 36771
rect 15761 36737 15795 36771
rect 15795 36737 15804 36771
rect 15752 36728 15804 36737
rect 12256 36592 12308 36644
rect 12992 36592 13044 36644
rect 9312 36524 9364 36576
rect 9404 36567 9456 36576
rect 9404 36533 9413 36567
rect 9413 36533 9447 36567
rect 9447 36533 9456 36567
rect 9404 36524 9456 36533
rect 10508 36524 10560 36576
rect 11428 36524 11480 36576
rect 11612 36524 11664 36576
rect 13176 36524 13228 36576
rect 14372 36592 14424 36644
rect 16856 36660 16908 36712
rect 24676 36796 24728 36848
rect 26608 36864 26660 36916
rect 25504 36796 25556 36848
rect 22560 36703 22612 36712
rect 22560 36669 22569 36703
rect 22569 36669 22603 36703
rect 22603 36669 22612 36703
rect 22560 36660 22612 36669
rect 24768 36703 24820 36712
rect 24768 36669 24777 36703
rect 24777 36669 24811 36703
rect 24811 36669 24820 36703
rect 24768 36660 24820 36669
rect 28264 36796 28316 36848
rect 29644 36864 29696 36916
rect 30380 36796 30432 36848
rect 30564 36796 30616 36848
rect 31668 36864 31720 36916
rect 32496 36864 32548 36916
rect 37372 36864 37424 36916
rect 32220 36796 32272 36848
rect 34060 36796 34112 36848
rect 36544 36796 36596 36848
rect 36728 36839 36780 36848
rect 36728 36805 36737 36839
rect 36737 36805 36771 36839
rect 36771 36805 36780 36839
rect 36728 36796 36780 36805
rect 37464 36771 37516 36780
rect 37464 36737 37473 36771
rect 37473 36737 37507 36771
rect 37507 36737 37516 36771
rect 37464 36728 37516 36737
rect 23940 36592 23992 36644
rect 24584 36592 24636 36644
rect 27160 36660 27212 36712
rect 27528 36703 27580 36712
rect 27528 36669 27537 36703
rect 27537 36669 27571 36703
rect 27571 36669 27580 36703
rect 27528 36660 27580 36669
rect 27804 36703 27856 36712
rect 27804 36669 27813 36703
rect 27813 36669 27847 36703
rect 27847 36669 27856 36703
rect 27804 36660 27856 36669
rect 29828 36703 29880 36712
rect 29828 36669 29837 36703
rect 29837 36669 29871 36703
rect 29871 36669 29880 36703
rect 29828 36660 29880 36669
rect 28816 36592 28868 36644
rect 19432 36567 19484 36576
rect 19432 36533 19441 36567
rect 19441 36533 19475 36567
rect 19475 36533 19484 36567
rect 19432 36524 19484 36533
rect 20260 36524 20312 36576
rect 25136 36524 25188 36576
rect 25228 36524 25280 36576
rect 29092 36524 29144 36576
rect 29828 36524 29880 36576
rect 33140 36592 33192 36644
rect 31300 36524 31352 36576
rect 32312 36567 32364 36576
rect 32312 36533 32321 36567
rect 32321 36533 32355 36567
rect 32355 36533 32364 36567
rect 32312 36524 32364 36533
rect 32404 36524 32456 36576
rect 35900 36567 35952 36576
rect 35900 36533 35909 36567
rect 35909 36533 35943 36567
rect 35943 36533 35952 36567
rect 35900 36524 35952 36533
rect 36084 36524 36136 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 8484 36363 8536 36372
rect 8484 36329 8493 36363
rect 8493 36329 8527 36363
rect 8527 36329 8536 36363
rect 8484 36320 8536 36329
rect 8668 36320 8720 36372
rect 9864 36320 9916 36372
rect 10600 36320 10652 36372
rect 11888 36320 11940 36372
rect 11980 36320 12032 36372
rect 17960 36320 18012 36372
rect 1584 36227 1636 36236
rect 1584 36193 1593 36227
rect 1593 36193 1627 36227
rect 1627 36193 1636 36227
rect 1584 36184 1636 36193
rect 4620 36116 4672 36168
rect 6736 36159 6788 36168
rect 6736 36125 6745 36159
rect 6745 36125 6779 36159
rect 6779 36125 6788 36159
rect 6736 36116 6788 36125
rect 11520 36184 11572 36236
rect 9588 36159 9640 36168
rect 1768 36091 1820 36100
rect 1768 36057 1777 36091
rect 1777 36057 1811 36091
rect 1811 36057 1820 36091
rect 1768 36048 1820 36057
rect 5448 36048 5500 36100
rect 9588 36125 9597 36159
rect 9597 36125 9631 36159
rect 9631 36125 9640 36159
rect 9588 36116 9640 36125
rect 10600 36116 10652 36168
rect 10692 36116 10744 36168
rect 13176 36184 13228 36236
rect 13820 36184 13872 36236
rect 12992 36116 13044 36168
rect 13084 36159 13136 36168
rect 13084 36125 13093 36159
rect 13093 36125 13127 36159
rect 13127 36125 13136 36159
rect 13084 36116 13136 36125
rect 11888 36048 11940 36100
rect 14464 36091 14516 36100
rect 6736 35980 6788 36032
rect 8024 35980 8076 36032
rect 9036 35980 9088 36032
rect 9404 35980 9456 36032
rect 9680 36023 9732 36032
rect 9680 35989 9689 36023
rect 9689 35989 9723 36023
rect 9723 35989 9732 36023
rect 9680 35980 9732 35989
rect 10416 36023 10468 36032
rect 10416 35989 10425 36023
rect 10425 35989 10459 36023
rect 10459 35989 10468 36023
rect 10416 35980 10468 35989
rect 11060 36023 11112 36032
rect 11060 35989 11069 36023
rect 11069 35989 11103 36023
rect 11103 35989 11112 36023
rect 11060 35980 11112 35989
rect 12072 35980 12124 36032
rect 13544 36023 13596 36032
rect 13544 35989 13553 36023
rect 13553 35989 13587 36023
rect 13587 35989 13596 36023
rect 13544 35980 13596 35989
rect 14464 36057 14473 36091
rect 14473 36057 14507 36091
rect 14507 36057 14516 36091
rect 14464 36048 14516 36057
rect 20628 36252 20680 36304
rect 23480 36320 23532 36372
rect 26608 36363 26660 36372
rect 24584 36252 24636 36304
rect 26608 36329 26617 36363
rect 26617 36329 26651 36363
rect 26651 36329 26660 36363
rect 26608 36320 26660 36329
rect 27068 36320 27120 36372
rect 32404 36320 32456 36372
rect 32496 36320 32548 36372
rect 35900 36320 35952 36372
rect 36176 36320 36228 36372
rect 16856 36184 16908 36236
rect 16948 36184 17000 36236
rect 20536 36184 20588 36236
rect 22284 36184 22336 36236
rect 22560 36184 22612 36236
rect 24768 36184 24820 36236
rect 25136 36227 25188 36236
rect 25136 36193 25145 36227
rect 25145 36193 25179 36227
rect 25179 36193 25188 36227
rect 25136 36184 25188 36193
rect 27988 36184 28040 36236
rect 28448 36184 28500 36236
rect 29092 36184 29144 36236
rect 17868 36116 17920 36168
rect 19432 36116 19484 36168
rect 22100 36116 22152 36168
rect 26240 36116 26292 36168
rect 27068 36159 27120 36168
rect 27068 36125 27077 36159
rect 27077 36125 27111 36159
rect 27111 36125 27120 36159
rect 27068 36116 27120 36125
rect 27712 36159 27764 36168
rect 27712 36125 27721 36159
rect 27721 36125 27755 36159
rect 27755 36125 27764 36159
rect 27712 36116 27764 36125
rect 28172 36116 28224 36168
rect 29000 36116 29052 36168
rect 36268 36252 36320 36304
rect 33692 36184 33744 36236
rect 30472 36116 30524 36168
rect 33508 36116 33560 36168
rect 16212 36091 16264 36100
rect 16212 36057 16221 36091
rect 16221 36057 16255 36091
rect 16255 36057 16264 36091
rect 16212 36048 16264 36057
rect 16672 36048 16724 36100
rect 17776 36048 17828 36100
rect 20996 36091 21048 36100
rect 20996 36057 21005 36091
rect 21005 36057 21039 36091
rect 21039 36057 21048 36091
rect 20996 36048 21048 36057
rect 23112 36048 23164 36100
rect 24584 36048 24636 36100
rect 25228 35980 25280 36032
rect 26424 36048 26476 36100
rect 31116 36048 31168 36100
rect 35256 36048 35308 36100
rect 36176 36116 36228 36168
rect 37832 36116 37884 36168
rect 37740 36048 37792 36100
rect 28356 35980 28408 36032
rect 28448 36023 28500 36032
rect 28448 35989 28457 36023
rect 28457 35989 28491 36023
rect 28491 35989 28500 36023
rect 28448 35980 28500 35989
rect 28632 35980 28684 36032
rect 29184 35980 29236 36032
rect 31300 35980 31352 36032
rect 32588 35980 32640 36032
rect 35532 35980 35584 36032
rect 38200 36023 38252 36032
rect 38200 35989 38209 36023
rect 38209 35989 38243 36023
rect 38243 35989 38252 36023
rect 38200 35980 38252 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1768 35776 1820 35828
rect 8300 35776 8352 35828
rect 10784 35776 10836 35828
rect 12348 35776 12400 35828
rect 13084 35776 13136 35828
rect 14464 35819 14516 35828
rect 14464 35785 14473 35819
rect 14473 35785 14507 35819
rect 14507 35785 14516 35819
rect 14464 35776 14516 35785
rect 3056 35751 3108 35760
rect 3056 35717 3065 35751
rect 3065 35717 3099 35751
rect 3099 35717 3108 35751
rect 3056 35708 3108 35717
rect 3976 35708 4028 35760
rect 9404 35708 9456 35760
rect 1492 35640 1544 35692
rect 2320 35683 2372 35692
rect 2320 35649 2329 35683
rect 2329 35649 2363 35683
rect 2363 35649 2372 35683
rect 2320 35640 2372 35649
rect 6552 35683 6604 35692
rect 6552 35649 6561 35683
rect 6561 35649 6595 35683
rect 6595 35649 6604 35683
rect 6552 35640 6604 35649
rect 8576 35640 8628 35692
rect 11520 35708 11572 35760
rect 11888 35751 11940 35760
rect 11888 35717 11906 35751
rect 11906 35717 11940 35751
rect 11888 35708 11940 35717
rect 12072 35708 12124 35760
rect 29276 35776 29328 35828
rect 31576 35776 31628 35828
rect 17592 35708 17644 35760
rect 18420 35708 18472 35760
rect 19708 35708 19760 35760
rect 20076 35708 20128 35760
rect 23296 35708 23348 35760
rect 33508 35751 33560 35760
rect 33508 35717 33517 35751
rect 33517 35717 33551 35751
rect 33551 35717 33560 35751
rect 33508 35708 33560 35717
rect 35624 35708 35676 35760
rect 10692 35640 10744 35692
rect 11336 35640 11388 35692
rect 8668 35572 8720 35624
rect 9404 35572 9456 35624
rect 10324 35572 10376 35624
rect 12716 35640 12768 35692
rect 16856 35683 16908 35692
rect 12624 35572 12676 35624
rect 12900 35572 12952 35624
rect 13084 35572 13136 35624
rect 16856 35649 16865 35683
rect 16865 35649 16899 35683
rect 16899 35649 16908 35683
rect 16856 35640 16908 35649
rect 22284 35683 22336 35692
rect 22284 35649 22293 35683
rect 22293 35649 22327 35683
rect 22327 35649 22336 35683
rect 22284 35640 22336 35649
rect 31484 35640 31536 35692
rect 34796 35640 34848 35692
rect 38384 35640 38436 35692
rect 17132 35615 17184 35624
rect 17132 35581 17141 35615
rect 17141 35581 17175 35615
rect 17175 35581 17184 35615
rect 17132 35572 17184 35581
rect 17500 35572 17552 35624
rect 19340 35615 19392 35624
rect 2872 35504 2924 35556
rect 8576 35504 8628 35556
rect 10048 35436 10100 35488
rect 10140 35479 10192 35488
rect 10140 35445 10149 35479
rect 10149 35445 10183 35479
rect 10183 35445 10192 35479
rect 16672 35504 16724 35556
rect 10140 35436 10192 35445
rect 16396 35436 16448 35488
rect 17224 35436 17276 35488
rect 19340 35581 19349 35615
rect 19349 35581 19383 35615
rect 19383 35581 19392 35615
rect 19340 35572 19392 35581
rect 19616 35615 19668 35624
rect 19616 35581 19625 35615
rect 19625 35581 19659 35615
rect 19659 35581 19668 35615
rect 19616 35572 19668 35581
rect 19708 35572 19760 35624
rect 23572 35572 23624 35624
rect 27344 35615 27396 35624
rect 27344 35581 27353 35615
rect 27353 35581 27387 35615
rect 27387 35581 27396 35615
rect 27344 35572 27396 35581
rect 23940 35436 23992 35488
rect 27436 35504 27488 35556
rect 33232 35615 33284 35624
rect 33232 35581 33241 35615
rect 33241 35581 33275 35615
rect 33275 35581 33284 35615
rect 33232 35572 33284 35581
rect 35716 35572 35768 35624
rect 28724 35436 28776 35488
rect 34704 35436 34756 35488
rect 37556 35436 37608 35488
rect 38200 35479 38252 35488
rect 38200 35445 38209 35479
rect 38209 35445 38243 35479
rect 38243 35445 38252 35479
rect 38200 35436 38252 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6552 35232 6604 35284
rect 6920 35164 6972 35216
rect 664 35096 716 35148
rect 1400 35028 1452 35080
rect 6460 35071 6512 35080
rect 6460 35037 6469 35071
rect 6469 35037 6503 35071
rect 6503 35037 6512 35071
rect 6460 35028 6512 35037
rect 15384 35232 15436 35284
rect 15568 35232 15620 35284
rect 19616 35232 19668 35284
rect 21824 35232 21876 35284
rect 22192 35232 22244 35284
rect 32312 35232 32364 35284
rect 35256 35232 35308 35284
rect 35716 35232 35768 35284
rect 39304 35232 39356 35284
rect 10508 35164 10560 35216
rect 9312 35096 9364 35148
rect 10048 35096 10100 35148
rect 10876 35096 10928 35148
rect 11336 35164 11388 35216
rect 11520 35164 11572 35216
rect 11888 35164 11940 35216
rect 20076 35164 20128 35216
rect 13176 35096 13228 35148
rect 16856 35096 16908 35148
rect 19340 35096 19392 35148
rect 22284 35096 22336 35148
rect 23480 35096 23532 35148
rect 29092 35096 29144 35148
rect 33232 35096 33284 35148
rect 14004 35028 14056 35080
rect 14372 35028 14424 35080
rect 14648 35028 14700 35080
rect 17316 35028 17368 35080
rect 17500 35028 17552 35080
rect 9312 35003 9364 35012
rect 9312 34969 9321 35003
rect 9321 34969 9355 35003
rect 9355 34969 9364 35003
rect 9312 34960 9364 34969
rect 9680 34960 9732 35012
rect 10784 34960 10836 35012
rect 12164 34960 12216 35012
rect 12256 34960 12308 35012
rect 13176 35003 13228 35012
rect 4988 34892 5040 34944
rect 6552 34935 6604 34944
rect 6552 34901 6561 34935
rect 6561 34901 6595 34935
rect 6595 34901 6604 34935
rect 6552 34892 6604 34901
rect 12808 34892 12860 34944
rect 13176 34969 13185 35003
rect 13185 34969 13219 35003
rect 13219 34969 13228 35003
rect 13176 34960 13228 34969
rect 13268 34960 13320 35012
rect 14556 34892 14608 34944
rect 14648 34892 14700 34944
rect 20352 35028 20404 35080
rect 22928 35071 22980 35080
rect 22928 35037 22937 35071
rect 22937 35037 22971 35071
rect 22971 35037 22980 35071
rect 22928 35028 22980 35037
rect 34428 35028 34480 35080
rect 37556 35071 37608 35080
rect 37556 35037 37565 35071
rect 37565 35037 37599 35071
rect 37599 35037 37608 35071
rect 37556 35028 37608 35037
rect 18788 34960 18840 35012
rect 19984 34960 20036 35012
rect 20720 35003 20772 35012
rect 20720 34969 20729 35003
rect 20729 34969 20763 35003
rect 20763 34969 20772 35003
rect 20720 34960 20772 34969
rect 20812 34960 20864 35012
rect 23112 34960 23164 35012
rect 30288 35003 30340 35012
rect 30288 34969 30297 35003
rect 30297 34969 30331 35003
rect 30331 34969 30340 35003
rect 31208 35003 31260 35012
rect 30288 34960 30340 34969
rect 31208 34969 31217 35003
rect 31217 34969 31251 35003
rect 31251 34969 31260 35003
rect 31208 34960 31260 34969
rect 32588 35003 32640 35012
rect 32588 34969 32597 35003
rect 32597 34969 32631 35003
rect 32631 34969 32640 35003
rect 32588 34960 32640 34969
rect 33324 34960 33376 35012
rect 34612 34960 34664 35012
rect 34704 34960 34756 35012
rect 36820 34960 36872 35012
rect 22100 34892 22152 34944
rect 33416 34892 33468 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2228 34688 2280 34740
rect 5448 34688 5500 34740
rect 10876 34688 10928 34740
rect 10968 34731 11020 34740
rect 10968 34697 10977 34731
rect 10977 34697 11011 34731
rect 11011 34697 11020 34731
rect 10968 34688 11020 34697
rect 3976 34663 4028 34672
rect 3976 34629 3985 34663
rect 3985 34629 4019 34663
rect 4019 34629 4028 34663
rect 3976 34620 4028 34629
rect 6552 34620 6604 34672
rect 10416 34620 10468 34672
rect 11888 34620 11940 34672
rect 12808 34620 12860 34672
rect 13912 34620 13964 34672
rect 14372 34620 14424 34672
rect 2320 34595 2372 34604
rect 2320 34561 2329 34595
rect 2329 34561 2363 34595
rect 2363 34561 2372 34595
rect 2320 34552 2372 34561
rect 3884 34595 3936 34604
rect 3884 34561 3893 34595
rect 3893 34561 3927 34595
rect 3927 34561 3936 34595
rect 3884 34552 3936 34561
rect 4988 34595 5040 34604
rect 4988 34561 4997 34595
rect 4997 34561 5031 34595
rect 5031 34561 5040 34595
rect 4988 34552 5040 34561
rect 8208 34595 8260 34604
rect 8208 34561 8217 34595
rect 8217 34561 8251 34595
rect 8251 34561 8260 34595
rect 8208 34552 8260 34561
rect 8300 34595 8352 34604
rect 8300 34561 8309 34595
rect 8309 34561 8343 34595
rect 8343 34561 8352 34595
rect 8300 34552 8352 34561
rect 10600 34552 10652 34604
rect 10876 34595 10928 34604
rect 10876 34561 10885 34595
rect 10885 34561 10919 34595
rect 10919 34561 10928 34595
rect 10876 34552 10928 34561
rect 11704 34595 11756 34604
rect 11704 34561 11713 34595
rect 11713 34561 11747 34595
rect 11747 34561 11756 34595
rect 11704 34552 11756 34561
rect 14188 34552 14240 34604
rect 15292 34620 15344 34672
rect 10048 34484 10100 34536
rect 10968 34484 11020 34536
rect 13084 34527 13136 34536
rect 13084 34493 13093 34527
rect 13093 34493 13127 34527
rect 13127 34493 13136 34527
rect 13084 34484 13136 34493
rect 14464 34416 14516 34468
rect 19432 34688 19484 34740
rect 19524 34688 19576 34740
rect 20720 34688 20772 34740
rect 18788 34663 18840 34672
rect 18788 34629 18797 34663
rect 18797 34629 18831 34663
rect 18831 34629 18840 34663
rect 18788 34620 18840 34629
rect 22192 34688 22244 34740
rect 20904 34663 20956 34672
rect 20904 34629 20913 34663
rect 20913 34629 20947 34663
rect 20947 34629 20956 34663
rect 31484 34731 31536 34740
rect 31484 34697 31493 34731
rect 31493 34697 31527 34731
rect 31527 34697 31536 34731
rect 31484 34688 31536 34697
rect 20904 34620 20956 34629
rect 24768 34620 24820 34672
rect 30472 34620 30524 34672
rect 19984 34484 20036 34536
rect 22284 34552 22336 34604
rect 27160 34595 27212 34604
rect 27160 34561 27169 34595
rect 27169 34561 27203 34595
rect 27203 34561 27212 34595
rect 27160 34552 27212 34561
rect 28540 34552 28592 34604
rect 30012 34595 30064 34604
rect 30012 34561 30021 34595
rect 30021 34561 30055 34595
rect 30055 34561 30064 34595
rect 30012 34552 30064 34561
rect 31024 34552 31076 34604
rect 33232 34688 33284 34740
rect 33968 34688 34020 34740
rect 38844 34688 38896 34740
rect 35256 34552 35308 34604
rect 35854 34620 35906 34672
rect 37924 34552 37976 34604
rect 29184 34527 29236 34536
rect 1768 34391 1820 34400
rect 1768 34357 1777 34391
rect 1777 34357 1811 34391
rect 1811 34357 1820 34391
rect 1768 34348 1820 34357
rect 11060 34348 11112 34400
rect 18236 34416 18288 34468
rect 29184 34493 29193 34527
rect 29193 34493 29227 34527
rect 29227 34493 29236 34527
rect 29184 34484 29236 34493
rect 29276 34484 29328 34536
rect 36176 34527 36228 34536
rect 36176 34493 36185 34527
rect 36185 34493 36219 34527
rect 36219 34493 36228 34527
rect 36176 34484 36228 34493
rect 16304 34391 16356 34400
rect 16304 34357 16313 34391
rect 16313 34357 16347 34391
rect 16347 34357 16356 34391
rect 16304 34348 16356 34357
rect 16672 34348 16724 34400
rect 24584 34416 24636 34468
rect 23572 34348 23624 34400
rect 24032 34348 24084 34400
rect 29000 34348 29052 34400
rect 32680 34348 32732 34400
rect 38200 34391 38252 34400
rect 38200 34357 38209 34391
rect 38209 34357 38243 34391
rect 38243 34357 38252 34391
rect 38200 34348 38252 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 9588 34144 9640 34196
rect 11428 34076 11480 34128
rect 12256 34076 12308 34128
rect 13176 34144 13228 34196
rect 13360 34144 13412 34196
rect 14280 34144 14332 34196
rect 15200 34144 15252 34196
rect 18236 34144 18288 34196
rect 19984 34144 20036 34196
rect 27344 34144 27396 34196
rect 30288 34144 30340 34196
rect 35716 34144 35768 34196
rect 2136 33983 2188 33992
rect 2136 33949 2145 33983
rect 2145 33949 2179 33983
rect 2179 33949 2188 33983
rect 2136 33940 2188 33949
rect 2780 33983 2832 33992
rect 2780 33949 2789 33983
rect 2789 33949 2823 33983
rect 2823 33949 2832 33983
rect 2780 33940 2832 33949
rect 6920 33940 6972 33992
rect 11704 33940 11756 33992
rect 12164 33940 12216 33992
rect 12256 33940 12308 33992
rect 13084 33940 13136 33992
rect 14556 33983 14608 33992
rect 14556 33949 14565 33983
rect 14565 33949 14599 33983
rect 14599 33949 14608 33983
rect 14556 33940 14608 33949
rect 1584 33804 1636 33856
rect 2872 33847 2924 33856
rect 2872 33813 2881 33847
rect 2881 33813 2915 33847
rect 2915 33813 2924 33847
rect 2872 33804 2924 33813
rect 11152 33804 11204 33856
rect 12072 33847 12124 33856
rect 12072 33813 12081 33847
rect 12081 33813 12115 33847
rect 12115 33813 12124 33847
rect 12072 33804 12124 33813
rect 13636 33804 13688 33856
rect 14464 33872 14516 33924
rect 16856 34008 16908 34060
rect 19340 34008 19392 34060
rect 32680 34076 32732 34128
rect 22100 34008 22152 34060
rect 22836 34008 22888 34060
rect 17684 33940 17736 33992
rect 18604 33940 18656 33992
rect 22008 33940 22060 33992
rect 25412 33983 25464 33992
rect 25412 33949 25421 33983
rect 25421 33949 25455 33983
rect 25455 33949 25464 33983
rect 25412 33940 25464 33949
rect 26148 33940 26200 33992
rect 15936 33872 15988 33924
rect 16120 33872 16172 33924
rect 15568 33804 15620 33856
rect 15752 33804 15804 33856
rect 19616 33872 19668 33924
rect 17132 33847 17184 33856
rect 17132 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17184 33847
rect 17132 33804 17184 33813
rect 17408 33804 17460 33856
rect 21180 33872 21232 33924
rect 22100 33872 22152 33924
rect 22468 33915 22520 33924
rect 22468 33881 22477 33915
rect 22477 33881 22511 33915
rect 22511 33881 22520 33915
rect 22468 33872 22520 33881
rect 24400 33872 24452 33924
rect 27436 33915 27488 33924
rect 27436 33881 27445 33915
rect 27445 33881 27479 33915
rect 27479 33881 27488 33915
rect 27436 33872 27488 33881
rect 27528 33915 27580 33924
rect 27528 33881 27537 33915
rect 27537 33881 27571 33915
rect 27571 33881 27580 33915
rect 28448 33915 28500 33924
rect 27528 33872 27580 33881
rect 28448 33881 28457 33915
rect 28457 33881 28491 33915
rect 28491 33881 28500 33915
rect 28448 33872 28500 33881
rect 30472 34008 30524 34060
rect 34428 34008 34480 34060
rect 31116 33940 31168 33992
rect 34704 33940 34756 33992
rect 32128 33872 32180 33924
rect 34520 33872 34572 33924
rect 35900 33872 35952 33924
rect 19892 33804 19944 33856
rect 24216 33804 24268 33856
rect 31116 33804 31168 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 9036 33600 9088 33652
rect 4620 33532 4672 33584
rect 8024 33575 8076 33584
rect 8024 33541 8033 33575
rect 8033 33541 8067 33575
rect 8067 33541 8076 33575
rect 8024 33532 8076 33541
rect 9220 33532 9272 33584
rect 10416 33575 10468 33584
rect 10416 33541 10425 33575
rect 10425 33541 10459 33575
rect 10459 33541 10468 33575
rect 10416 33532 10468 33541
rect 11980 33600 12032 33652
rect 13084 33600 13136 33652
rect 8668 33507 8720 33516
rect 8668 33473 8677 33507
rect 8677 33473 8711 33507
rect 8711 33473 8720 33507
rect 8668 33464 8720 33473
rect 5080 33396 5132 33448
rect 5356 33439 5408 33448
rect 5356 33405 5365 33439
rect 5365 33405 5399 33439
rect 5399 33405 5408 33439
rect 5356 33396 5408 33405
rect 6736 33396 6788 33448
rect 12164 33464 12216 33516
rect 16120 33532 16172 33584
rect 17132 33600 17184 33652
rect 18604 33643 18656 33652
rect 18604 33609 18613 33643
rect 18613 33609 18647 33643
rect 18647 33609 18656 33643
rect 18604 33600 18656 33609
rect 19064 33600 19116 33652
rect 22100 33600 22152 33652
rect 24952 33643 25004 33652
rect 24952 33609 24961 33643
rect 24961 33609 24995 33643
rect 24995 33609 25004 33643
rect 24952 33600 25004 33609
rect 27436 33600 27488 33652
rect 19984 33532 20036 33584
rect 24492 33532 24544 33584
rect 25044 33532 25096 33584
rect 30012 33532 30064 33584
rect 34428 33532 34480 33584
rect 35532 33532 35584 33584
rect 13728 33464 13780 33516
rect 16672 33464 16724 33516
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 10140 33396 10192 33448
rect 10508 33396 10560 33448
rect 10692 33396 10744 33448
rect 12256 33396 12308 33448
rect 13176 33328 13228 33380
rect 14648 33396 14700 33448
rect 15936 33396 15988 33448
rect 16396 33396 16448 33448
rect 17776 33396 17828 33448
rect 15752 33328 15804 33380
rect 9588 33260 9640 33312
rect 13268 33303 13320 33312
rect 13268 33269 13277 33303
rect 13277 33269 13311 33303
rect 13311 33269 13320 33303
rect 13268 33260 13320 33269
rect 13360 33260 13412 33312
rect 27160 33464 27212 33516
rect 29828 33464 29880 33516
rect 31116 33464 31168 33516
rect 32956 33507 33008 33516
rect 32956 33473 32965 33507
rect 32965 33473 32999 33507
rect 32999 33473 33008 33507
rect 32956 33464 33008 33473
rect 21732 33396 21784 33448
rect 22008 33396 22060 33448
rect 24216 33396 24268 33448
rect 25596 33439 25648 33448
rect 25596 33405 25605 33439
rect 25605 33405 25639 33439
rect 25639 33405 25648 33439
rect 25596 33396 25648 33405
rect 26240 33439 26292 33448
rect 26240 33405 26249 33439
rect 26249 33405 26283 33439
rect 26283 33405 26292 33439
rect 26240 33396 26292 33405
rect 28724 33439 28776 33448
rect 28724 33405 28733 33439
rect 28733 33405 28767 33439
rect 28767 33405 28776 33439
rect 28724 33396 28776 33405
rect 29920 33396 29972 33448
rect 35900 33439 35952 33448
rect 35900 33405 35909 33439
rect 35909 33405 35943 33439
rect 35943 33405 35952 33439
rect 36176 33439 36228 33448
rect 35900 33396 35952 33405
rect 36176 33405 36185 33439
rect 36185 33405 36219 33439
rect 36219 33405 36228 33439
rect 36176 33396 36228 33405
rect 38108 33328 38160 33380
rect 20812 33260 20864 33312
rect 20904 33260 20956 33312
rect 25412 33260 25464 33312
rect 27620 33260 27672 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 3884 33056 3936 33108
rect 8208 33056 8260 33108
rect 9220 33099 9272 33108
rect 9220 33065 9229 33099
rect 9229 33065 9263 33099
rect 9263 33065 9272 33099
rect 9220 33056 9272 33065
rect 10324 33099 10376 33108
rect 10324 33065 10333 33099
rect 10333 33065 10367 33099
rect 10367 33065 10376 33099
rect 10324 33056 10376 33065
rect 11520 33056 11572 33108
rect 34060 33056 34112 33108
rect 34520 33056 34572 33108
rect 5080 32920 5132 32972
rect 13820 32988 13872 33040
rect 14096 32988 14148 33040
rect 14924 32988 14976 33040
rect 20168 32988 20220 33040
rect 22100 32988 22152 33040
rect 25044 33031 25096 33040
rect 25044 32997 25053 33031
rect 25053 32997 25087 33031
rect 25087 32997 25096 33031
rect 25044 32988 25096 32997
rect 1584 32895 1636 32904
rect 1584 32861 1593 32895
rect 1593 32861 1627 32895
rect 1627 32861 1636 32895
rect 1584 32852 1636 32861
rect 8392 32852 8444 32904
rect 10232 32895 10284 32904
rect 1768 32759 1820 32768
rect 1768 32725 1777 32759
rect 1777 32725 1811 32759
rect 1811 32725 1820 32759
rect 1768 32716 1820 32725
rect 7288 32716 7340 32768
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 10876 32895 10928 32904
rect 10876 32861 10885 32895
rect 10885 32861 10919 32895
rect 10919 32861 10928 32895
rect 10876 32852 10928 32861
rect 11520 32895 11572 32904
rect 11520 32861 11529 32895
rect 11529 32861 11563 32895
rect 11563 32861 11572 32895
rect 11520 32852 11572 32861
rect 12348 32852 12400 32904
rect 11336 32716 11388 32768
rect 12348 32716 12400 32768
rect 12532 32784 12584 32836
rect 13360 32784 13412 32836
rect 17500 32920 17552 32972
rect 20260 32920 20312 32972
rect 20812 32963 20864 32972
rect 20812 32929 20821 32963
rect 20821 32929 20855 32963
rect 20855 32929 20864 32963
rect 20812 32920 20864 32929
rect 25596 32920 25648 32972
rect 27620 32920 27672 32972
rect 28448 32963 28500 32972
rect 28448 32929 28457 32963
rect 28457 32929 28491 32963
rect 28491 32929 28500 32963
rect 28448 32920 28500 32929
rect 16948 32852 17000 32904
rect 24584 32852 24636 32904
rect 37464 32895 37516 32904
rect 13084 32716 13136 32768
rect 13176 32716 13228 32768
rect 17408 32784 17460 32836
rect 21548 32784 21600 32836
rect 37464 32861 37473 32895
rect 37473 32861 37507 32895
rect 37507 32861 37516 32895
rect 37464 32852 37516 32861
rect 38752 32852 38804 32904
rect 28356 32784 28408 32836
rect 28448 32784 28500 32836
rect 37280 32784 37332 32836
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 10416 32512 10468 32564
rect 14924 32512 14976 32564
rect 15200 32512 15252 32564
rect 7288 32487 7340 32496
rect 7288 32453 7297 32487
rect 7297 32453 7331 32487
rect 7331 32453 7340 32487
rect 7288 32444 7340 32453
rect 10140 32444 10192 32496
rect 2044 32376 2096 32428
rect 12992 32444 13044 32496
rect 13084 32444 13136 32496
rect 15844 32444 15896 32496
rect 17224 32444 17276 32496
rect 18420 32444 18472 32496
rect 10876 32376 10928 32428
rect 11704 32419 11756 32428
rect 11704 32385 11713 32419
rect 11713 32385 11747 32419
rect 11747 32385 11756 32419
rect 11704 32376 11756 32385
rect 12256 32376 12308 32428
rect 14924 32376 14976 32428
rect 16856 32419 16908 32428
rect 7196 32351 7248 32360
rect 7196 32317 7205 32351
rect 7205 32317 7239 32351
rect 7239 32317 7248 32351
rect 7196 32308 7248 32317
rect 10232 32240 10284 32292
rect 1768 32215 1820 32224
rect 1768 32181 1777 32215
rect 1777 32181 1811 32215
rect 1811 32181 1820 32215
rect 1768 32172 1820 32181
rect 10140 32172 10192 32224
rect 10600 32172 10652 32224
rect 14556 32308 14608 32360
rect 15108 32308 15160 32360
rect 16856 32385 16865 32419
rect 16865 32385 16899 32419
rect 16899 32385 16908 32419
rect 16856 32376 16908 32385
rect 18236 32376 18288 32428
rect 21088 32376 21140 32428
rect 15384 32240 15436 32292
rect 19248 32308 19300 32360
rect 21456 32512 21508 32564
rect 28724 32512 28776 32564
rect 38108 32555 38160 32564
rect 38108 32521 38117 32555
rect 38117 32521 38151 32555
rect 38151 32521 38160 32555
rect 38108 32512 38160 32521
rect 23112 32419 23164 32428
rect 23112 32385 23121 32419
rect 23121 32385 23155 32419
rect 23155 32385 23164 32419
rect 23112 32376 23164 32385
rect 26148 32376 26200 32428
rect 38292 32419 38344 32428
rect 38292 32385 38301 32419
rect 38301 32385 38335 32419
rect 38335 32385 38344 32419
rect 38292 32376 38344 32385
rect 21732 32308 21784 32360
rect 22008 32308 22060 32360
rect 26240 32308 26292 32360
rect 15016 32172 15068 32224
rect 16764 32172 16816 32224
rect 16856 32172 16908 32224
rect 18512 32172 18564 32224
rect 18604 32215 18656 32224
rect 18604 32181 18613 32215
rect 18613 32181 18647 32215
rect 18647 32181 18656 32215
rect 22652 32240 22704 32292
rect 21456 32215 21508 32224
rect 18604 32172 18656 32181
rect 21456 32181 21465 32215
rect 21465 32181 21499 32215
rect 21499 32181 21508 32215
rect 21456 32172 21508 32181
rect 26332 32172 26384 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 12072 31968 12124 32020
rect 11152 31875 11204 31884
rect 11152 31841 11161 31875
rect 11161 31841 11195 31875
rect 11195 31841 11204 31875
rect 11152 31832 11204 31841
rect 12532 31832 12584 31884
rect 21088 31968 21140 32020
rect 27528 31968 27580 32020
rect 35900 31968 35952 32020
rect 12808 31900 12860 31952
rect 15016 31900 15068 31952
rect 16672 31900 16724 31952
rect 24032 31943 24084 31952
rect 13360 31875 13412 31884
rect 13360 31841 13369 31875
rect 13369 31841 13403 31875
rect 13403 31841 13412 31875
rect 13360 31832 13412 31841
rect 15384 31875 15436 31884
rect 15384 31841 15393 31875
rect 15393 31841 15427 31875
rect 15427 31841 15436 31875
rect 15384 31832 15436 31841
rect 17868 31832 17920 31884
rect 18512 31832 18564 31884
rect 19248 31832 19300 31884
rect 24032 31909 24041 31943
rect 24041 31909 24075 31943
rect 24075 31909 24084 31943
rect 24032 31900 24084 31909
rect 33508 31900 33560 31952
rect 34060 31900 34112 31952
rect 20076 31832 20128 31884
rect 21640 31832 21692 31884
rect 22652 31832 22704 31884
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 9772 31807 9824 31816
rect 9772 31773 9781 31807
rect 9781 31773 9815 31807
rect 9815 31773 9824 31807
rect 9772 31764 9824 31773
rect 9864 31807 9916 31816
rect 9864 31773 9873 31807
rect 9873 31773 9907 31807
rect 9907 31773 9916 31807
rect 15108 31807 15160 31816
rect 9864 31764 9916 31773
rect 15108 31773 15117 31807
rect 15117 31773 15151 31807
rect 15151 31773 15160 31807
rect 15108 31764 15160 31773
rect 16764 31764 16816 31816
rect 17408 31764 17460 31816
rect 21088 31764 21140 31816
rect 11244 31739 11296 31748
rect 11244 31705 11253 31739
rect 11253 31705 11287 31739
rect 11287 31705 11296 31739
rect 11244 31696 11296 31705
rect 12808 31739 12860 31748
rect 12808 31705 12817 31739
rect 12817 31705 12851 31739
rect 12851 31705 12860 31739
rect 12808 31696 12860 31705
rect 15844 31696 15896 31748
rect 20168 31696 20220 31748
rect 22008 31764 22060 31816
rect 24952 31764 25004 31816
rect 28080 31832 28132 31884
rect 32312 31875 32364 31884
rect 32312 31841 32321 31875
rect 32321 31841 32355 31875
rect 32355 31841 32364 31875
rect 32312 31832 32364 31841
rect 35532 31832 35584 31884
rect 27712 31764 27764 31816
rect 30380 31764 30432 31816
rect 33600 31764 33652 31816
rect 34060 31807 34112 31816
rect 34060 31773 34069 31807
rect 34069 31773 34103 31807
rect 34103 31773 34112 31807
rect 34060 31764 34112 31773
rect 36084 31807 36136 31816
rect 36084 31773 36093 31807
rect 36093 31773 36127 31807
rect 36127 31773 36136 31807
rect 36084 31764 36136 31773
rect 9404 31628 9456 31680
rect 22468 31628 22520 31680
rect 23848 31628 23900 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4620 31424 4672 31476
rect 7196 31424 7248 31476
rect 12808 31424 12860 31476
rect 5264 31288 5316 31340
rect 6644 31288 6696 31340
rect 11060 31356 11112 31408
rect 11704 31331 11756 31340
rect 6368 31220 6420 31272
rect 10416 31152 10468 31204
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 12440 31220 12492 31272
rect 14096 31263 14148 31272
rect 14096 31229 14105 31263
rect 14105 31229 14139 31263
rect 14139 31229 14148 31263
rect 14096 31220 14148 31229
rect 23940 31424 23992 31476
rect 32588 31424 32640 31476
rect 35808 31424 35860 31476
rect 20536 31356 20588 31408
rect 25412 31356 25464 31408
rect 33416 31356 33468 31408
rect 37372 31356 37424 31408
rect 18512 31288 18564 31340
rect 35808 31288 35860 31340
rect 19248 31220 19300 31272
rect 32220 31220 32272 31272
rect 36636 31220 36688 31272
rect 9680 31084 9732 31136
rect 10784 31084 10836 31136
rect 14556 31152 14608 31204
rect 16120 31152 16172 31204
rect 20168 31084 20220 31136
rect 27436 31084 27488 31136
rect 35532 31084 35584 31136
rect 36452 31084 36504 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 8392 30880 8444 30932
rect 10232 30812 10284 30864
rect 11704 30880 11756 30932
rect 24676 30880 24728 30932
rect 26700 30880 26752 30932
rect 34244 30880 34296 30932
rect 9588 30744 9640 30796
rect 13268 30744 13320 30796
rect 13452 30787 13504 30796
rect 13452 30753 13461 30787
rect 13461 30753 13495 30787
rect 13495 30753 13504 30787
rect 13452 30744 13504 30753
rect 4712 30676 4764 30728
rect 12164 30719 12216 30728
rect 12164 30685 12173 30719
rect 12173 30685 12207 30719
rect 12207 30685 12216 30719
rect 12164 30676 12216 30685
rect 14464 30719 14516 30728
rect 14464 30685 14473 30719
rect 14473 30685 14507 30719
rect 14507 30685 14516 30719
rect 14464 30676 14516 30685
rect 9588 30651 9640 30660
rect 9588 30617 9597 30651
rect 9597 30617 9631 30651
rect 9631 30617 9640 30651
rect 9588 30608 9640 30617
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 10784 30651 10836 30660
rect 10784 30617 10793 30651
rect 10793 30617 10827 30651
rect 10827 30617 10836 30651
rect 10784 30608 10836 30617
rect 10600 30540 10652 30592
rect 12808 30540 12860 30592
rect 12992 30540 13044 30592
rect 14832 30608 14884 30660
rect 15108 30744 15160 30796
rect 15568 30744 15620 30796
rect 16764 30744 16816 30796
rect 18512 30744 18564 30796
rect 21824 30787 21876 30796
rect 21824 30753 21833 30787
rect 21833 30753 21867 30787
rect 21867 30753 21876 30787
rect 21824 30744 21876 30753
rect 23848 30787 23900 30796
rect 23848 30753 23857 30787
rect 23857 30753 23891 30787
rect 23891 30753 23900 30787
rect 23848 30744 23900 30753
rect 26148 30744 26200 30796
rect 32220 30744 32272 30796
rect 35900 30744 35952 30796
rect 36452 30787 36504 30796
rect 36452 30753 36461 30787
rect 36461 30753 36495 30787
rect 36495 30753 36504 30787
rect 36452 30744 36504 30753
rect 37280 30787 37332 30796
rect 37280 30753 37289 30787
rect 37289 30753 37323 30787
rect 37323 30753 37332 30787
rect 37280 30744 37332 30753
rect 16856 30676 16908 30728
rect 32956 30676 33008 30728
rect 15752 30608 15804 30660
rect 19984 30608 20036 30660
rect 17408 30540 17460 30592
rect 17868 30540 17920 30592
rect 21456 30608 21508 30660
rect 20904 30540 20956 30592
rect 21272 30540 21324 30592
rect 21916 30540 21968 30592
rect 25228 30540 25280 30592
rect 25872 30540 25924 30592
rect 26240 30540 26292 30592
rect 28632 30608 28684 30660
rect 32772 30651 32824 30660
rect 32772 30617 32781 30651
rect 32781 30617 32815 30651
rect 32815 30617 32824 30651
rect 32772 30608 32824 30617
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 8392 30336 8444 30388
rect 8668 30336 8720 30388
rect 9588 30336 9640 30388
rect 12808 30336 12860 30388
rect 16580 30336 16632 30388
rect 24676 30336 24728 30388
rect 29644 30336 29696 30388
rect 10232 30268 10284 30320
rect 11520 30268 11572 30320
rect 8208 30200 8260 30252
rect 9128 30243 9180 30252
rect 9128 30209 9137 30243
rect 9137 30209 9171 30243
rect 9171 30209 9180 30243
rect 9128 30200 9180 30209
rect 9772 30243 9824 30252
rect 9772 30209 9781 30243
rect 9781 30209 9815 30243
rect 9815 30209 9824 30243
rect 9772 30200 9824 30209
rect 14372 30200 14424 30252
rect 15108 30268 15160 30320
rect 15292 30268 15344 30320
rect 16120 30268 16172 30320
rect 36268 30268 36320 30320
rect 18512 30200 18564 30252
rect 23112 30200 23164 30252
rect 27620 30200 27672 30252
rect 30012 30200 30064 30252
rect 38292 30243 38344 30252
rect 38292 30209 38301 30243
rect 38301 30209 38335 30243
rect 38335 30209 38344 30243
rect 38292 30200 38344 30209
rect 11796 30175 11848 30184
rect 10416 30064 10468 30116
rect 11796 30141 11805 30175
rect 11805 30141 11839 30175
rect 11839 30141 11848 30175
rect 11796 30132 11848 30141
rect 13912 30132 13964 30184
rect 12256 30064 12308 30116
rect 14280 30064 14332 30116
rect 18604 30132 18656 30184
rect 16028 30064 16080 30116
rect 16764 30064 16816 30116
rect 18328 30064 18380 30116
rect 19064 30132 19116 30184
rect 29736 30132 29788 30184
rect 30380 30132 30432 30184
rect 34796 30132 34848 30184
rect 35256 30175 35308 30184
rect 35256 30141 35265 30175
rect 35265 30141 35299 30175
rect 35299 30141 35308 30175
rect 35256 30132 35308 30141
rect 10876 29996 10928 30048
rect 12164 29996 12216 30048
rect 16120 29996 16172 30048
rect 16304 30039 16356 30048
rect 16304 30005 16313 30039
rect 16313 30005 16347 30039
rect 16347 30005 16356 30039
rect 16304 29996 16356 30005
rect 19156 29996 19208 30048
rect 26884 29996 26936 30048
rect 37556 30064 37608 30116
rect 36636 29996 36688 30048
rect 38476 29996 38528 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 11520 29835 11572 29844
rect 11520 29801 11529 29835
rect 11529 29801 11563 29835
rect 11563 29801 11572 29835
rect 11520 29792 11572 29801
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 2136 29724 2188 29776
rect 9772 29724 9824 29776
rect 19340 29792 19392 29844
rect 9956 29656 10008 29708
rect 11796 29656 11848 29708
rect 12256 29699 12308 29708
rect 12256 29665 12265 29699
rect 12265 29665 12299 29699
rect 12299 29665 12308 29699
rect 12256 29656 12308 29665
rect 1860 29588 1912 29640
rect 10876 29588 10928 29640
rect 11428 29631 11480 29640
rect 11428 29597 11437 29631
rect 11437 29597 11471 29631
rect 11471 29597 11480 29631
rect 11428 29588 11480 29597
rect 15384 29724 15436 29776
rect 16764 29724 16816 29776
rect 29184 29792 29236 29844
rect 26332 29724 26384 29776
rect 31208 29792 31260 29844
rect 15660 29699 15712 29708
rect 15660 29665 15669 29699
rect 15669 29665 15703 29699
rect 15703 29665 15712 29699
rect 15660 29656 15712 29665
rect 16028 29656 16080 29708
rect 16120 29656 16172 29708
rect 23020 29656 23072 29708
rect 26148 29656 26200 29708
rect 29736 29699 29788 29708
rect 29736 29665 29745 29699
rect 29745 29665 29779 29699
rect 29779 29665 29788 29699
rect 29736 29656 29788 29665
rect 30472 29656 30524 29708
rect 15108 29588 15160 29640
rect 17408 29631 17460 29640
rect 17408 29597 17417 29631
rect 17417 29597 17451 29631
rect 17451 29597 17460 29631
rect 17408 29588 17460 29597
rect 20628 29631 20680 29640
rect 20628 29597 20637 29631
rect 20637 29597 20671 29631
rect 20671 29597 20680 29631
rect 20628 29588 20680 29597
rect 27620 29588 27672 29640
rect 7748 29520 7800 29572
rect 9128 29520 9180 29572
rect 12348 29563 12400 29572
rect 1768 29495 1820 29504
rect 1768 29461 1777 29495
rect 1777 29461 1811 29495
rect 1811 29461 1820 29495
rect 1768 29452 1820 29461
rect 9864 29452 9916 29504
rect 12348 29529 12357 29563
rect 12357 29529 12391 29563
rect 12391 29529 12400 29563
rect 12348 29520 12400 29529
rect 13452 29520 13504 29572
rect 15660 29520 15712 29572
rect 13636 29452 13688 29504
rect 16948 29520 17000 29572
rect 21180 29520 21232 29572
rect 23940 29520 23992 29572
rect 16672 29452 16724 29504
rect 26884 29452 26936 29504
rect 29644 29520 29696 29572
rect 31392 29520 31444 29572
rect 32220 29699 32272 29708
rect 32220 29665 32229 29699
rect 32229 29665 32263 29699
rect 32263 29665 32272 29699
rect 32220 29656 32272 29665
rect 34796 29656 34848 29708
rect 32956 29520 33008 29572
rect 35164 29563 35216 29572
rect 35164 29529 35173 29563
rect 35173 29529 35207 29563
rect 35207 29529 35216 29563
rect 35164 29520 35216 29529
rect 36912 29563 36964 29572
rect 35440 29452 35492 29504
rect 36912 29529 36921 29563
rect 36921 29529 36955 29563
rect 36955 29529 36964 29563
rect 36912 29520 36964 29529
rect 38108 29563 38160 29572
rect 38108 29529 38117 29563
rect 38117 29529 38151 29563
rect 38151 29529 38160 29563
rect 38108 29520 38160 29529
rect 37004 29452 37056 29504
rect 38200 29495 38252 29504
rect 38200 29461 38209 29495
rect 38209 29461 38243 29495
rect 38243 29461 38252 29495
rect 38200 29452 38252 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4712 29291 4764 29300
rect 4712 29257 4721 29291
rect 4721 29257 4755 29291
rect 4755 29257 4764 29291
rect 4712 29248 4764 29257
rect 8024 29180 8076 29232
rect 11704 29248 11756 29300
rect 12348 29248 12400 29300
rect 9864 29180 9916 29232
rect 16672 29248 16724 29300
rect 16856 29248 16908 29300
rect 13176 29223 13228 29232
rect 13176 29189 13185 29223
rect 13185 29189 13219 29223
rect 13219 29189 13228 29223
rect 13176 29180 13228 29189
rect 14096 29223 14148 29232
rect 14096 29189 14105 29223
rect 14105 29189 14139 29223
rect 14139 29189 14148 29223
rect 14096 29180 14148 29189
rect 16580 29180 16632 29232
rect 23112 29248 23164 29300
rect 31300 29248 31352 29300
rect 35164 29248 35216 29300
rect 28264 29180 28316 29232
rect 34060 29180 34112 29232
rect 6828 29112 6880 29164
rect 11060 29112 11112 29164
rect 12256 29112 12308 29164
rect 14648 29112 14700 29164
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 22008 29155 22060 29164
rect 22008 29121 22017 29155
rect 22017 29121 22051 29155
rect 22051 29121 22060 29155
rect 22008 29112 22060 29121
rect 26148 29112 26200 29164
rect 32220 29112 32272 29164
rect 38292 29155 38344 29164
rect 38292 29121 38301 29155
rect 38301 29121 38335 29155
rect 38335 29121 38344 29155
rect 38292 29112 38344 29121
rect 1584 29087 1636 29096
rect 1584 29053 1593 29087
rect 1593 29053 1627 29087
rect 1627 29053 1636 29087
rect 1584 29044 1636 29053
rect 1952 29044 2004 29096
rect 12716 29044 12768 29096
rect 16396 29044 16448 29096
rect 16948 29044 17000 29096
rect 17776 29044 17828 29096
rect 18144 29044 18196 29096
rect 13452 28976 13504 29028
rect 14648 29019 14700 29028
rect 14648 28985 14657 29019
rect 14657 28985 14691 29019
rect 14691 28985 14700 29019
rect 14648 28976 14700 28985
rect 16120 28976 16172 29028
rect 11428 28908 11480 28960
rect 16488 28908 16540 28960
rect 17500 28976 17552 29028
rect 20720 29044 20772 29096
rect 33140 29044 33192 29096
rect 36544 29044 36596 29096
rect 39212 29044 39264 29096
rect 29000 29019 29052 29028
rect 29000 28985 29009 29019
rect 29009 28985 29043 29019
rect 29043 28985 29052 29019
rect 29000 28976 29052 28985
rect 29276 28976 29328 29028
rect 38108 29019 38160 29028
rect 38108 28985 38117 29019
rect 38117 28985 38151 29019
rect 38151 28985 38160 29019
rect 38108 28976 38160 28985
rect 16764 28908 16816 28960
rect 17960 28908 18012 28960
rect 19156 28908 19208 28960
rect 20076 28951 20128 28960
rect 20076 28917 20085 28951
rect 20085 28917 20119 28951
rect 20119 28917 20128 28951
rect 20076 28908 20128 28917
rect 27344 28908 27396 28960
rect 35440 28908 35492 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6828 28704 6880 28756
rect 11244 28747 11296 28756
rect 11244 28713 11253 28747
rect 11253 28713 11287 28747
rect 11287 28713 11296 28747
rect 11244 28704 11296 28713
rect 32864 28704 32916 28756
rect 12532 28636 12584 28688
rect 16120 28636 16172 28688
rect 11888 28568 11940 28620
rect 12440 28611 12492 28620
rect 12440 28577 12449 28611
rect 12449 28577 12483 28611
rect 12483 28577 12492 28611
rect 12440 28568 12492 28577
rect 15108 28568 15160 28620
rect 17776 28568 17828 28620
rect 4620 28500 4672 28552
rect 7196 28500 7248 28552
rect 7564 28543 7616 28552
rect 7564 28509 7573 28543
rect 7573 28509 7607 28543
rect 7607 28509 7616 28543
rect 7564 28500 7616 28509
rect 11796 28500 11848 28552
rect 13544 28543 13596 28552
rect 13544 28509 13553 28543
rect 13553 28509 13587 28543
rect 13587 28509 13596 28543
rect 13544 28500 13596 28509
rect 18144 28500 18196 28552
rect 20720 28568 20772 28620
rect 32220 28568 32272 28620
rect 8392 28432 8444 28484
rect 10048 28432 10100 28484
rect 10784 28432 10836 28484
rect 4988 28407 5040 28416
rect 4988 28373 4997 28407
rect 4997 28373 5031 28407
rect 5031 28373 5040 28407
rect 4988 28364 5040 28373
rect 12256 28432 12308 28484
rect 16488 28475 16540 28484
rect 16488 28441 16497 28475
rect 16497 28441 16531 28475
rect 16531 28441 16540 28475
rect 16488 28432 16540 28441
rect 18512 28432 18564 28484
rect 19432 28432 19484 28484
rect 20076 28432 20128 28484
rect 32772 28475 32824 28484
rect 19340 28364 19392 28416
rect 32772 28441 32781 28475
rect 32781 28441 32815 28475
rect 32815 28441 32824 28475
rect 32772 28432 32824 28441
rect 33048 28432 33100 28484
rect 33784 28432 33836 28484
rect 20812 28364 20864 28416
rect 34244 28407 34296 28416
rect 34244 28373 34253 28407
rect 34253 28373 34287 28407
rect 34287 28373 34296 28407
rect 34244 28364 34296 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 7472 28024 7524 28076
rect 11888 28160 11940 28212
rect 9312 28092 9364 28144
rect 12532 28160 12584 28212
rect 4988 27956 5040 28008
rect 16304 28160 16356 28212
rect 16488 28160 16540 28212
rect 23296 28160 23348 28212
rect 14372 28092 14424 28144
rect 15108 28092 15160 28144
rect 17500 28092 17552 28144
rect 20536 28092 20588 28144
rect 21364 28092 21416 28144
rect 26884 28092 26936 28144
rect 27436 28135 27488 28144
rect 27436 28101 27445 28135
rect 27445 28101 27479 28135
rect 27479 28101 27488 28135
rect 27436 28092 27488 28101
rect 28724 28092 28776 28144
rect 29184 28135 29236 28144
rect 29184 28101 29193 28135
rect 29193 28101 29227 28135
rect 29227 28101 29236 28135
rect 29184 28092 29236 28101
rect 29644 28092 29696 28144
rect 32496 28092 32548 28144
rect 34796 28092 34848 28144
rect 14556 28067 14608 28076
rect 14556 28033 14565 28067
rect 14565 28033 14599 28067
rect 14599 28033 14608 28067
rect 14556 28024 14608 28033
rect 20720 28024 20772 28076
rect 13084 27956 13136 28008
rect 13360 27999 13412 28008
rect 13360 27965 13369 27999
rect 13369 27965 13403 27999
rect 13403 27965 13412 27999
rect 13360 27956 13412 27965
rect 14832 27999 14884 28008
rect 14832 27965 14841 27999
rect 14841 27965 14875 27999
rect 14875 27965 14884 27999
rect 14832 27956 14884 27965
rect 15568 27956 15620 28008
rect 17224 27956 17276 28008
rect 17776 27999 17828 28008
rect 17776 27965 17785 27999
rect 17785 27965 17819 27999
rect 17819 27965 17828 27999
rect 17776 27956 17828 27965
rect 7840 27863 7892 27872
rect 7840 27829 7849 27863
rect 7849 27829 7883 27863
rect 7883 27829 7892 27863
rect 7840 27820 7892 27829
rect 7932 27820 7984 27872
rect 10324 27863 10376 27872
rect 10324 27829 10333 27863
rect 10333 27829 10367 27863
rect 10367 27829 10376 27863
rect 10324 27820 10376 27829
rect 11520 27820 11572 27872
rect 11888 27820 11940 27872
rect 18420 27956 18472 28008
rect 20168 27956 20220 28008
rect 26332 27956 26384 28008
rect 26424 27956 26476 28008
rect 33140 27999 33192 28008
rect 33140 27965 33149 27999
rect 33149 27965 33183 27999
rect 33183 27965 33192 27999
rect 33140 27956 33192 27965
rect 19248 27888 19300 27940
rect 20812 27888 20864 27940
rect 30472 27820 30524 27872
rect 30932 27820 30984 27872
rect 33876 27820 33928 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4620 27616 4672 27668
rect 7104 27616 7156 27668
rect 7196 27616 7248 27668
rect 13544 27616 13596 27668
rect 25964 27616 26016 27668
rect 27160 27616 27212 27668
rect 34612 27616 34664 27668
rect 36912 27616 36964 27668
rect 12900 27548 12952 27600
rect 14372 27591 14424 27600
rect 14372 27557 14381 27591
rect 14381 27557 14415 27591
rect 14415 27557 14424 27591
rect 14372 27548 14424 27557
rect 14832 27548 14884 27600
rect 15384 27548 15436 27600
rect 7840 27480 7892 27532
rect 13176 27480 13228 27532
rect 14096 27480 14148 27532
rect 17776 27480 17828 27532
rect 23204 27480 23256 27532
rect 23296 27480 23348 27532
rect 31116 27480 31168 27532
rect 33232 27480 33284 27532
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 7932 27455 7984 27464
rect 7932 27421 7941 27455
rect 7941 27421 7975 27455
rect 7975 27421 7984 27455
rect 7932 27412 7984 27421
rect 12348 27412 12400 27464
rect 12808 27412 12860 27464
rect 15568 27412 15620 27464
rect 26424 27412 26476 27464
rect 32404 27412 32456 27464
rect 37280 27480 37332 27532
rect 34428 27412 34480 27464
rect 38292 27455 38344 27464
rect 38292 27421 38301 27455
rect 38301 27421 38335 27455
rect 38335 27421 38344 27455
rect 38292 27412 38344 27421
rect 1676 27387 1728 27396
rect 1676 27353 1685 27387
rect 1685 27353 1719 27387
rect 1719 27353 1728 27387
rect 1676 27344 1728 27353
rect 5448 27344 5500 27396
rect 10232 27344 10284 27396
rect 11520 27387 11572 27396
rect 11520 27353 11529 27387
rect 11529 27353 11563 27387
rect 11563 27353 11572 27387
rect 13084 27387 13136 27396
rect 11520 27344 11572 27353
rect 13084 27353 13093 27387
rect 13093 27353 13127 27387
rect 13127 27353 13136 27387
rect 13084 27344 13136 27353
rect 7012 27276 7064 27328
rect 12072 27276 12124 27328
rect 17408 27319 17460 27328
rect 17408 27285 17417 27319
rect 17417 27285 17451 27319
rect 17451 27285 17460 27319
rect 17408 27276 17460 27285
rect 22468 27344 22520 27396
rect 26976 27387 27028 27396
rect 26976 27353 26985 27387
rect 26985 27353 27019 27387
rect 27019 27353 27028 27387
rect 26976 27344 27028 27353
rect 29092 27344 29144 27396
rect 30472 27344 30524 27396
rect 31668 27344 31720 27396
rect 39580 27344 39632 27396
rect 21548 27319 21600 27328
rect 21548 27285 21557 27319
rect 21557 27285 21591 27319
rect 21591 27285 21600 27319
rect 21548 27276 21600 27285
rect 31760 27276 31812 27328
rect 32312 27276 32364 27328
rect 35532 27276 35584 27328
rect 39304 27276 39356 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 12072 27115 12124 27124
rect 12072 27081 12081 27115
rect 12081 27081 12115 27115
rect 12115 27081 12124 27115
rect 12072 27072 12124 27081
rect 13084 27072 13136 27124
rect 20536 27072 20588 27124
rect 21548 27072 21600 27124
rect 31668 27072 31720 27124
rect 6828 27004 6880 27056
rect 10324 27004 10376 27056
rect 11520 27004 11572 27056
rect 12716 27004 12768 27056
rect 14188 27004 14240 27056
rect 18880 27004 18932 27056
rect 7012 26979 7064 26988
rect 7012 26945 7021 26979
rect 7021 26945 7055 26979
rect 7055 26945 7064 26979
rect 7012 26936 7064 26945
rect 12808 26936 12860 26988
rect 14556 26979 14608 26988
rect 14556 26945 14565 26979
rect 14565 26945 14599 26979
rect 14599 26945 14608 26979
rect 14556 26936 14608 26945
rect 17960 26936 18012 26988
rect 18144 26979 18196 26988
rect 18144 26945 18153 26979
rect 18153 26945 18187 26979
rect 18187 26945 18196 26979
rect 18144 26936 18196 26945
rect 22008 26936 22060 26988
rect 27620 26979 27672 26988
rect 27620 26945 27629 26979
rect 27629 26945 27663 26979
rect 27663 26945 27672 26979
rect 27620 26936 27672 26945
rect 6000 26868 6052 26920
rect 10048 26868 10100 26920
rect 10692 26868 10744 26920
rect 7196 26843 7248 26852
rect 7196 26809 7205 26843
rect 7205 26809 7239 26843
rect 7239 26809 7248 26843
rect 7196 26800 7248 26809
rect 14096 26868 14148 26920
rect 16304 26868 16356 26920
rect 18052 26868 18104 26920
rect 18420 26911 18472 26920
rect 18420 26877 18429 26911
rect 18429 26877 18463 26911
rect 18463 26877 18472 26911
rect 18420 26868 18472 26877
rect 26424 26868 26476 26920
rect 29368 26868 29420 26920
rect 15844 26800 15896 26852
rect 17316 26800 17368 26852
rect 7104 26732 7156 26784
rect 10876 26732 10928 26784
rect 11796 26732 11848 26784
rect 15936 26732 15988 26784
rect 16396 26732 16448 26784
rect 18788 26732 18840 26784
rect 21456 26800 21508 26852
rect 30380 26868 30432 26920
rect 31024 26868 31076 26920
rect 20536 26732 20588 26784
rect 30840 26800 30892 26852
rect 34612 27072 34664 27124
rect 33048 27004 33100 27056
rect 38568 27004 38620 27056
rect 33140 26868 33192 26920
rect 30196 26732 30248 26784
rect 31300 26775 31352 26784
rect 31300 26741 31309 26775
rect 31309 26741 31343 26775
rect 31343 26741 31352 26775
rect 31300 26732 31352 26741
rect 35624 26868 35676 26920
rect 33600 26732 33652 26784
rect 34428 26732 34480 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 7564 26528 7616 26580
rect 10232 26460 10284 26512
rect 6828 26392 6880 26444
rect 1768 26367 1820 26376
rect 1768 26333 1777 26367
rect 1777 26333 1811 26367
rect 1811 26333 1820 26367
rect 1768 26324 1820 26333
rect 4712 26324 4764 26376
rect 5448 26324 5500 26376
rect 8852 26324 8904 26376
rect 22744 26528 22796 26580
rect 34704 26528 34756 26580
rect 12716 26460 12768 26512
rect 15568 26460 15620 26512
rect 27436 26460 27488 26512
rect 30840 26460 30892 26512
rect 33048 26460 33100 26512
rect 39396 26460 39448 26512
rect 10692 26392 10744 26444
rect 13360 26435 13412 26444
rect 13360 26401 13369 26435
rect 13369 26401 13403 26435
rect 13403 26401 13412 26435
rect 13360 26392 13412 26401
rect 14556 26392 14608 26444
rect 15936 26435 15988 26444
rect 15936 26401 15945 26435
rect 15945 26401 15979 26435
rect 15979 26401 15988 26435
rect 15936 26392 15988 26401
rect 17408 26392 17460 26444
rect 20720 26435 20772 26444
rect 20720 26401 20729 26435
rect 20729 26401 20763 26435
rect 20763 26401 20772 26435
rect 20720 26392 20772 26401
rect 22836 26392 22888 26444
rect 26424 26392 26476 26444
rect 30564 26392 30616 26444
rect 31116 26392 31168 26444
rect 33600 26392 33652 26444
rect 34428 26392 34480 26444
rect 10876 26367 10928 26376
rect 10876 26333 10885 26367
rect 10885 26333 10919 26367
rect 10919 26333 10928 26367
rect 10876 26324 10928 26333
rect 37648 26324 37700 26376
rect 38292 26367 38344 26376
rect 38292 26333 38301 26367
rect 38301 26333 38335 26367
rect 38335 26333 38344 26367
rect 38292 26324 38344 26333
rect 8300 26256 8352 26308
rect 12716 26299 12768 26308
rect 12716 26265 12725 26299
rect 12725 26265 12759 26299
rect 12759 26265 12768 26299
rect 12716 26256 12768 26265
rect 5448 26231 5500 26240
rect 5448 26197 5457 26231
rect 5457 26197 5491 26231
rect 5491 26197 5500 26231
rect 5448 26188 5500 26197
rect 14832 26256 14884 26308
rect 20352 26256 20404 26308
rect 22560 26256 22612 26308
rect 26332 26299 26384 26308
rect 26332 26265 26341 26299
rect 26341 26265 26375 26299
rect 26375 26265 26384 26299
rect 26332 26256 26384 26265
rect 29552 26256 29604 26308
rect 31760 26299 31812 26308
rect 31760 26265 31769 26299
rect 31769 26265 31803 26299
rect 31803 26265 31812 26299
rect 31760 26256 31812 26265
rect 34520 26256 34572 26308
rect 13820 26188 13872 26240
rect 16764 26188 16816 26240
rect 25044 26188 25096 26240
rect 25872 26188 25924 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 5264 25984 5316 26036
rect 10968 25984 11020 26036
rect 11704 25984 11756 26036
rect 13820 26027 13872 26036
rect 13820 25993 13829 26027
rect 13829 25993 13863 26027
rect 13863 25993 13872 26027
rect 13820 25984 13872 25993
rect 15936 25984 15988 26036
rect 20168 25984 20220 26036
rect 19064 25916 19116 25968
rect 24676 25916 24728 25968
rect 5448 25848 5500 25900
rect 7104 25848 7156 25900
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 5540 25823 5592 25832
rect 5540 25789 5549 25823
rect 5549 25789 5583 25823
rect 5583 25789 5592 25823
rect 5540 25780 5592 25789
rect 9220 25780 9272 25832
rect 9680 25780 9732 25832
rect 10876 25712 10928 25764
rect 6000 25687 6052 25696
rect 6000 25653 6009 25687
rect 6009 25653 6043 25687
rect 6043 25653 6052 25687
rect 6000 25644 6052 25653
rect 7564 25687 7616 25696
rect 7564 25653 7573 25687
rect 7573 25653 7607 25687
rect 7607 25653 7616 25687
rect 7564 25644 7616 25653
rect 7840 25644 7892 25696
rect 14280 25848 14332 25900
rect 15292 25780 15344 25832
rect 19432 25780 19484 25832
rect 19524 25712 19576 25764
rect 22928 25823 22980 25832
rect 22928 25789 22937 25823
rect 22937 25789 22971 25823
rect 22971 25789 22980 25823
rect 22928 25780 22980 25789
rect 23204 25823 23256 25832
rect 23204 25789 23213 25823
rect 23213 25789 23247 25823
rect 23247 25789 23256 25823
rect 23204 25780 23256 25789
rect 26608 25984 26660 26036
rect 37740 26027 37792 26036
rect 28080 25916 28132 25968
rect 37740 25993 37749 26027
rect 37749 25993 37783 26027
rect 37783 25993 37792 26027
rect 37740 25984 37792 25993
rect 33876 25916 33928 25968
rect 35716 25916 35768 25968
rect 26424 25848 26476 25900
rect 29368 25891 29420 25900
rect 29368 25857 29377 25891
rect 29377 25857 29411 25891
rect 29411 25857 29420 25891
rect 29368 25848 29420 25857
rect 30748 25848 30800 25900
rect 33600 25848 33652 25900
rect 38660 25848 38712 25900
rect 24860 25780 24912 25832
rect 28540 25712 28592 25764
rect 14372 25644 14424 25696
rect 19248 25644 19300 25696
rect 20996 25644 21048 25696
rect 27436 25644 27488 25696
rect 30840 25644 30892 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7932 25483 7984 25492
rect 7932 25449 7941 25483
rect 7941 25449 7975 25483
rect 7975 25449 7984 25483
rect 7932 25440 7984 25449
rect 9404 25440 9456 25492
rect 21640 25440 21692 25492
rect 22836 25440 22888 25492
rect 30380 25440 30432 25492
rect 35348 25440 35400 25492
rect 20260 25372 20312 25424
rect 2872 25304 2924 25356
rect 8024 25304 8076 25356
rect 9220 25347 9272 25356
rect 9220 25313 9229 25347
rect 9229 25313 9263 25347
rect 9263 25313 9272 25347
rect 9220 25304 9272 25313
rect 10968 25304 11020 25356
rect 5080 25279 5132 25288
rect 5080 25245 5089 25279
rect 5089 25245 5123 25279
rect 5123 25245 5132 25279
rect 5080 25236 5132 25245
rect 8300 25236 8352 25288
rect 14372 25236 14424 25288
rect 25044 25304 25096 25356
rect 26424 25304 26476 25356
rect 30564 25347 30616 25356
rect 30564 25313 30573 25347
rect 30573 25313 30607 25347
rect 30607 25313 30616 25347
rect 30564 25304 30616 25313
rect 34704 25304 34756 25356
rect 9864 25211 9916 25220
rect 5632 25100 5684 25152
rect 9864 25177 9873 25211
rect 9873 25177 9907 25211
rect 9907 25177 9916 25211
rect 9864 25168 9916 25177
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 16856 25236 16908 25288
rect 15752 25100 15804 25152
rect 16948 25168 17000 25220
rect 18144 25168 18196 25220
rect 34612 25236 34664 25288
rect 37096 25279 37148 25288
rect 37096 25245 37105 25279
rect 37105 25245 37139 25279
rect 37139 25245 37148 25279
rect 37096 25236 37148 25245
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 22284 25168 22336 25220
rect 24952 25168 25004 25220
rect 25044 25168 25096 25220
rect 25412 25211 25464 25220
rect 25412 25177 25421 25211
rect 25421 25177 25455 25211
rect 25455 25177 25464 25211
rect 25412 25168 25464 25177
rect 27528 25168 27580 25220
rect 30840 25211 30892 25220
rect 30840 25177 30849 25211
rect 30849 25177 30883 25211
rect 30883 25177 30892 25211
rect 30840 25168 30892 25177
rect 31852 25168 31904 25220
rect 36176 25168 36228 25220
rect 16856 25100 16908 25152
rect 21180 25100 21232 25152
rect 21364 25100 21416 25152
rect 25596 25100 25648 25152
rect 35348 25100 35400 25152
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 5080 24896 5132 24948
rect 16304 24896 16356 24948
rect 18696 24896 18748 24948
rect 23848 24896 23900 24948
rect 38016 24896 38068 24948
rect 3976 24760 4028 24812
rect 4620 24760 4672 24812
rect 5816 24803 5868 24812
rect 5816 24769 5825 24803
rect 5825 24769 5859 24803
rect 5859 24769 5868 24803
rect 5816 24760 5868 24769
rect 6828 24803 6880 24812
rect 6828 24769 6837 24803
rect 6837 24769 6871 24803
rect 6871 24769 6880 24803
rect 6828 24760 6880 24769
rect 7564 24760 7616 24812
rect 7748 24760 7800 24812
rect 7932 24803 7984 24812
rect 7932 24769 7941 24803
rect 7941 24769 7975 24803
rect 7975 24769 7984 24803
rect 7932 24760 7984 24769
rect 9128 24760 9180 24812
rect 8576 24692 8628 24744
rect 10232 24692 10284 24744
rect 11152 24735 11204 24744
rect 11152 24701 11161 24735
rect 11161 24701 11195 24735
rect 11195 24701 11204 24735
rect 11152 24692 11204 24701
rect 18328 24828 18380 24880
rect 22928 24828 22980 24880
rect 36452 24828 36504 24880
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 19524 24760 19576 24812
rect 15568 24692 15620 24744
rect 18420 24735 18472 24744
rect 18420 24701 18429 24735
rect 18429 24701 18463 24735
rect 18463 24701 18472 24735
rect 18420 24692 18472 24701
rect 19432 24692 19484 24744
rect 29828 24760 29880 24812
rect 5540 24624 5592 24676
rect 6000 24624 6052 24676
rect 9864 24624 9916 24676
rect 13176 24624 13228 24676
rect 14556 24624 14608 24676
rect 1768 24599 1820 24608
rect 1768 24565 1777 24599
rect 1777 24565 1811 24599
rect 1811 24565 1820 24599
rect 1768 24556 1820 24565
rect 6736 24556 6788 24608
rect 8024 24599 8076 24608
rect 8024 24565 8033 24599
rect 8033 24565 8067 24599
rect 8067 24565 8076 24599
rect 8024 24556 8076 24565
rect 15844 24556 15896 24608
rect 18052 24556 18104 24608
rect 20076 24624 20128 24676
rect 27620 24692 27672 24744
rect 28540 24735 28592 24744
rect 22284 24624 22336 24676
rect 22928 24624 22980 24676
rect 20168 24556 20220 24608
rect 28540 24701 28549 24735
rect 28549 24701 28583 24735
rect 28583 24701 28592 24735
rect 28540 24692 28592 24701
rect 31944 24692 31996 24744
rect 33048 24692 33100 24744
rect 33968 24692 34020 24744
rect 29644 24624 29696 24676
rect 29000 24556 29052 24608
rect 30012 24599 30064 24608
rect 30012 24565 30021 24599
rect 30021 24565 30055 24599
rect 30055 24565 30064 24599
rect 30012 24556 30064 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8576 24352 8628 24404
rect 15844 24352 15896 24404
rect 16028 24395 16080 24404
rect 16028 24361 16058 24395
rect 16058 24361 16080 24395
rect 16028 24352 16080 24361
rect 8392 24284 8444 24336
rect 18420 24352 18472 24404
rect 26516 24352 26568 24404
rect 30012 24352 30064 24404
rect 34428 24352 34480 24404
rect 35808 24352 35860 24404
rect 18696 24284 18748 24336
rect 26700 24284 26752 24336
rect 29644 24284 29696 24336
rect 5816 24216 5868 24268
rect 9864 24216 9916 24268
rect 10784 24216 10836 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 27620 24216 27672 24268
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 7288 24191 7340 24200
rect 7288 24157 7297 24191
rect 7297 24157 7331 24191
rect 7331 24157 7340 24191
rect 7288 24148 7340 24157
rect 10140 24148 10192 24200
rect 15568 24148 15620 24200
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 15752 24148 15804 24157
rect 20812 24148 20864 24200
rect 33048 24216 33100 24268
rect 34612 24216 34664 24268
rect 35256 24216 35308 24268
rect 4896 24080 4948 24132
rect 6276 24123 6328 24132
rect 6276 24089 6285 24123
rect 6285 24089 6319 24123
rect 6319 24089 6328 24123
rect 6276 24080 6328 24089
rect 9496 24080 9548 24132
rect 11980 24080 12032 24132
rect 12256 24123 12308 24132
rect 12256 24089 12265 24123
rect 12265 24089 12299 24123
rect 12299 24089 12308 24123
rect 12256 24080 12308 24089
rect 8300 24012 8352 24064
rect 10784 24012 10836 24064
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 14372 24080 14424 24132
rect 16304 24080 16356 24132
rect 17684 24080 17736 24132
rect 18328 24080 18380 24132
rect 16672 24012 16724 24064
rect 17500 24012 17552 24064
rect 29000 24123 29052 24132
rect 29000 24089 29009 24123
rect 29009 24089 29043 24123
rect 29043 24089 29052 24123
rect 34520 24148 34572 24200
rect 38292 24191 38344 24200
rect 38292 24157 38301 24191
rect 38301 24157 38335 24191
rect 38335 24157 38344 24191
rect 38292 24148 38344 24157
rect 29000 24080 29052 24089
rect 19340 24012 19392 24064
rect 19524 24012 19576 24064
rect 24308 24012 24360 24064
rect 30564 24080 30616 24132
rect 35900 24080 35952 24132
rect 31484 24055 31536 24064
rect 31484 24021 31493 24055
rect 31493 24021 31527 24055
rect 31527 24021 31536 24055
rect 31484 24012 31536 24021
rect 33232 24012 33284 24064
rect 38200 24012 38252 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 6276 23808 6328 23860
rect 12256 23808 12308 23860
rect 8300 23783 8352 23792
rect 8300 23749 8309 23783
rect 8309 23749 8343 23783
rect 8343 23749 8352 23783
rect 8300 23740 8352 23749
rect 10968 23740 11020 23792
rect 15752 23808 15804 23860
rect 1952 23672 2004 23724
rect 6736 23715 6788 23724
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 9128 23604 9180 23656
rect 3976 23536 4028 23588
rect 14372 23672 14424 23724
rect 16212 23740 16264 23792
rect 18144 23808 18196 23860
rect 18604 23851 18656 23860
rect 18604 23817 18613 23851
rect 18613 23817 18647 23851
rect 18647 23817 18656 23851
rect 18604 23808 18656 23817
rect 18696 23808 18748 23860
rect 20720 23740 20772 23792
rect 18236 23672 18288 23724
rect 16764 23604 16816 23656
rect 14556 23536 14608 23588
rect 17500 23604 17552 23656
rect 18144 23604 18196 23656
rect 20168 23604 20220 23656
rect 20260 23604 20312 23656
rect 24860 23808 24912 23860
rect 26976 23808 27028 23860
rect 32680 23808 32732 23860
rect 33508 23808 33560 23860
rect 33968 23808 34020 23860
rect 23940 23783 23992 23792
rect 23940 23749 23949 23783
rect 23949 23749 23983 23783
rect 23983 23749 23992 23783
rect 23940 23740 23992 23749
rect 25688 23740 25740 23792
rect 30288 23740 30340 23792
rect 34336 23740 34388 23792
rect 37464 23740 37516 23792
rect 22284 23672 22336 23724
rect 34520 23715 34572 23724
rect 34520 23681 34529 23715
rect 34529 23681 34563 23715
rect 34563 23681 34572 23715
rect 34520 23672 34572 23681
rect 25504 23604 25556 23656
rect 28908 23647 28960 23656
rect 9956 23468 10008 23520
rect 14372 23468 14424 23520
rect 16672 23468 16724 23520
rect 20996 23468 21048 23520
rect 28908 23613 28917 23647
rect 28917 23613 28951 23647
rect 28951 23613 28960 23647
rect 28908 23604 28960 23613
rect 31944 23604 31996 23656
rect 33324 23604 33376 23656
rect 36728 23604 36780 23656
rect 29000 23468 29052 23520
rect 30380 23511 30432 23520
rect 30380 23477 30389 23511
rect 30389 23477 30423 23511
rect 30423 23477 30432 23511
rect 30380 23468 30432 23477
rect 30656 23468 30708 23520
rect 32588 23468 32640 23520
rect 32680 23468 32732 23520
rect 36360 23468 36412 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 9772 23264 9824 23316
rect 13360 23264 13412 23316
rect 15384 23264 15436 23316
rect 16764 23307 16816 23316
rect 8392 23196 8444 23248
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 37832 23307 37884 23316
rect 9496 23128 9548 23180
rect 10324 23171 10376 23180
rect 10324 23137 10333 23171
rect 10333 23137 10367 23171
rect 10367 23137 10376 23171
rect 10324 23128 10376 23137
rect 8116 23060 8168 23112
rect 11796 23060 11848 23112
rect 15752 23128 15804 23180
rect 19432 23128 19484 23180
rect 9772 23035 9824 23044
rect 9772 23001 9781 23035
rect 9781 23001 9815 23035
rect 9815 23001 9824 23035
rect 9772 22992 9824 23001
rect 11888 22992 11940 23044
rect 9404 22924 9456 22976
rect 11244 22924 11296 22976
rect 11796 22924 11848 22976
rect 12164 22924 12216 22976
rect 12532 22967 12584 22976
rect 12532 22933 12541 22967
rect 12541 22933 12575 22967
rect 12575 22933 12584 22967
rect 15292 23035 15344 23044
rect 15292 23001 15301 23035
rect 15301 23001 15335 23035
rect 15335 23001 15344 23035
rect 15292 22992 15344 23001
rect 17408 22992 17460 23044
rect 17684 22992 17736 23044
rect 18696 22992 18748 23044
rect 20076 23035 20128 23044
rect 20076 23001 20085 23035
rect 20085 23001 20119 23035
rect 20119 23001 20128 23035
rect 20076 22992 20128 23001
rect 21364 22992 21416 23044
rect 21824 22992 21876 23044
rect 33324 23196 33376 23248
rect 33692 23239 33744 23248
rect 33692 23205 33701 23239
rect 33701 23205 33735 23239
rect 33735 23205 33744 23239
rect 33692 23196 33744 23205
rect 22284 23171 22336 23180
rect 22284 23137 22293 23171
rect 22293 23137 22327 23171
rect 22327 23137 22336 23171
rect 22284 23128 22336 23137
rect 23756 23128 23808 23180
rect 29000 23128 29052 23180
rect 30472 23128 30524 23180
rect 30656 23128 30708 23180
rect 33232 23128 33284 23180
rect 34612 23128 34664 23180
rect 35624 23128 35676 23180
rect 35808 23128 35860 23180
rect 37832 23273 37841 23307
rect 37841 23273 37875 23307
rect 37875 23273 37884 23307
rect 37832 23264 37884 23273
rect 25780 23103 25832 23112
rect 25780 23069 25789 23103
rect 25789 23069 25823 23103
rect 25823 23069 25832 23103
rect 25780 23060 25832 23069
rect 31576 23060 31628 23112
rect 31944 23103 31996 23112
rect 31944 23069 31953 23103
rect 31953 23069 31987 23103
rect 31987 23069 31996 23103
rect 31944 23060 31996 23069
rect 38200 23060 38252 23112
rect 39028 23060 39080 23112
rect 25964 22992 26016 23044
rect 27068 22992 27120 23044
rect 12532 22924 12584 22933
rect 21456 22924 21508 22976
rect 29368 22992 29420 23044
rect 29920 22992 29972 23044
rect 33876 22992 33928 23044
rect 37832 22992 37884 23044
rect 32036 22924 32088 22976
rect 32496 22924 32548 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 7288 22720 7340 22772
rect 8392 22720 8444 22772
rect 8668 22720 8720 22772
rect 15200 22720 15252 22772
rect 9404 22695 9456 22704
rect 9404 22661 9413 22695
rect 9413 22661 9447 22695
rect 9447 22661 9456 22695
rect 9404 22652 9456 22661
rect 11888 22695 11940 22704
rect 11888 22661 11897 22695
rect 11897 22661 11931 22695
rect 11931 22661 11940 22695
rect 11888 22652 11940 22661
rect 12532 22652 12584 22704
rect 20996 22720 21048 22772
rect 21364 22720 21416 22772
rect 22376 22720 22428 22772
rect 26516 22720 26568 22772
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 11060 22584 11112 22636
rect 12808 22584 12860 22636
rect 12992 22584 13044 22636
rect 17868 22652 17920 22704
rect 19432 22652 19484 22704
rect 20260 22652 20312 22704
rect 24492 22652 24544 22704
rect 22008 22627 22060 22636
rect 22008 22593 22017 22627
rect 22017 22593 22051 22627
rect 22051 22593 22060 22627
rect 22008 22584 22060 22593
rect 22284 22584 22336 22636
rect 24308 22584 24360 22636
rect 25780 22584 25832 22636
rect 29000 22720 29052 22772
rect 27436 22695 27488 22704
rect 27436 22661 27445 22695
rect 27445 22661 27479 22695
rect 27479 22661 27488 22695
rect 27436 22652 27488 22661
rect 28448 22652 28500 22704
rect 36084 22720 36136 22772
rect 36544 22720 36596 22772
rect 36728 22763 36780 22772
rect 36728 22729 36737 22763
rect 36737 22729 36771 22763
rect 36771 22729 36780 22763
rect 36728 22720 36780 22729
rect 37556 22652 37608 22704
rect 31944 22584 31996 22636
rect 34612 22584 34664 22636
rect 37648 22584 37700 22636
rect 4620 22516 4672 22568
rect 9128 22516 9180 22568
rect 11152 22516 11204 22568
rect 11796 22559 11848 22568
rect 11796 22525 11805 22559
rect 11805 22525 11839 22559
rect 11839 22525 11848 22559
rect 11796 22516 11848 22525
rect 11704 22448 11756 22500
rect 18052 22516 18104 22568
rect 18328 22516 18380 22568
rect 12348 22448 12400 22500
rect 12808 22448 12860 22500
rect 9680 22380 9732 22432
rect 13636 22380 13688 22432
rect 20076 22448 20128 22500
rect 22376 22448 22428 22500
rect 28908 22559 28960 22568
rect 28908 22525 28917 22559
rect 28917 22525 28951 22559
rect 28951 22525 28960 22559
rect 28908 22516 28960 22525
rect 31484 22516 31536 22568
rect 31668 22516 31720 22568
rect 33140 22516 33192 22568
rect 25504 22448 25556 22500
rect 38200 22491 38252 22500
rect 38200 22457 38209 22491
rect 38209 22457 38243 22491
rect 38243 22457 38252 22491
rect 38200 22448 38252 22457
rect 23388 22380 23440 22432
rect 33140 22380 33192 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 15568 22176 15620 22228
rect 18420 22176 18472 22228
rect 18696 22219 18748 22228
rect 18696 22185 18705 22219
rect 18705 22185 18739 22219
rect 18739 22185 18748 22219
rect 18696 22176 18748 22185
rect 20076 22176 20128 22228
rect 20260 22176 20312 22228
rect 25596 22176 25648 22228
rect 34704 22176 34756 22228
rect 34888 22176 34940 22228
rect 36452 22176 36504 22228
rect 4620 22108 4672 22160
rect 12072 22108 12124 22160
rect 4804 21972 4856 22024
rect 8392 22015 8444 22024
rect 8392 21981 8401 22015
rect 8401 21981 8435 22015
rect 8435 21981 8444 22015
rect 9220 22040 9272 22092
rect 10600 22040 10652 22092
rect 10876 22040 10928 22092
rect 12532 22040 12584 22092
rect 12808 22083 12860 22092
rect 12808 22049 12817 22083
rect 12817 22049 12851 22083
rect 12851 22049 12860 22083
rect 12808 22040 12860 22049
rect 20720 22083 20772 22092
rect 20720 22049 20729 22083
rect 20729 22049 20763 22083
rect 20763 22049 20772 22083
rect 20720 22040 20772 22049
rect 24492 22108 24544 22160
rect 24768 22108 24820 22160
rect 23020 22083 23072 22092
rect 8392 21972 8444 21981
rect 8024 21904 8076 21956
rect 5632 21836 5684 21888
rect 7564 21836 7616 21888
rect 9036 21904 9088 21956
rect 9680 21904 9732 21956
rect 10416 21904 10468 21956
rect 10968 21904 11020 21956
rect 12348 21947 12400 21956
rect 12348 21913 12357 21947
rect 12357 21913 12391 21947
rect 12391 21913 12400 21947
rect 12348 21904 12400 21913
rect 12256 21836 12308 21888
rect 12532 21836 12584 21888
rect 14740 21947 14792 21956
rect 14740 21913 14749 21947
rect 14749 21913 14783 21947
rect 14783 21913 14792 21947
rect 14740 21904 14792 21913
rect 16764 21904 16816 21956
rect 16948 21904 17000 21956
rect 17132 21904 17184 21956
rect 19248 21972 19300 22024
rect 20444 21972 20496 22024
rect 23020 22049 23029 22083
rect 23029 22049 23063 22083
rect 23063 22049 23072 22083
rect 23020 22040 23072 22049
rect 25780 22040 25832 22092
rect 31944 22040 31996 22092
rect 32312 22040 32364 22092
rect 32864 22040 32916 22092
rect 37464 22083 37516 22092
rect 37464 22049 37473 22083
rect 37473 22049 37507 22083
rect 37507 22049 37516 22083
rect 37464 22040 37516 22049
rect 23296 21972 23348 22024
rect 36452 21972 36504 22024
rect 37188 21972 37240 22024
rect 38016 22015 38068 22024
rect 38016 21981 38025 22015
rect 38025 21981 38059 22015
rect 38059 21981 38068 22015
rect 38016 21972 38068 21981
rect 22192 21904 22244 21956
rect 27436 21904 27488 21956
rect 31208 21904 31260 21956
rect 34796 21904 34848 21956
rect 34980 21947 35032 21956
rect 34980 21913 34989 21947
rect 34989 21913 35023 21947
rect 35023 21913 35032 21947
rect 34980 21904 35032 21913
rect 35072 21947 35124 21956
rect 35072 21913 35081 21947
rect 35081 21913 35115 21947
rect 35115 21913 35124 21947
rect 35072 21904 35124 21913
rect 35440 21904 35492 21956
rect 21272 21836 21324 21888
rect 26792 21836 26844 21888
rect 27160 21836 27212 21888
rect 32864 21836 32916 21888
rect 36544 21836 36596 21888
rect 36912 21836 36964 21888
rect 38200 21879 38252 21888
rect 38200 21845 38209 21879
rect 38209 21845 38243 21879
rect 38243 21845 38252 21879
rect 38200 21836 38252 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 1952 21496 2004 21548
rect 12256 21632 12308 21684
rect 16764 21632 16816 21684
rect 23940 21632 23992 21684
rect 24768 21632 24820 21684
rect 30564 21632 30616 21684
rect 35072 21632 35124 21684
rect 35716 21675 35768 21684
rect 35716 21641 35725 21675
rect 35725 21641 35759 21675
rect 35759 21641 35768 21675
rect 35716 21632 35768 21641
rect 8576 21564 8628 21616
rect 12164 21564 12216 21616
rect 13636 21564 13688 21616
rect 16212 21564 16264 21616
rect 7656 21539 7708 21548
rect 7656 21505 7665 21539
rect 7665 21505 7699 21539
rect 7699 21505 7708 21539
rect 7656 21496 7708 21505
rect 10508 21496 10560 21548
rect 11796 21496 11848 21548
rect 12532 21496 12584 21548
rect 9220 21428 9272 21480
rect 9772 21428 9824 21480
rect 10140 21471 10192 21480
rect 10140 21437 10149 21471
rect 10149 21437 10183 21471
rect 10183 21437 10192 21471
rect 10140 21428 10192 21437
rect 12256 21360 12308 21412
rect 16948 21496 17000 21548
rect 17684 21539 17736 21548
rect 17684 21505 17693 21539
rect 17693 21505 17727 21539
rect 17727 21505 17736 21539
rect 17684 21496 17736 21505
rect 22192 21496 22244 21548
rect 28908 21564 28960 21616
rect 33324 21607 33376 21616
rect 33324 21573 33333 21607
rect 33333 21573 33367 21607
rect 33367 21573 33376 21607
rect 33324 21564 33376 21573
rect 34060 21564 34112 21616
rect 37556 21675 37608 21684
rect 37556 21641 37565 21675
rect 37565 21641 37599 21675
rect 37599 21641 37608 21675
rect 37556 21632 37608 21641
rect 36360 21564 36412 21616
rect 15844 21428 15896 21480
rect 19984 21428 20036 21480
rect 22652 21428 22704 21480
rect 22836 21471 22888 21480
rect 22836 21437 22845 21471
rect 22845 21437 22879 21471
rect 22879 21437 22888 21471
rect 22836 21428 22888 21437
rect 31024 21496 31076 21548
rect 31208 21496 31260 21548
rect 34152 21496 34204 21548
rect 36544 21539 36596 21548
rect 28908 21428 28960 21480
rect 32680 21428 32732 21480
rect 13452 21360 13504 21412
rect 1952 21292 2004 21344
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 12532 21292 12584 21344
rect 12992 21292 13044 21344
rect 17132 21292 17184 21344
rect 19156 21360 19208 21412
rect 26240 21360 26292 21412
rect 30472 21360 30524 21412
rect 34980 21428 35032 21480
rect 36544 21505 36553 21539
rect 36553 21505 36587 21539
rect 36587 21505 36596 21539
rect 36544 21496 36596 21505
rect 37096 21496 37148 21548
rect 37188 21496 37240 21548
rect 22376 21292 22428 21344
rect 23204 21292 23256 21344
rect 25136 21292 25188 21344
rect 31944 21292 31996 21344
rect 34520 21292 34572 21344
rect 34888 21292 34940 21344
rect 35532 21292 35584 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 10876 21088 10928 21140
rect 12256 21088 12308 21140
rect 14740 21088 14792 21140
rect 15200 21088 15252 21140
rect 17040 21088 17092 21140
rect 19340 21088 19392 21140
rect 19432 21088 19484 21140
rect 21180 21131 21232 21140
rect 21180 21097 21189 21131
rect 21189 21097 21223 21131
rect 21223 21097 21232 21131
rect 21180 21088 21232 21097
rect 29092 21088 29144 21140
rect 29828 21131 29880 21140
rect 29828 21097 29837 21131
rect 29837 21097 29871 21131
rect 29871 21097 29880 21131
rect 29828 21088 29880 21097
rect 30748 21131 30800 21140
rect 30748 21097 30757 21131
rect 30757 21097 30791 21131
rect 30791 21097 30800 21131
rect 30748 21088 30800 21097
rect 31852 21088 31904 21140
rect 34152 21131 34204 21140
rect 34152 21097 34161 21131
rect 34161 21097 34195 21131
rect 34195 21097 34204 21131
rect 34152 21088 34204 21097
rect 34796 21088 34848 21140
rect 37372 21088 37424 21140
rect 12624 21020 12676 21072
rect 8484 20952 8536 21004
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 7472 20859 7524 20868
rect 7472 20825 7481 20859
rect 7481 20825 7515 20859
rect 7515 20825 7524 20859
rect 7472 20816 7524 20825
rect 7564 20859 7616 20868
rect 7564 20825 7573 20859
rect 7573 20825 7607 20859
rect 7607 20825 7616 20859
rect 7564 20816 7616 20825
rect 9128 20816 9180 20868
rect 10232 20952 10284 21004
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 10600 20952 10652 21004
rect 11796 20952 11848 21004
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 11060 20884 11112 20936
rect 11428 20884 11480 20936
rect 13452 20884 13504 20936
rect 14372 20884 14424 20936
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 12624 20748 12676 20800
rect 12992 20748 13044 20800
rect 14096 20748 14148 20800
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 18052 20927 18104 20936
rect 14648 20884 14700 20893
rect 18052 20893 18061 20927
rect 18061 20893 18095 20927
rect 18095 20893 18104 20927
rect 18052 20884 18104 20893
rect 18696 20927 18748 20936
rect 18696 20893 18705 20927
rect 18705 20893 18739 20927
rect 18739 20893 18748 20927
rect 18696 20884 18748 20893
rect 19248 20884 19300 20936
rect 21088 21020 21140 21072
rect 20444 20952 20496 21004
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 17040 20859 17092 20868
rect 17040 20825 17049 20859
rect 17049 20825 17083 20859
rect 17083 20825 17092 20859
rect 17040 20816 17092 20825
rect 17224 20816 17276 20868
rect 21272 20816 21324 20868
rect 17868 20748 17920 20800
rect 21548 20748 21600 20800
rect 22008 20952 22060 21004
rect 26424 21020 26476 21072
rect 23940 20952 23992 21004
rect 30472 20952 30524 21004
rect 22192 20884 22244 20936
rect 22652 20884 22704 20936
rect 23296 20927 23348 20936
rect 23296 20893 23305 20927
rect 23305 20893 23339 20927
rect 23339 20893 23348 20927
rect 23296 20884 23348 20893
rect 26056 20884 26108 20936
rect 26332 20884 26384 20936
rect 28908 20927 28960 20936
rect 28908 20893 28917 20927
rect 28917 20893 28951 20927
rect 28951 20893 28960 20927
rect 28908 20884 28960 20893
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 33416 21020 33468 21072
rect 33784 21020 33836 21072
rect 33140 20952 33192 21004
rect 34796 20952 34848 21004
rect 35256 20995 35308 21004
rect 35256 20961 35265 20995
rect 35265 20961 35299 20995
rect 35299 20961 35308 20995
rect 35256 20952 35308 20961
rect 35440 20952 35492 21004
rect 29736 20884 29788 20893
rect 31944 20927 31996 20936
rect 24492 20816 24544 20868
rect 25136 20816 25188 20868
rect 25780 20816 25832 20868
rect 25872 20816 25924 20868
rect 27896 20816 27948 20868
rect 31944 20893 31953 20927
rect 31953 20893 31987 20927
rect 31987 20893 31996 20927
rect 31944 20884 31996 20893
rect 34612 20884 34664 20936
rect 32680 20859 32732 20868
rect 29920 20748 29972 20800
rect 30012 20748 30064 20800
rect 32680 20825 32689 20859
rect 32689 20825 32723 20859
rect 32723 20825 32732 20859
rect 32680 20816 32732 20825
rect 34060 20816 34112 20868
rect 36452 20927 36504 20936
rect 36452 20893 36461 20927
rect 36461 20893 36495 20927
rect 36495 20893 36504 20927
rect 36452 20884 36504 20893
rect 36544 20884 36596 20936
rect 34704 20748 34756 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 1860 20544 1912 20596
rect 5356 20544 5408 20596
rect 6644 20476 6696 20528
rect 9956 20476 10008 20528
rect 1860 20408 1912 20460
rect 7840 20408 7892 20460
rect 11796 20476 11848 20528
rect 10692 20408 10744 20460
rect 5632 20340 5684 20392
rect 7288 20383 7340 20392
rect 7288 20349 7297 20383
rect 7297 20349 7331 20383
rect 7331 20349 7340 20383
rect 7288 20340 7340 20349
rect 10048 20340 10100 20392
rect 12164 20544 12216 20596
rect 16396 20544 16448 20596
rect 18236 20544 18288 20596
rect 18880 20587 18932 20596
rect 18880 20553 18889 20587
rect 18889 20553 18923 20587
rect 18923 20553 18932 20587
rect 18880 20544 18932 20553
rect 12808 20476 12860 20528
rect 13176 20476 13228 20528
rect 14556 20476 14608 20528
rect 14740 20476 14792 20528
rect 16764 20476 16816 20528
rect 17592 20476 17644 20528
rect 22836 20544 22888 20596
rect 23388 20544 23440 20596
rect 20996 20476 21048 20528
rect 23572 20476 23624 20528
rect 23940 20519 23992 20528
rect 23940 20485 23949 20519
rect 23949 20485 23983 20519
rect 23983 20485 23992 20519
rect 23940 20476 23992 20485
rect 7748 20272 7800 20324
rect 10876 20315 10928 20324
rect 5080 20204 5132 20256
rect 8024 20204 8076 20256
rect 8760 20204 8812 20256
rect 10876 20281 10885 20315
rect 10885 20281 10919 20315
rect 10919 20281 10928 20315
rect 12808 20340 12860 20392
rect 17684 20408 17736 20460
rect 18052 20408 18104 20460
rect 13452 20340 13504 20392
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 22008 20408 22060 20460
rect 24124 20408 24176 20460
rect 25412 20544 25464 20596
rect 25688 20544 25740 20596
rect 26516 20544 26568 20596
rect 27160 20544 27212 20596
rect 28172 20544 28224 20596
rect 29736 20544 29788 20596
rect 31116 20587 31168 20596
rect 24676 20476 24728 20528
rect 28540 20519 28592 20528
rect 28540 20485 28549 20519
rect 28549 20485 28583 20519
rect 28583 20485 28592 20519
rect 28540 20476 28592 20485
rect 28632 20476 28684 20528
rect 25688 20451 25740 20460
rect 23204 20340 23256 20392
rect 23296 20340 23348 20392
rect 25688 20417 25697 20451
rect 25697 20417 25731 20451
rect 25731 20417 25740 20451
rect 25688 20408 25740 20417
rect 26516 20408 26568 20460
rect 25136 20340 25188 20392
rect 25412 20340 25464 20392
rect 26056 20340 26108 20392
rect 26240 20340 26292 20392
rect 28172 20340 28224 20392
rect 10876 20272 10928 20281
rect 16672 20272 16724 20324
rect 20812 20272 20864 20324
rect 23020 20272 23072 20324
rect 28816 20408 28868 20460
rect 29460 20408 29512 20460
rect 30380 20451 30432 20460
rect 30380 20417 30389 20451
rect 30389 20417 30423 20451
rect 30423 20417 30432 20451
rect 30380 20408 30432 20417
rect 31116 20553 31125 20587
rect 31125 20553 31159 20587
rect 31159 20553 31168 20587
rect 31116 20544 31168 20553
rect 32588 20544 32640 20596
rect 33140 20544 33192 20596
rect 31944 20476 31996 20528
rect 34520 20519 34572 20528
rect 34520 20485 34529 20519
rect 34529 20485 34563 20519
rect 34563 20485 34572 20519
rect 34520 20476 34572 20485
rect 35900 20544 35952 20596
rect 36084 20544 36136 20596
rect 37280 20544 37332 20596
rect 37740 20544 37792 20596
rect 28908 20340 28960 20392
rect 33048 20408 33100 20460
rect 36268 20451 36320 20460
rect 35348 20340 35400 20392
rect 31300 20272 31352 20324
rect 18788 20204 18840 20256
rect 23388 20204 23440 20256
rect 26424 20204 26476 20256
rect 26516 20204 26568 20256
rect 29736 20204 29788 20256
rect 31208 20204 31260 20256
rect 34796 20204 34848 20256
rect 35440 20272 35492 20324
rect 36268 20417 36277 20451
rect 36277 20417 36311 20451
rect 36311 20417 36320 20451
rect 36268 20408 36320 20417
rect 37188 20408 37240 20460
rect 36084 20204 36136 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6644 20043 6696 20052
rect 6644 20009 6653 20043
rect 6653 20009 6687 20043
rect 6687 20009 6696 20043
rect 6644 20000 6696 20009
rect 10876 20000 10928 20052
rect 11152 20000 11204 20052
rect 14832 20000 14884 20052
rect 16764 20043 16816 20052
rect 16764 20009 16773 20043
rect 16773 20009 16807 20043
rect 16807 20009 16816 20043
rect 16764 20000 16816 20009
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 22560 20000 22612 20052
rect 23204 20000 23256 20052
rect 25136 20000 25188 20052
rect 27528 20000 27580 20052
rect 28908 20043 28960 20052
rect 28908 20009 28917 20043
rect 28917 20009 28951 20043
rect 28951 20009 28960 20043
rect 28908 20000 28960 20009
rect 31392 20043 31444 20052
rect 31392 20009 31401 20043
rect 31401 20009 31435 20043
rect 31435 20009 31444 20043
rect 31392 20000 31444 20009
rect 32680 20000 32732 20052
rect 33324 20000 33376 20052
rect 34060 20000 34112 20052
rect 35440 20000 35492 20052
rect 35716 20000 35768 20052
rect 36176 20043 36228 20052
rect 36176 20009 36185 20043
rect 36185 20009 36219 20043
rect 36219 20009 36228 20043
rect 36176 20000 36228 20009
rect 36728 20000 36780 20052
rect 37924 20000 37976 20052
rect 5448 19932 5500 19984
rect 10324 19932 10376 19984
rect 1860 19864 1912 19916
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 8024 19864 8076 19916
rect 12072 19864 12124 19916
rect 12532 19864 12584 19916
rect 13084 19864 13136 19916
rect 13176 19864 13228 19916
rect 14372 19932 14424 19984
rect 20444 19932 20496 19984
rect 21364 19975 21416 19984
rect 21364 19941 21373 19975
rect 21373 19941 21407 19975
rect 21407 19941 21416 19975
rect 21364 19932 21416 19941
rect 27436 19932 27488 19984
rect 28356 19932 28408 19984
rect 29736 19932 29788 19984
rect 31944 19932 31996 19984
rect 34428 19932 34480 19984
rect 36452 19932 36504 19984
rect 39212 19932 39264 19984
rect 16304 19864 16356 19916
rect 9404 19796 9456 19848
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 12624 19796 12676 19848
rect 14096 19796 14148 19848
rect 1492 19728 1544 19780
rect 11888 19771 11940 19780
rect 9864 19660 9916 19712
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 11888 19737 11897 19771
rect 11897 19737 11931 19771
rect 11931 19737 11940 19771
rect 11888 19728 11940 19737
rect 12992 19771 13044 19780
rect 12992 19737 13001 19771
rect 13001 19737 13035 19771
rect 13035 19737 13044 19771
rect 12992 19728 13044 19737
rect 13084 19771 13136 19780
rect 13084 19737 13093 19771
rect 13093 19737 13127 19771
rect 13127 19737 13136 19771
rect 15936 19796 15988 19848
rect 16580 19796 16632 19848
rect 19156 19864 19208 19916
rect 20996 19864 21048 19916
rect 23020 19864 23072 19916
rect 25320 19864 25372 19916
rect 29460 19864 29512 19916
rect 29828 19907 29880 19916
rect 29828 19873 29837 19907
rect 29837 19873 29871 19907
rect 29871 19873 29880 19907
rect 29828 19864 29880 19873
rect 30472 19907 30524 19916
rect 30472 19873 30481 19907
rect 30481 19873 30515 19907
rect 30515 19873 30524 19907
rect 30472 19864 30524 19873
rect 31024 19864 31076 19916
rect 17684 19796 17736 19848
rect 13084 19728 13136 19737
rect 16764 19728 16816 19780
rect 16948 19728 17000 19780
rect 20812 19728 20864 19780
rect 12072 19660 12124 19712
rect 13912 19660 13964 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 15384 19660 15436 19712
rect 20260 19660 20312 19712
rect 25872 19796 25924 19848
rect 26240 19796 26292 19848
rect 28816 19839 28868 19848
rect 23388 19771 23440 19780
rect 23388 19737 23397 19771
rect 23397 19737 23431 19771
rect 23431 19737 23440 19771
rect 23388 19728 23440 19737
rect 23480 19771 23532 19780
rect 23480 19737 23489 19771
rect 23489 19737 23523 19771
rect 23523 19737 23532 19771
rect 23480 19728 23532 19737
rect 25412 19728 25464 19780
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 30748 19796 30800 19848
rect 31300 19839 31352 19848
rect 31300 19805 31309 19839
rect 31309 19805 31343 19839
rect 31343 19805 31352 19839
rect 31300 19796 31352 19805
rect 31484 19796 31536 19848
rect 36268 19864 36320 19916
rect 33416 19796 33468 19848
rect 36084 19839 36136 19848
rect 36084 19805 36093 19839
rect 36093 19805 36127 19839
rect 36127 19805 36136 19839
rect 36084 19796 36136 19805
rect 36544 19796 36596 19848
rect 37188 19796 37240 19848
rect 37464 19796 37516 19848
rect 29000 19728 29052 19780
rect 29920 19771 29972 19780
rect 29920 19737 29929 19771
rect 29929 19737 29963 19771
rect 29963 19737 29972 19771
rect 29920 19728 29972 19737
rect 32680 19771 32732 19780
rect 32680 19737 32689 19771
rect 32689 19737 32723 19771
rect 32723 19737 32732 19771
rect 32680 19728 32732 19737
rect 35072 19771 35124 19780
rect 35072 19737 35081 19771
rect 35081 19737 35115 19771
rect 35115 19737 35124 19771
rect 35072 19728 35124 19737
rect 35440 19728 35492 19780
rect 24860 19660 24912 19712
rect 28632 19660 28684 19712
rect 33232 19660 33284 19712
rect 33876 19660 33928 19712
rect 34244 19660 34296 19712
rect 34888 19660 34940 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 6828 19456 6880 19508
rect 7656 19456 7708 19508
rect 8760 19431 8812 19440
rect 8760 19397 8769 19431
rect 8769 19397 8803 19431
rect 8803 19397 8812 19431
rect 8760 19388 8812 19397
rect 10968 19388 11020 19440
rect 1768 19363 1820 19372
rect 1768 19329 1777 19363
rect 1777 19329 1811 19363
rect 1811 19329 1820 19363
rect 1768 19320 1820 19329
rect 7748 19320 7800 19372
rect 8116 19320 8168 19372
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 13084 19456 13136 19508
rect 13452 19456 13504 19508
rect 14188 19499 14240 19508
rect 14188 19465 14197 19499
rect 14197 19465 14231 19499
rect 14231 19465 14240 19499
rect 14188 19456 14240 19465
rect 17500 19456 17552 19508
rect 17776 19456 17828 19508
rect 19064 19456 19116 19508
rect 20260 19499 20312 19508
rect 20260 19465 20269 19499
rect 20269 19465 20303 19499
rect 20303 19465 20312 19499
rect 20260 19456 20312 19465
rect 20904 19499 20956 19508
rect 20904 19465 20913 19499
rect 20913 19465 20947 19499
rect 20947 19465 20956 19499
rect 20904 19456 20956 19465
rect 24584 19499 24636 19508
rect 24584 19465 24593 19499
rect 24593 19465 24627 19499
rect 24627 19465 24636 19499
rect 24584 19456 24636 19465
rect 24952 19456 25004 19508
rect 25964 19456 26016 19508
rect 11152 19388 11204 19440
rect 13176 19388 13228 19440
rect 13544 19388 13596 19440
rect 15384 19431 15436 19440
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 12808 19295 12860 19304
rect 12808 19261 12817 19295
rect 12817 19261 12851 19295
rect 12851 19261 12860 19295
rect 12808 19252 12860 19261
rect 15384 19397 15393 19431
rect 15393 19397 15427 19431
rect 15427 19397 15436 19431
rect 15384 19388 15436 19397
rect 16304 19431 16356 19440
rect 16304 19397 16313 19431
rect 16313 19397 16347 19431
rect 16347 19397 16356 19431
rect 16304 19388 16356 19397
rect 20720 19388 20772 19440
rect 16764 19320 16816 19372
rect 17592 19363 17644 19372
rect 17592 19329 17601 19363
rect 17601 19329 17635 19363
rect 17635 19329 17644 19363
rect 17592 19320 17644 19329
rect 17684 19320 17736 19372
rect 19432 19320 19484 19372
rect 20536 19320 20588 19372
rect 20812 19363 20864 19372
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 25320 19388 25372 19440
rect 29000 19456 29052 19508
rect 30196 19456 30248 19508
rect 30288 19456 30340 19508
rect 33232 19499 33284 19508
rect 33232 19465 33241 19499
rect 33241 19465 33275 19499
rect 33275 19465 33284 19499
rect 33232 19456 33284 19465
rect 34336 19456 34388 19508
rect 34796 19456 34848 19508
rect 35256 19456 35308 19508
rect 35992 19456 36044 19508
rect 36820 19499 36872 19508
rect 36820 19465 36829 19499
rect 36829 19465 36863 19499
rect 36863 19465 36872 19499
rect 36820 19456 36872 19465
rect 20812 19320 20864 19329
rect 21640 19320 21692 19372
rect 22652 19320 22704 19372
rect 24124 19320 24176 19372
rect 12440 19184 12492 19236
rect 12624 19116 12676 19168
rect 14004 19184 14056 19236
rect 23020 19252 23072 19304
rect 23940 19252 23992 19304
rect 24768 19320 24820 19372
rect 25412 19363 25464 19372
rect 24860 19252 24912 19304
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 26976 19388 27028 19440
rect 26240 19320 26292 19372
rect 26700 19320 26752 19372
rect 27252 19363 27304 19372
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 27436 19320 27488 19372
rect 29276 19388 29328 19440
rect 31576 19388 31628 19440
rect 34244 19388 34296 19440
rect 35532 19388 35584 19440
rect 31116 19320 31168 19372
rect 31944 19320 31996 19372
rect 22836 19184 22888 19236
rect 25964 19184 26016 19236
rect 22100 19159 22152 19168
rect 22100 19125 22109 19159
rect 22109 19125 22143 19159
rect 22143 19125 22152 19159
rect 22100 19116 22152 19125
rect 24584 19116 24636 19168
rect 28908 19252 28960 19304
rect 29000 19295 29052 19304
rect 29000 19261 29009 19295
rect 29009 19261 29043 19295
rect 29043 19261 29052 19295
rect 29000 19252 29052 19261
rect 30564 19252 30616 19304
rect 34152 19320 34204 19372
rect 34428 19320 34480 19372
rect 35992 19320 36044 19372
rect 36176 19320 36228 19372
rect 37188 19320 37240 19372
rect 36360 19252 36412 19304
rect 28172 19184 28224 19236
rect 33232 19184 33284 19236
rect 26332 19116 26384 19168
rect 29000 19116 29052 19168
rect 31300 19116 31352 19168
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 15568 18955 15620 18964
rect 15568 18921 15577 18955
rect 15577 18921 15611 18955
rect 15611 18921 15620 18955
rect 15568 18912 15620 18921
rect 18512 18912 18564 18964
rect 12900 18844 12952 18896
rect 13728 18844 13780 18896
rect 16948 18844 17000 18896
rect 17868 18844 17920 18896
rect 20904 18844 20956 18896
rect 23388 18844 23440 18896
rect 23572 18912 23624 18964
rect 24216 18912 24268 18964
rect 24768 18912 24820 18964
rect 26332 18955 26384 18964
rect 26332 18921 26341 18955
rect 26341 18921 26375 18955
rect 26375 18921 26384 18955
rect 26332 18912 26384 18921
rect 27804 18912 27856 18964
rect 28816 18912 28868 18964
rect 29552 18912 29604 18964
rect 32312 18912 32364 18964
rect 9588 18819 9640 18828
rect 9588 18785 9597 18819
rect 9597 18785 9631 18819
rect 9631 18785 9640 18819
rect 9588 18776 9640 18785
rect 10048 18776 10100 18828
rect 11980 18776 12032 18828
rect 7748 18708 7800 18760
rect 10600 18640 10652 18692
rect 12256 18683 12308 18692
rect 12256 18649 12265 18683
rect 12265 18649 12299 18683
rect 12299 18649 12308 18683
rect 13176 18683 13228 18692
rect 12256 18640 12308 18649
rect 13176 18649 13185 18683
rect 13185 18649 13219 18683
rect 13219 18649 13228 18683
rect 13176 18640 13228 18649
rect 9312 18572 9364 18624
rect 15200 18708 15252 18760
rect 19984 18776 20036 18828
rect 21272 18819 21324 18828
rect 21272 18785 21281 18819
rect 21281 18785 21315 18819
rect 21315 18785 21324 18819
rect 21272 18776 21324 18785
rect 21548 18776 21600 18828
rect 22468 18776 22520 18828
rect 16948 18708 17000 18760
rect 17684 18708 17736 18760
rect 24584 18751 24636 18760
rect 22100 18640 22152 18692
rect 22836 18683 22888 18692
rect 22836 18649 22845 18683
rect 22845 18649 22879 18683
rect 22879 18649 22888 18683
rect 22836 18640 22888 18649
rect 17040 18572 17092 18624
rect 23664 18572 23716 18624
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 24768 18708 24820 18760
rect 26424 18776 26476 18828
rect 27436 18776 27488 18828
rect 27988 18819 28040 18828
rect 27988 18785 27997 18819
rect 27997 18785 28031 18819
rect 28031 18785 28040 18819
rect 27988 18776 28040 18785
rect 27896 18708 27948 18760
rect 30564 18776 30616 18828
rect 33508 18912 33560 18964
rect 34060 18912 34112 18964
rect 34704 18912 34756 18964
rect 35256 18912 35308 18964
rect 38844 18912 38896 18964
rect 34612 18844 34664 18896
rect 37556 18844 37608 18896
rect 32864 18776 32916 18828
rect 29736 18751 29788 18760
rect 29736 18717 29745 18751
rect 29745 18717 29779 18751
rect 29779 18717 29788 18751
rect 29736 18708 29788 18717
rect 30748 18708 30800 18760
rect 31116 18708 31168 18760
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 34152 18708 34204 18760
rect 37740 18776 37792 18828
rect 23848 18640 23900 18692
rect 25964 18640 26016 18692
rect 26976 18683 27028 18692
rect 26240 18572 26292 18624
rect 26976 18649 26985 18683
rect 26985 18649 27019 18683
rect 27019 18649 27028 18683
rect 26976 18640 27028 18649
rect 27436 18640 27488 18692
rect 32864 18640 32916 18692
rect 33048 18640 33100 18692
rect 35900 18708 35952 18760
rect 36176 18708 36228 18760
rect 37280 18683 37332 18692
rect 37280 18649 37289 18683
rect 37289 18649 37323 18683
rect 37323 18649 37332 18683
rect 37280 18640 37332 18649
rect 37372 18683 37424 18692
rect 37372 18649 37381 18683
rect 37381 18649 37415 18683
rect 37415 18649 37424 18683
rect 37372 18640 37424 18649
rect 30012 18572 30064 18624
rect 32404 18572 32456 18624
rect 37924 18572 37976 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 7472 18368 7524 18420
rect 9772 18368 9824 18420
rect 11520 18368 11572 18420
rect 4620 18232 4672 18284
rect 10508 18300 10560 18352
rect 19248 18368 19300 18420
rect 23480 18368 23532 18420
rect 24400 18411 24452 18420
rect 24400 18377 24409 18411
rect 24409 18377 24443 18411
rect 24443 18377 24452 18411
rect 24400 18368 24452 18377
rect 26056 18411 26108 18420
rect 26056 18377 26065 18411
rect 26065 18377 26099 18411
rect 26099 18377 26108 18411
rect 26056 18368 26108 18377
rect 27436 18411 27488 18420
rect 27436 18377 27445 18411
rect 27445 18377 27479 18411
rect 27479 18377 27488 18411
rect 27436 18368 27488 18377
rect 28724 18411 28776 18420
rect 28724 18377 28733 18411
rect 28733 18377 28767 18411
rect 28767 18377 28776 18411
rect 28724 18368 28776 18377
rect 28908 18368 28960 18420
rect 32128 18368 32180 18420
rect 33600 18411 33652 18420
rect 13912 18343 13964 18352
rect 13912 18309 13921 18343
rect 13921 18309 13955 18343
rect 13955 18309 13964 18343
rect 13912 18300 13964 18309
rect 21916 18300 21968 18352
rect 24768 18300 24820 18352
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 7932 18164 7984 18216
rect 9404 18232 9456 18284
rect 10784 18275 10836 18284
rect 10784 18241 10793 18275
rect 10793 18241 10827 18275
rect 10827 18241 10836 18275
rect 10784 18232 10836 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 19432 18275 19484 18284
rect 19432 18241 19441 18275
rect 19441 18241 19475 18275
rect 19475 18241 19484 18275
rect 19432 18232 19484 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 12624 18164 12676 18216
rect 13268 18207 13320 18216
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 21640 18164 21692 18216
rect 23940 18232 23992 18284
rect 25964 18275 26016 18284
rect 23388 18164 23440 18216
rect 25964 18241 25973 18275
rect 25973 18241 26007 18275
rect 26007 18241 26016 18275
rect 25964 18232 26016 18241
rect 27068 18300 27120 18352
rect 28172 18232 28224 18284
rect 30748 18300 30800 18352
rect 31208 18343 31260 18352
rect 31208 18309 31217 18343
rect 31217 18309 31251 18343
rect 31251 18309 31260 18343
rect 31208 18300 31260 18309
rect 31300 18300 31352 18352
rect 33600 18377 33609 18411
rect 33609 18377 33643 18411
rect 33643 18377 33652 18411
rect 33600 18368 33652 18377
rect 34612 18368 34664 18420
rect 35440 18368 35492 18420
rect 37004 18368 37056 18420
rect 37832 18368 37884 18420
rect 28816 18232 28868 18284
rect 30472 18232 30524 18284
rect 33140 18232 33192 18284
rect 34152 18232 34204 18284
rect 34612 18232 34664 18284
rect 36544 18300 36596 18352
rect 10416 18028 10468 18080
rect 14004 18071 14056 18080
rect 14004 18037 14013 18071
rect 14013 18037 14047 18071
rect 14047 18037 14056 18071
rect 14004 18028 14056 18037
rect 14096 18028 14148 18080
rect 19616 18028 19668 18080
rect 21456 18028 21508 18080
rect 25320 18028 25372 18080
rect 31392 18207 31444 18216
rect 31392 18173 31401 18207
rect 31401 18173 31435 18207
rect 31435 18173 31444 18207
rect 31392 18164 31444 18173
rect 28448 18028 28500 18080
rect 32864 18164 32916 18216
rect 36360 18232 36412 18284
rect 37188 18232 37240 18284
rect 37832 18275 37884 18284
rect 37832 18241 37841 18275
rect 37841 18241 37875 18275
rect 37875 18241 37884 18275
rect 37832 18232 37884 18241
rect 31668 18096 31720 18148
rect 33048 18096 33100 18148
rect 36452 18164 36504 18216
rect 38476 18164 38528 18216
rect 38016 18096 38068 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 11520 17824 11572 17876
rect 12348 17824 12400 17876
rect 20076 17824 20128 17876
rect 24584 17824 24636 17876
rect 25228 17824 25280 17876
rect 28080 17824 28132 17876
rect 28632 17867 28684 17876
rect 28632 17833 28641 17867
rect 28641 17833 28675 17867
rect 28675 17833 28684 17867
rect 28632 17824 28684 17833
rect 30472 17824 30524 17876
rect 34152 17824 34204 17876
rect 38568 17824 38620 17876
rect 21364 17756 21416 17808
rect 30564 17756 30616 17808
rect 31024 17756 31076 17808
rect 7288 17688 7340 17740
rect 7932 17688 7984 17740
rect 9864 17688 9916 17740
rect 13084 17731 13136 17740
rect 13084 17697 13093 17731
rect 13093 17697 13127 17731
rect 13127 17697 13136 17731
rect 13084 17688 13136 17697
rect 20628 17688 20680 17740
rect 30380 17731 30432 17740
rect 14280 17663 14332 17672
rect 8852 17484 8904 17536
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 15660 17620 15712 17672
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 22560 17620 22612 17672
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 23940 17620 23992 17672
rect 25136 17620 25188 17672
rect 25688 17663 25740 17672
rect 25688 17629 25697 17663
rect 25697 17629 25731 17663
rect 25731 17629 25740 17663
rect 25688 17620 25740 17629
rect 9220 17595 9272 17604
rect 9220 17561 9229 17595
rect 9229 17561 9263 17595
rect 9263 17561 9272 17595
rect 9220 17552 9272 17561
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 11152 17595 11204 17604
rect 11152 17561 11161 17595
rect 11161 17561 11195 17595
rect 11195 17561 11204 17595
rect 12072 17595 12124 17604
rect 11152 17552 11204 17561
rect 12072 17561 12081 17595
rect 12081 17561 12115 17595
rect 12115 17561 12124 17595
rect 12072 17552 12124 17561
rect 10784 17484 10836 17536
rect 15108 17552 15160 17604
rect 16672 17552 16724 17604
rect 27252 17552 27304 17604
rect 30380 17697 30389 17731
rect 30389 17697 30423 17731
rect 30423 17697 30432 17731
rect 30380 17688 30432 17697
rect 31392 17688 31444 17740
rect 31668 17688 31720 17740
rect 27896 17663 27948 17672
rect 27896 17629 27905 17663
rect 27905 17629 27939 17663
rect 27939 17629 27948 17663
rect 27896 17620 27948 17629
rect 28172 17620 28224 17672
rect 35348 17688 35400 17740
rect 35900 17731 35952 17740
rect 35900 17697 35909 17731
rect 35909 17697 35943 17731
rect 35943 17697 35952 17731
rect 35900 17688 35952 17697
rect 39580 17756 39632 17808
rect 37740 17688 37792 17740
rect 29000 17552 29052 17604
rect 29828 17595 29880 17604
rect 29828 17561 29837 17595
rect 29837 17561 29871 17595
rect 29871 17561 29880 17595
rect 29828 17552 29880 17561
rect 33508 17663 33560 17672
rect 33508 17629 33517 17663
rect 33517 17629 33551 17663
rect 33551 17629 33560 17663
rect 33508 17620 33560 17629
rect 34152 17663 34204 17672
rect 34152 17629 34161 17663
rect 34161 17629 34195 17663
rect 34195 17629 34204 17663
rect 34152 17620 34204 17629
rect 34796 17620 34848 17672
rect 37188 17663 37240 17672
rect 37188 17629 37197 17663
rect 37197 17629 37231 17663
rect 37231 17629 37240 17663
rect 37188 17620 37240 17629
rect 37832 17663 37884 17672
rect 37832 17629 37841 17663
rect 37841 17629 37875 17663
rect 37875 17629 37884 17663
rect 37832 17620 37884 17629
rect 14096 17484 14148 17536
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 18512 17484 18564 17536
rect 20076 17484 20128 17536
rect 22928 17484 22980 17536
rect 26332 17484 26384 17536
rect 27528 17484 27580 17536
rect 33416 17552 33468 17604
rect 32864 17484 32916 17536
rect 33508 17484 33560 17536
rect 35348 17484 35400 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 11152 17280 11204 17332
rect 19248 17280 19300 17332
rect 20444 17280 20496 17332
rect 8852 17255 8904 17264
rect 8852 17221 8861 17255
rect 8861 17221 8895 17255
rect 8895 17221 8904 17255
rect 8852 17212 8904 17221
rect 20076 17255 20128 17264
rect 20076 17221 20085 17255
rect 20085 17221 20119 17255
rect 20119 17221 20128 17255
rect 20076 17212 20128 17221
rect 21364 17212 21416 17264
rect 22468 17212 22520 17264
rect 22928 17255 22980 17264
rect 22928 17221 22937 17255
rect 22937 17221 22971 17255
rect 22971 17221 22980 17255
rect 22928 17212 22980 17221
rect 23848 17212 23900 17264
rect 26148 17280 26200 17332
rect 29184 17323 29236 17332
rect 29184 17289 29193 17323
rect 29193 17289 29227 17323
rect 29227 17289 29236 17323
rect 29184 17280 29236 17289
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 19248 17187 19300 17196
rect 8576 17076 8628 17128
rect 9036 17076 9088 17128
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 25688 17144 25740 17196
rect 30196 17212 30248 17264
rect 33508 17255 33560 17264
rect 33508 17221 33517 17255
rect 33517 17221 33551 17255
rect 33551 17221 33560 17255
rect 33508 17212 33560 17221
rect 35348 17255 35400 17264
rect 35348 17221 35357 17255
rect 35357 17221 35391 17255
rect 35391 17221 35400 17255
rect 35348 17212 35400 17221
rect 37464 17212 37516 17264
rect 19984 17119 20036 17128
rect 19984 17085 19993 17119
rect 19993 17085 20027 17119
rect 20027 17085 20036 17119
rect 19984 17076 20036 17085
rect 21456 17008 21508 17060
rect 24308 17008 24360 17060
rect 32036 17144 32088 17196
rect 30288 17076 30340 17128
rect 30564 17119 30616 17128
rect 30564 17085 30573 17119
rect 30573 17085 30607 17119
rect 30607 17085 30616 17119
rect 30564 17076 30616 17085
rect 32128 17076 32180 17128
rect 9772 16940 9824 16992
rect 20996 16940 21048 16992
rect 29920 16983 29972 16992
rect 29920 16949 29929 16983
rect 29929 16949 29963 16983
rect 29963 16949 29972 16983
rect 29920 16940 29972 16949
rect 30380 17008 30432 17060
rect 34612 17076 34664 17128
rect 35348 17076 35400 17128
rect 36084 17119 36136 17128
rect 36084 17085 36093 17119
rect 36093 17085 36127 17119
rect 36127 17085 36136 17119
rect 36084 17076 36136 17085
rect 36360 17076 36412 17128
rect 31116 16940 31168 16992
rect 33048 16940 33100 16992
rect 38200 17051 38252 17060
rect 38200 17017 38209 17051
rect 38209 17017 38243 17051
rect 38243 17017 38252 17051
rect 38200 17008 38252 17017
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19248 16736 19300 16788
rect 27436 16736 27488 16788
rect 28264 16736 28316 16788
rect 31024 16736 31076 16788
rect 34796 16736 34848 16788
rect 23664 16668 23716 16720
rect 13544 16600 13596 16652
rect 14464 16600 14516 16652
rect 20168 16600 20220 16652
rect 22744 16600 22796 16652
rect 23480 16600 23532 16652
rect 21180 16551 21181 16584
rect 21181 16551 21215 16584
rect 21215 16551 21232 16584
rect 21180 16532 21232 16551
rect 21548 16532 21600 16584
rect 22192 16464 22244 16516
rect 23204 16575 23256 16584
rect 23204 16541 23213 16575
rect 23213 16541 23247 16575
rect 23247 16541 23256 16575
rect 26332 16600 26384 16652
rect 28356 16668 28408 16720
rect 27344 16600 27396 16652
rect 29092 16600 29144 16652
rect 31392 16600 31444 16652
rect 34888 16668 34940 16720
rect 35716 16668 35768 16720
rect 35348 16600 35400 16652
rect 39396 16736 39448 16788
rect 23204 16532 23256 16541
rect 35992 16575 36044 16584
rect 35992 16541 36001 16575
rect 36001 16541 36035 16575
rect 36035 16541 36044 16575
rect 35992 16532 36044 16541
rect 38108 16668 38160 16720
rect 37004 16532 37056 16584
rect 39304 16600 39356 16652
rect 11888 16396 11940 16448
rect 20168 16396 20220 16448
rect 22652 16396 22704 16448
rect 23572 16396 23624 16448
rect 30288 16507 30340 16516
rect 30288 16473 30297 16507
rect 30297 16473 30331 16507
rect 30331 16473 30340 16507
rect 30288 16464 30340 16473
rect 31852 16507 31904 16516
rect 31852 16473 31861 16507
rect 31861 16473 31895 16507
rect 31895 16473 31904 16507
rect 32772 16507 32824 16516
rect 31852 16464 31904 16473
rect 32772 16473 32781 16507
rect 32781 16473 32815 16507
rect 32815 16473 32824 16507
rect 32772 16464 32824 16473
rect 32864 16464 32916 16516
rect 34336 16507 34388 16516
rect 34336 16473 34345 16507
rect 34345 16473 34379 16507
rect 34379 16473 34388 16507
rect 34336 16464 34388 16473
rect 27252 16396 27304 16448
rect 27620 16396 27672 16448
rect 29460 16396 29512 16448
rect 29828 16396 29880 16448
rect 37924 16532 37976 16584
rect 38752 16464 38804 16516
rect 35532 16396 35584 16448
rect 37648 16396 37700 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 13728 16192 13780 16244
rect 15016 16192 15068 16244
rect 17040 16167 17092 16176
rect 17040 16133 17049 16167
rect 17049 16133 17083 16167
rect 17083 16133 17092 16167
rect 17040 16124 17092 16133
rect 18512 16167 18564 16176
rect 18512 16133 18521 16167
rect 18521 16133 18555 16167
rect 18555 16133 18564 16167
rect 18512 16124 18564 16133
rect 18972 16192 19024 16244
rect 22100 16192 22152 16244
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 12256 15988 12308 16040
rect 17776 15988 17828 16040
rect 22376 16056 22428 16108
rect 25596 16192 25648 16244
rect 25320 16167 25372 16176
rect 25320 16133 25329 16167
rect 25329 16133 25363 16167
rect 25363 16133 25372 16167
rect 25320 16124 25372 16133
rect 20996 16031 21048 16040
rect 15108 15920 15160 15972
rect 17500 15963 17552 15972
rect 17500 15929 17509 15963
rect 17509 15929 17543 15963
rect 17543 15929 17552 15963
rect 17500 15920 17552 15929
rect 1768 15895 1820 15904
rect 1768 15861 1777 15895
rect 1777 15861 1811 15895
rect 1811 15861 1820 15895
rect 1768 15852 1820 15861
rect 12440 15852 12492 15904
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 22284 15988 22336 16040
rect 29828 16192 29880 16244
rect 30288 16192 30340 16244
rect 27804 16167 27856 16176
rect 27804 16133 27813 16167
rect 27813 16133 27847 16167
rect 27847 16133 27856 16167
rect 27804 16124 27856 16133
rect 27988 16124 28040 16176
rect 28448 16124 28500 16176
rect 29460 16167 29512 16176
rect 29460 16133 29469 16167
rect 29469 16133 29503 16167
rect 29503 16133 29512 16167
rect 29460 16124 29512 16133
rect 31576 16124 31628 16176
rect 35992 16192 36044 16244
rect 32680 16124 32732 16176
rect 34428 16167 34480 16176
rect 31024 16056 31076 16108
rect 34428 16133 34437 16167
rect 34437 16133 34471 16167
rect 34471 16133 34480 16167
rect 34428 16124 34480 16133
rect 34520 16124 34572 16176
rect 35624 16056 35676 16108
rect 37372 16124 37424 16176
rect 36728 16099 36780 16108
rect 36728 16065 36737 16099
rect 36737 16065 36771 16099
rect 36771 16065 36780 16099
rect 36728 16056 36780 16065
rect 38016 16099 38068 16108
rect 38016 16065 38025 16099
rect 38025 16065 38059 16099
rect 38059 16065 38068 16099
rect 38016 16056 38068 16065
rect 21272 15920 21324 15972
rect 23940 15920 23992 15972
rect 29460 15988 29512 16040
rect 29920 15988 29972 16040
rect 30380 15988 30432 16040
rect 33048 16031 33100 16040
rect 33048 15997 33057 16031
rect 33057 15997 33091 16031
rect 33091 15997 33100 16031
rect 33048 15988 33100 15997
rect 34520 15920 34572 15972
rect 37648 15920 37700 15972
rect 21180 15895 21232 15904
rect 21180 15861 21189 15895
rect 21189 15861 21223 15895
rect 21223 15861 21232 15895
rect 21180 15852 21232 15861
rect 24676 15852 24728 15904
rect 25964 15852 26016 15904
rect 26792 15852 26844 15904
rect 27436 15852 27488 15904
rect 30932 15852 30984 15904
rect 37096 15852 37148 15904
rect 38200 15895 38252 15904
rect 38200 15861 38209 15895
rect 38209 15861 38243 15895
rect 38243 15861 38252 15895
rect 38200 15852 38252 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 11704 15648 11756 15700
rect 24032 15648 24084 15700
rect 25228 15648 25280 15700
rect 26148 15648 26200 15700
rect 27804 15648 27856 15700
rect 29276 15648 29328 15700
rect 31024 15691 31076 15700
rect 31024 15657 31033 15691
rect 31033 15657 31067 15691
rect 31067 15657 31076 15691
rect 31024 15648 31076 15657
rect 34520 15648 34572 15700
rect 35624 15648 35676 15700
rect 13176 15512 13228 15564
rect 33048 15580 33100 15632
rect 8760 15444 8812 15496
rect 14556 15444 14608 15496
rect 16764 15444 16816 15496
rect 20628 15444 20680 15496
rect 22284 15444 22336 15496
rect 22468 15487 22520 15496
rect 22468 15453 22477 15487
rect 22477 15453 22511 15487
rect 22511 15453 22520 15487
rect 22468 15444 22520 15453
rect 22652 15487 22704 15496
rect 22652 15453 22661 15487
rect 22661 15453 22695 15487
rect 22695 15453 22704 15487
rect 22652 15444 22704 15453
rect 24216 15444 24268 15496
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 25964 15444 26016 15496
rect 26148 15487 26200 15496
rect 26148 15453 26157 15487
rect 26157 15453 26191 15487
rect 26191 15453 26200 15487
rect 27252 15487 27304 15496
rect 26148 15444 26200 15453
rect 27252 15453 27261 15487
rect 27261 15453 27295 15487
rect 27295 15453 27304 15487
rect 27252 15444 27304 15453
rect 28172 15444 28224 15496
rect 29184 15444 29236 15496
rect 30932 15444 30984 15496
rect 31208 15487 31260 15496
rect 31208 15453 31217 15487
rect 31217 15453 31251 15487
rect 31251 15453 31260 15487
rect 31208 15444 31260 15453
rect 31668 15487 31720 15496
rect 31668 15453 31677 15487
rect 31677 15453 31711 15487
rect 31711 15453 31720 15487
rect 31668 15444 31720 15453
rect 31852 15512 31904 15564
rect 31944 15444 31996 15496
rect 32772 15444 32824 15496
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 10324 15419 10376 15428
rect 10324 15385 10333 15419
rect 10333 15385 10367 15419
rect 10367 15385 10376 15419
rect 10324 15376 10376 15385
rect 10416 15419 10468 15428
rect 10416 15385 10425 15419
rect 10425 15385 10459 15419
rect 10459 15385 10468 15419
rect 10416 15376 10468 15385
rect 12716 15376 12768 15428
rect 17224 15376 17276 15428
rect 17500 15376 17552 15428
rect 23296 15376 23348 15428
rect 28448 15419 28500 15428
rect 28448 15385 28457 15419
rect 28457 15385 28491 15419
rect 28491 15385 28500 15419
rect 28448 15376 28500 15385
rect 28908 15376 28960 15428
rect 34152 15512 34204 15564
rect 36636 15512 36688 15564
rect 37556 15512 37608 15564
rect 35900 15444 35952 15496
rect 33692 15419 33744 15428
rect 33692 15385 33701 15419
rect 33701 15385 33735 15419
rect 33735 15385 33744 15419
rect 33692 15376 33744 15385
rect 36360 15419 36412 15428
rect 1768 15308 1820 15360
rect 16304 15308 16356 15360
rect 20536 15308 20588 15360
rect 21640 15308 21692 15360
rect 23112 15351 23164 15360
rect 23112 15317 23121 15351
rect 23121 15317 23155 15351
rect 23155 15317 23164 15351
rect 23112 15308 23164 15317
rect 23204 15308 23256 15360
rect 25412 15308 25464 15360
rect 27804 15308 27856 15360
rect 28172 15308 28224 15360
rect 30472 15351 30524 15360
rect 30472 15317 30481 15351
rect 30481 15317 30515 15351
rect 30515 15317 30524 15351
rect 30472 15308 30524 15317
rect 31116 15308 31168 15360
rect 32404 15351 32456 15360
rect 32404 15317 32413 15351
rect 32413 15317 32447 15351
rect 32447 15317 32456 15351
rect 32404 15308 32456 15317
rect 36360 15385 36369 15419
rect 36369 15385 36403 15419
rect 36403 15385 36412 15419
rect 36360 15376 36412 15385
rect 37648 15419 37700 15428
rect 37648 15385 37657 15419
rect 37657 15385 37691 15419
rect 37691 15385 37700 15419
rect 37648 15376 37700 15385
rect 37740 15308 37792 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 8116 15147 8168 15156
rect 8116 15113 8125 15147
rect 8125 15113 8159 15147
rect 8159 15113 8168 15147
rect 8116 15104 8168 15113
rect 12992 15104 13044 15156
rect 13636 15147 13688 15156
rect 13636 15113 13645 15147
rect 13645 15113 13679 15147
rect 13679 15113 13688 15147
rect 13636 15104 13688 15113
rect 17040 15104 17092 15156
rect 19984 15104 20036 15156
rect 23112 15104 23164 15156
rect 23388 15104 23440 15156
rect 28816 15104 28868 15156
rect 29000 15104 29052 15156
rect 35900 15147 35952 15156
rect 2044 15036 2096 15088
rect 7564 15036 7616 15088
rect 14372 15079 14424 15088
rect 14372 15045 14381 15079
rect 14381 15045 14415 15079
rect 14415 15045 14424 15079
rect 14372 15036 14424 15045
rect 15016 15036 15068 15088
rect 16672 15036 16724 15088
rect 16948 15079 17000 15088
rect 16948 15045 16957 15079
rect 16957 15045 16991 15079
rect 16991 15045 17000 15079
rect 16948 15036 17000 15045
rect 8024 15011 8076 15020
rect 8024 14977 8033 15011
rect 8033 14977 8067 15011
rect 8067 14977 8076 15011
rect 8024 14968 8076 14977
rect 9772 15011 9824 15020
rect 9772 14977 9781 15011
rect 9781 14977 9815 15011
rect 9815 14977 9824 15011
rect 9772 14968 9824 14977
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 17592 14968 17644 15020
rect 20168 14968 20220 15020
rect 30472 15036 30524 15088
rect 32220 15036 32272 15088
rect 23572 15011 23624 15020
rect 23572 14977 23581 15011
rect 23581 14977 23615 15011
rect 23615 14977 23624 15011
rect 23572 14968 23624 14977
rect 25044 15011 25096 15020
rect 25044 14977 25053 15011
rect 25053 14977 25087 15011
rect 25087 14977 25096 15011
rect 25044 14968 25096 14977
rect 26608 15011 26660 15020
rect 26608 14977 26617 15011
rect 26617 14977 26651 15011
rect 26651 14977 26660 15011
rect 26608 14968 26660 14977
rect 26884 14968 26936 15020
rect 27528 14968 27580 15020
rect 27712 14968 27764 15020
rect 15200 14900 15252 14952
rect 21548 14900 21600 14952
rect 28540 14943 28592 14952
rect 26884 14832 26936 14884
rect 28540 14909 28549 14943
rect 28549 14909 28583 14943
rect 28583 14909 28592 14943
rect 28540 14900 28592 14909
rect 29276 14968 29328 15020
rect 30288 14968 30340 15020
rect 32312 15011 32364 15020
rect 32312 14977 32321 15011
rect 32321 14977 32355 15011
rect 32355 14977 32364 15011
rect 32312 14968 32364 14977
rect 34612 15036 34664 15088
rect 34888 15036 34940 15088
rect 35900 15113 35909 15147
rect 35909 15113 35943 15147
rect 35943 15113 35952 15147
rect 35900 15104 35952 15113
rect 30840 14900 30892 14952
rect 31024 14943 31076 14952
rect 31024 14909 31033 14943
rect 31033 14909 31067 14943
rect 31067 14909 31076 14943
rect 31024 14900 31076 14909
rect 10784 14764 10836 14816
rect 24952 14764 25004 14816
rect 25044 14764 25096 14816
rect 30288 14832 30340 14884
rect 33968 14900 34020 14952
rect 29460 14764 29512 14816
rect 30564 14764 30616 14816
rect 34520 14900 34572 14952
rect 37004 14968 37056 15020
rect 38108 15011 38160 15020
rect 38108 14977 38117 15011
rect 38117 14977 38151 15011
rect 38151 14977 38160 15011
rect 38108 14968 38160 14977
rect 35624 14832 35676 14884
rect 31300 14764 31352 14816
rect 33692 14764 33744 14816
rect 34888 14764 34940 14816
rect 35808 14764 35860 14816
rect 35900 14764 35952 14816
rect 36912 14764 36964 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1860 14560 1912 14612
rect 7564 14560 7616 14612
rect 12072 14492 12124 14544
rect 20812 14560 20864 14612
rect 22744 14560 22796 14612
rect 25136 14560 25188 14612
rect 28448 14560 28500 14612
rect 28540 14560 28592 14612
rect 30288 14560 30340 14612
rect 31300 14560 31352 14612
rect 33692 14560 33744 14612
rect 36912 14560 36964 14612
rect 17868 14492 17920 14544
rect 21272 14492 21324 14544
rect 16948 14424 17000 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 8668 14356 8720 14408
rect 9036 14356 9088 14408
rect 14924 14399 14976 14408
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 15200 14356 15252 14408
rect 19432 14424 19484 14476
rect 20720 14424 20772 14476
rect 23296 14492 23348 14544
rect 26608 14492 26660 14544
rect 29736 14492 29788 14544
rect 30380 14492 30432 14544
rect 31024 14492 31076 14544
rect 21548 14467 21600 14476
rect 21548 14433 21557 14467
rect 21557 14433 21591 14467
rect 21591 14433 21600 14467
rect 21548 14424 21600 14433
rect 21824 14424 21876 14476
rect 23112 14424 23164 14476
rect 26700 14424 26752 14476
rect 26884 14424 26936 14476
rect 8852 14220 8904 14272
rect 11888 14220 11940 14272
rect 15292 14288 15344 14340
rect 17132 14288 17184 14340
rect 17592 14331 17644 14340
rect 17592 14297 17601 14331
rect 17601 14297 17635 14331
rect 17635 14297 17644 14331
rect 17592 14288 17644 14297
rect 16856 14220 16908 14272
rect 23664 14399 23716 14408
rect 23664 14365 23673 14399
rect 23673 14365 23707 14399
rect 23707 14365 23716 14399
rect 23664 14356 23716 14365
rect 26792 14356 26844 14408
rect 28448 14356 28500 14408
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 21640 14331 21692 14340
rect 21640 14297 21649 14331
rect 21649 14297 21683 14331
rect 21683 14297 21692 14331
rect 21640 14288 21692 14297
rect 21824 14288 21876 14340
rect 22376 14288 22428 14340
rect 22836 14288 22888 14340
rect 24860 14288 24912 14340
rect 27620 14331 27672 14340
rect 27620 14297 27629 14331
rect 27629 14297 27663 14331
rect 27663 14297 27672 14331
rect 28540 14331 28592 14340
rect 27620 14288 27672 14297
rect 28540 14297 28549 14331
rect 28549 14297 28583 14331
rect 28583 14297 28592 14331
rect 28540 14288 28592 14297
rect 30472 14331 30524 14340
rect 22928 14220 22980 14272
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 23572 14220 23624 14272
rect 24768 14220 24820 14272
rect 24952 14220 25004 14272
rect 30472 14297 30481 14331
rect 30481 14297 30515 14331
rect 30515 14297 30524 14331
rect 30472 14288 30524 14297
rect 30564 14331 30616 14340
rect 30564 14297 30573 14331
rect 30573 14297 30607 14331
rect 30607 14297 30616 14331
rect 30564 14288 30616 14297
rect 29460 14220 29512 14272
rect 30012 14220 30064 14272
rect 32404 14424 32456 14476
rect 37648 14492 37700 14544
rect 34152 14399 34204 14408
rect 34152 14365 34161 14399
rect 34161 14365 34195 14399
rect 34195 14365 34204 14399
rect 34152 14356 34204 14365
rect 34244 14356 34296 14408
rect 35348 14424 35400 14476
rect 36728 14424 36780 14476
rect 35900 14356 35952 14408
rect 36452 14399 36504 14408
rect 36452 14365 36461 14399
rect 36461 14365 36495 14399
rect 36495 14365 36504 14399
rect 36452 14356 36504 14365
rect 30840 14220 30892 14272
rect 35624 14288 35676 14340
rect 37280 14331 37332 14340
rect 37280 14297 37289 14331
rect 37289 14297 37323 14331
rect 37323 14297 37332 14331
rect 37280 14288 37332 14297
rect 38016 14220 38068 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9220 14016 9272 14068
rect 11888 13991 11940 14000
rect 11888 13957 11897 13991
rect 11897 13957 11931 13991
rect 11931 13957 11940 13991
rect 11888 13948 11940 13957
rect 17868 13991 17920 14000
rect 17868 13957 17877 13991
rect 17877 13957 17911 13991
rect 17911 13957 17920 13991
rect 17868 13948 17920 13957
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 10508 13880 10560 13932
rect 11060 13880 11112 13932
rect 13636 13880 13688 13932
rect 10324 13812 10376 13864
rect 10784 13812 10836 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 18420 13855 18472 13864
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 23020 14016 23072 14068
rect 30196 14059 30248 14068
rect 30196 14025 30205 14059
rect 30205 14025 30239 14059
rect 30239 14025 30248 14059
rect 30196 14016 30248 14025
rect 21180 13948 21232 14000
rect 22192 13991 22244 14000
rect 22192 13957 22201 13991
rect 22201 13957 22235 13991
rect 22235 13957 22244 13991
rect 22192 13948 22244 13957
rect 22928 13948 22980 14000
rect 24768 13991 24820 14000
rect 21824 13880 21876 13932
rect 23480 13880 23532 13932
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 20168 13855 20220 13864
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 23296 13812 23348 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 15844 13744 15896 13796
rect 21916 13744 21968 13796
rect 24768 13957 24777 13991
rect 24777 13957 24811 13991
rect 24811 13957 24820 13991
rect 24768 13948 24820 13957
rect 27804 13948 27856 14000
rect 30012 13948 30064 14000
rect 30564 13948 30616 14000
rect 29092 13880 29144 13932
rect 30104 13923 30156 13932
rect 30104 13889 30113 13923
rect 30113 13889 30147 13923
rect 30147 13889 30156 13923
rect 30104 13880 30156 13889
rect 34520 14059 34572 14068
rect 34520 14025 34529 14059
rect 34529 14025 34563 14059
rect 34563 14025 34572 14059
rect 34520 14016 34572 14025
rect 35808 13991 35860 14000
rect 32588 13923 32640 13932
rect 32588 13889 32597 13923
rect 32597 13889 32631 13923
rect 32631 13889 32640 13923
rect 32588 13880 32640 13889
rect 32772 13880 32824 13932
rect 35808 13957 35817 13991
rect 35817 13957 35851 13991
rect 35851 13957 35860 13991
rect 35808 13948 35860 13957
rect 36360 13880 36412 13932
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 27620 13812 27672 13864
rect 30380 13812 30432 13864
rect 31024 13855 31076 13864
rect 31024 13821 31033 13855
rect 31033 13821 31067 13855
rect 31067 13821 31076 13855
rect 31024 13812 31076 13821
rect 35716 13855 35768 13864
rect 35716 13821 35725 13855
rect 35725 13821 35759 13855
rect 35759 13821 35768 13855
rect 35716 13812 35768 13821
rect 35900 13812 35952 13864
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 18972 13719 19024 13728
rect 18972 13685 18981 13719
rect 18981 13685 19015 13719
rect 19015 13685 19024 13719
rect 18972 13676 19024 13685
rect 21180 13676 21232 13728
rect 26332 13676 26384 13728
rect 29276 13719 29328 13728
rect 29276 13685 29285 13719
rect 29285 13685 29319 13719
rect 29319 13685 29328 13719
rect 29276 13676 29328 13685
rect 31300 13676 31352 13728
rect 38200 13719 38252 13728
rect 38200 13685 38209 13719
rect 38209 13685 38243 13719
rect 38243 13685 38252 13719
rect 38200 13676 38252 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 14464 13472 14516 13524
rect 21088 13472 21140 13524
rect 28264 13472 28316 13524
rect 28448 13472 28500 13524
rect 28632 13472 28684 13524
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 11060 13379 11112 13388
rect 11060 13345 11069 13379
rect 11069 13345 11103 13379
rect 11103 13345 11112 13379
rect 18604 13404 18656 13456
rect 16948 13379 17000 13388
rect 11060 13336 11112 13345
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 17224 13379 17276 13388
rect 17224 13345 17233 13379
rect 17233 13345 17267 13379
rect 17267 13345 17276 13379
rect 17224 13336 17276 13345
rect 19984 13379 20036 13388
rect 19984 13345 19993 13379
rect 19993 13345 20027 13379
rect 20027 13345 20036 13379
rect 19984 13336 20036 13345
rect 26332 13379 26384 13388
rect 14832 13268 14884 13320
rect 22100 13268 22152 13320
rect 26332 13345 26341 13379
rect 26341 13345 26375 13379
rect 26375 13345 26384 13379
rect 26332 13336 26384 13345
rect 26700 13404 26752 13456
rect 30472 13472 30524 13524
rect 35808 13472 35860 13524
rect 38660 13472 38712 13524
rect 37556 13447 37608 13456
rect 29276 13336 29328 13388
rect 29460 13336 29512 13388
rect 31208 13379 31260 13388
rect 31208 13345 31217 13379
rect 31217 13345 31251 13379
rect 31251 13345 31260 13379
rect 31208 13336 31260 13345
rect 10876 13243 10928 13252
rect 10876 13209 10885 13243
rect 10885 13209 10919 13243
rect 10919 13209 10928 13243
rect 10876 13200 10928 13209
rect 17040 13243 17092 13252
rect 17040 13209 17049 13243
rect 17049 13209 17083 13243
rect 17083 13209 17092 13243
rect 17040 13200 17092 13209
rect 18144 13200 18196 13252
rect 13084 13132 13136 13184
rect 21640 13175 21692 13184
rect 21640 13141 21649 13175
rect 21649 13141 21683 13175
rect 21683 13141 21692 13175
rect 21640 13132 21692 13141
rect 22744 13175 22796 13184
rect 22744 13141 22753 13175
rect 22753 13141 22787 13175
rect 22787 13141 22796 13175
rect 22744 13132 22796 13141
rect 27160 13268 27212 13320
rect 31024 13268 31076 13320
rect 37556 13413 37565 13447
rect 37565 13413 37599 13447
rect 37599 13413 37608 13447
rect 37556 13404 37608 13413
rect 35348 13336 35400 13388
rect 32312 13311 32364 13320
rect 32312 13277 32321 13311
rect 32321 13277 32355 13311
rect 32355 13277 32364 13311
rect 32312 13268 32364 13277
rect 32956 13311 33008 13320
rect 32956 13277 32965 13311
rect 32965 13277 32999 13311
rect 32999 13277 33008 13311
rect 32956 13268 33008 13277
rect 33324 13268 33376 13320
rect 34520 13268 34572 13320
rect 30472 13200 30524 13252
rect 34796 13200 34848 13252
rect 35624 13200 35676 13252
rect 37004 13243 37056 13252
rect 37004 13209 37013 13243
rect 37013 13209 37047 13243
rect 37047 13209 37056 13243
rect 37004 13200 37056 13209
rect 37096 13243 37148 13252
rect 37096 13209 37105 13243
rect 37105 13209 37139 13243
rect 37139 13209 37148 13243
rect 37096 13200 37148 13209
rect 26976 13175 27028 13184
rect 26976 13141 26985 13175
rect 26985 13141 27019 13175
rect 27019 13141 27028 13175
rect 26976 13132 27028 13141
rect 29000 13132 29052 13184
rect 31300 13132 31352 13184
rect 34888 13175 34940 13184
rect 34888 13141 34897 13175
rect 34897 13141 34931 13175
rect 34931 13141 34940 13175
rect 34888 13132 34940 13141
rect 35532 13175 35584 13184
rect 35532 13141 35541 13175
rect 35541 13141 35575 13175
rect 35575 13141 35584 13175
rect 35532 13132 35584 13141
rect 36176 13175 36228 13184
rect 36176 13141 36185 13175
rect 36185 13141 36219 13175
rect 36219 13141 36228 13175
rect 36176 13132 36228 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1584 12928 1636 12980
rect 5448 12860 5500 12912
rect 10876 12860 10928 12912
rect 12256 12903 12308 12912
rect 12256 12869 12265 12903
rect 12265 12869 12299 12903
rect 12299 12869 12308 12903
rect 12256 12860 12308 12869
rect 18972 12860 19024 12912
rect 22744 12860 22796 12912
rect 24768 12860 24820 12912
rect 25044 12903 25096 12912
rect 25044 12869 25053 12903
rect 25053 12869 25087 12903
rect 25087 12869 25096 12903
rect 25044 12860 25096 12869
rect 29092 12928 29144 12980
rect 32588 12971 32640 12980
rect 32588 12937 32597 12971
rect 32597 12937 32631 12971
rect 32631 12937 32640 12971
rect 32588 12928 32640 12937
rect 32128 12860 32180 12912
rect 34888 12903 34940 12912
rect 4712 12792 4764 12844
rect 12164 12835 12216 12844
rect 12164 12801 12173 12835
rect 12173 12801 12207 12835
rect 12207 12801 12216 12835
rect 12164 12792 12216 12801
rect 15844 12792 15896 12844
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 23112 12792 23164 12844
rect 13084 12724 13136 12776
rect 17408 12724 17460 12776
rect 18420 12724 18472 12776
rect 14832 12699 14884 12708
rect 14832 12665 14841 12699
rect 14841 12665 14875 12699
rect 14875 12665 14884 12699
rect 14832 12656 14884 12665
rect 20168 12656 20220 12708
rect 23572 12767 23624 12776
rect 23572 12733 23581 12767
rect 23581 12733 23615 12767
rect 23615 12733 23624 12767
rect 23572 12724 23624 12733
rect 24676 12724 24728 12776
rect 22376 12699 22428 12708
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 4068 12631 4120 12640
rect 4068 12597 4077 12631
rect 4077 12597 4111 12631
rect 4111 12597 4120 12631
rect 4068 12588 4120 12597
rect 22376 12665 22385 12699
rect 22385 12665 22419 12699
rect 22419 12665 22428 12699
rect 22376 12656 22428 12665
rect 27620 12792 27672 12844
rect 28264 12835 28316 12844
rect 28264 12801 28273 12835
rect 28273 12801 28307 12835
rect 28307 12801 28316 12835
rect 28264 12792 28316 12801
rect 29000 12792 29052 12844
rect 31300 12792 31352 12844
rect 30380 12767 30432 12776
rect 29184 12656 29236 12708
rect 30380 12733 30389 12767
rect 30389 12733 30423 12767
rect 30423 12733 30432 12767
rect 30380 12724 30432 12733
rect 31208 12724 31260 12776
rect 31484 12792 31536 12844
rect 32312 12792 32364 12844
rect 33600 12792 33652 12844
rect 34888 12869 34897 12903
rect 34897 12869 34931 12903
rect 34931 12869 34940 12903
rect 34888 12860 34940 12869
rect 34980 12860 35032 12912
rect 35624 12860 35676 12912
rect 36176 12903 36228 12912
rect 36176 12869 36185 12903
rect 36185 12869 36219 12903
rect 36219 12869 36228 12903
rect 36176 12860 36228 12869
rect 37372 12792 37424 12844
rect 35532 12724 35584 12776
rect 35808 12724 35860 12776
rect 26976 12588 27028 12640
rect 31576 12588 31628 12640
rect 33048 12588 33100 12640
rect 36176 12588 36228 12640
rect 38200 12631 38252 12640
rect 38200 12597 38209 12631
rect 38209 12597 38243 12631
rect 38243 12597 38252 12631
rect 38200 12588 38252 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4896 12427 4948 12436
rect 4896 12393 4905 12427
rect 4905 12393 4939 12427
rect 4939 12393 4948 12427
rect 4896 12384 4948 12393
rect 16948 12384 17000 12436
rect 19892 12384 19944 12436
rect 31024 12384 31076 12436
rect 18604 12316 18656 12368
rect 24492 12316 24544 12368
rect 30656 12316 30708 12368
rect 31392 12316 31444 12368
rect 34520 12384 34572 12436
rect 34704 12384 34756 12436
rect 35348 12384 35400 12436
rect 37004 12384 37056 12436
rect 1492 12180 1544 12232
rect 13176 12180 13228 12232
rect 22008 12248 22060 12300
rect 23940 12291 23992 12300
rect 23940 12257 23949 12291
rect 23949 12257 23983 12291
rect 23983 12257 23992 12291
rect 23940 12248 23992 12257
rect 25228 12248 25280 12300
rect 29828 12291 29880 12300
rect 29828 12257 29837 12291
rect 29837 12257 29871 12291
rect 29871 12257 29880 12291
rect 29828 12248 29880 12257
rect 34704 12248 34756 12300
rect 35624 12291 35676 12300
rect 35624 12257 35633 12291
rect 35633 12257 35667 12291
rect 35667 12257 35676 12291
rect 35624 12248 35676 12257
rect 29644 12180 29696 12232
rect 22284 12112 22336 12164
rect 23204 12112 23256 12164
rect 24676 12155 24728 12164
rect 24676 12121 24685 12155
rect 24685 12121 24719 12155
rect 24719 12121 24728 12155
rect 24676 12112 24728 12121
rect 25688 12155 25740 12164
rect 20076 12044 20128 12096
rect 23664 12044 23716 12096
rect 25688 12121 25697 12155
rect 25697 12121 25731 12155
rect 25731 12121 25740 12155
rect 25688 12112 25740 12121
rect 26608 12044 26660 12096
rect 31116 12155 31168 12164
rect 31116 12121 31125 12155
rect 31125 12121 31159 12155
rect 31159 12121 31168 12155
rect 31116 12112 31168 12121
rect 31392 12112 31444 12164
rect 32956 12180 33008 12232
rect 32128 12087 32180 12096
rect 32128 12053 32137 12087
rect 32137 12053 32171 12087
rect 32171 12053 32180 12087
rect 32128 12044 32180 12053
rect 32220 12044 32272 12096
rect 35072 12155 35124 12164
rect 35072 12121 35081 12155
rect 35081 12121 35115 12155
rect 35115 12121 35124 12155
rect 39028 12180 39080 12232
rect 35072 12112 35124 12121
rect 37740 12112 37792 12164
rect 33232 12087 33284 12096
rect 33232 12053 33241 12087
rect 33241 12053 33275 12087
rect 33275 12053 33284 12087
rect 33232 12044 33284 12053
rect 34612 12044 34664 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 12624 11883 12676 11892
rect 12624 11849 12633 11883
rect 12633 11849 12667 11883
rect 12667 11849 12676 11883
rect 12624 11840 12676 11849
rect 17040 11840 17092 11892
rect 21456 11840 21508 11892
rect 16028 11772 16080 11824
rect 9036 11704 9088 11756
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 16764 11704 16816 11756
rect 18604 11815 18656 11824
rect 18604 11781 18613 11815
rect 18613 11781 18647 11815
rect 18647 11781 18656 11815
rect 18604 11772 18656 11781
rect 20076 11815 20128 11824
rect 20076 11781 20085 11815
rect 20085 11781 20119 11815
rect 20119 11781 20128 11815
rect 20076 11772 20128 11781
rect 20904 11772 20956 11824
rect 23756 11772 23808 11824
rect 25412 11815 25464 11824
rect 25412 11781 25421 11815
rect 25421 11781 25455 11815
rect 25455 11781 25464 11815
rect 25412 11772 25464 11781
rect 30380 11840 30432 11892
rect 32956 11883 33008 11892
rect 32956 11849 32965 11883
rect 32965 11849 32999 11883
rect 32999 11849 33008 11883
rect 32956 11840 33008 11849
rect 30748 11772 30800 11824
rect 30932 11772 30984 11824
rect 31576 11772 31628 11824
rect 31668 11772 31720 11824
rect 34520 11840 34572 11892
rect 35716 11840 35768 11892
rect 34428 11772 34480 11824
rect 18788 11636 18840 11688
rect 20076 11636 20128 11688
rect 27252 11636 27304 11688
rect 31300 11636 31352 11688
rect 24860 11568 24912 11620
rect 25872 11611 25924 11620
rect 25872 11577 25881 11611
rect 25881 11577 25915 11611
rect 25915 11577 25924 11611
rect 25872 11568 25924 11577
rect 30196 11568 30248 11620
rect 32220 11636 32272 11688
rect 33232 11704 33284 11756
rect 34612 11679 34664 11688
rect 34612 11645 34621 11679
rect 34621 11645 34655 11679
rect 34655 11645 34664 11679
rect 34612 11636 34664 11645
rect 35440 11704 35492 11756
rect 36452 11747 36504 11756
rect 36452 11713 36461 11747
rect 36461 11713 36495 11747
rect 36495 11713 36504 11747
rect 36452 11704 36504 11713
rect 37556 11704 37608 11756
rect 7564 11500 7616 11552
rect 9036 11500 9088 11552
rect 13544 11500 13596 11552
rect 21272 11500 21324 11552
rect 23480 11500 23532 11552
rect 27344 11500 27396 11552
rect 30748 11500 30800 11552
rect 33048 11568 33100 11620
rect 34796 11568 34848 11620
rect 32404 11543 32456 11552
rect 32404 11509 32413 11543
rect 32413 11509 32447 11543
rect 32447 11509 32456 11543
rect 32404 11500 32456 11509
rect 37832 11543 37884 11552
rect 37832 11509 37841 11543
rect 37841 11509 37875 11543
rect 37875 11509 37884 11543
rect 37832 11500 37884 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 9036 11296 9088 11348
rect 9128 11296 9180 11348
rect 10324 11296 10376 11348
rect 8576 11160 8628 11212
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 29644 11296 29696 11348
rect 31116 11296 31168 11348
rect 18788 11228 18840 11280
rect 20996 11228 21048 11280
rect 25688 11228 25740 11280
rect 35992 11296 36044 11348
rect 38016 11228 38068 11280
rect 21272 11203 21324 11212
rect 3424 11092 3476 11144
rect 7564 11135 7616 11144
rect 7564 11101 7573 11135
rect 7573 11101 7607 11135
rect 7607 11101 7616 11135
rect 7564 11092 7616 11101
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 1676 11067 1728 11076
rect 1676 11033 1685 11067
rect 1685 11033 1719 11067
rect 1719 11033 1728 11067
rect 1676 11024 1728 11033
rect 3976 11024 4028 11076
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 12992 11092 13044 11144
rect 14924 11092 14976 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 18144 11092 18196 11144
rect 22376 11160 22428 11212
rect 31300 11203 31352 11212
rect 31300 11169 31309 11203
rect 31309 11169 31343 11203
rect 31343 11169 31352 11203
rect 31300 11160 31352 11169
rect 37556 11160 37608 11212
rect 22100 11092 22152 11144
rect 30656 11135 30708 11144
rect 13360 11024 13412 11076
rect 22560 11024 22612 11076
rect 30656 11101 30665 11135
rect 30665 11101 30699 11135
rect 30699 11101 30708 11135
rect 30656 11092 30708 11101
rect 34796 11092 34848 11144
rect 36820 11135 36872 11144
rect 36820 11101 36829 11135
rect 36829 11101 36863 11135
rect 36863 11101 36872 11135
rect 36820 11092 36872 11101
rect 32128 11024 32180 11076
rect 36728 11024 36780 11076
rect 37556 11067 37608 11076
rect 37556 11033 37565 11067
rect 37565 11033 37599 11067
rect 37599 11033 37608 11067
rect 37556 11024 37608 11033
rect 37648 11067 37700 11076
rect 37648 11033 37657 11067
rect 37657 11033 37691 11067
rect 37691 11033 37700 11067
rect 37648 11024 37700 11033
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 28908 10999 28960 11008
rect 28908 10965 28917 10999
rect 28917 10965 28951 10999
rect 28951 10965 28960 10999
rect 28908 10956 28960 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4620 10752 4672 10804
rect 8944 10752 8996 10804
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 16028 10752 16080 10804
rect 24676 10752 24728 10804
rect 29828 10752 29880 10804
rect 36360 10752 36412 10804
rect 38200 10795 38252 10804
rect 38200 10761 38209 10795
rect 38209 10761 38243 10795
rect 38243 10761 38252 10795
rect 38200 10752 38252 10761
rect 14924 10684 14976 10736
rect 22560 10684 22612 10736
rect 27344 10727 27396 10736
rect 27344 10693 27353 10727
rect 27353 10693 27387 10727
rect 27387 10693 27396 10727
rect 27344 10684 27396 10693
rect 28356 10684 28408 10736
rect 35440 10684 35492 10736
rect 15200 10659 15252 10668
rect 15200 10625 15209 10659
rect 15209 10625 15243 10659
rect 15243 10625 15252 10659
rect 15200 10616 15252 10625
rect 15936 10616 15988 10668
rect 14280 10548 14332 10600
rect 22284 10616 22336 10668
rect 25228 10616 25280 10668
rect 28908 10659 28960 10668
rect 28908 10625 28917 10659
rect 28917 10625 28951 10659
rect 28951 10625 28960 10659
rect 28908 10616 28960 10625
rect 36176 10659 36228 10668
rect 27252 10591 27304 10600
rect 27252 10557 27261 10591
rect 27261 10557 27295 10591
rect 27295 10557 27304 10591
rect 29092 10591 29144 10600
rect 27252 10548 27304 10557
rect 16856 10480 16908 10532
rect 17776 10480 17828 10532
rect 25504 10480 25556 10532
rect 29092 10557 29101 10591
rect 29101 10557 29135 10591
rect 29135 10557 29144 10591
rect 29092 10548 29144 10557
rect 36176 10625 36185 10659
rect 36185 10625 36219 10659
rect 36219 10625 36228 10659
rect 36176 10616 36228 10625
rect 38016 10659 38068 10668
rect 38016 10625 38025 10659
rect 38025 10625 38059 10659
rect 38059 10625 38068 10659
rect 38016 10616 38068 10625
rect 38108 10548 38160 10600
rect 14648 10455 14700 10464
rect 14648 10421 14657 10455
rect 14657 10421 14691 10455
rect 14691 10421 14700 10455
rect 14648 10412 14700 10421
rect 16120 10412 16172 10464
rect 22652 10412 22704 10464
rect 24768 10412 24820 10464
rect 37924 10412 37976 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 17868 10208 17920 10260
rect 26240 10208 26292 10260
rect 30472 10251 30524 10260
rect 30472 10217 30481 10251
rect 30481 10217 30515 10251
rect 30515 10217 30524 10251
rect 30472 10208 30524 10217
rect 37372 10208 37424 10260
rect 38200 10251 38252 10260
rect 38200 10217 38209 10251
rect 38209 10217 38243 10251
rect 38243 10217 38252 10251
rect 38200 10208 38252 10217
rect 22468 10140 22520 10192
rect 22560 10115 22612 10124
rect 22560 10081 22569 10115
rect 22569 10081 22603 10115
rect 22603 10081 22612 10115
rect 22560 10072 22612 10081
rect 29828 10140 29880 10192
rect 10140 10004 10192 10056
rect 12440 10047 12492 10056
rect 12440 10013 12449 10047
rect 12449 10013 12483 10047
rect 12483 10013 12492 10047
rect 12440 10004 12492 10013
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 17776 10047 17828 10056
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 24952 10004 25004 10056
rect 30380 10047 30432 10056
rect 22652 9979 22704 9988
rect 22652 9945 22661 9979
rect 22661 9945 22695 9979
rect 22695 9945 22704 9979
rect 22652 9936 22704 9945
rect 2044 9868 2096 9920
rect 14924 9868 14976 9920
rect 17040 9868 17092 9920
rect 22192 9868 22244 9920
rect 24676 9936 24728 9988
rect 30380 10013 30389 10047
rect 30389 10013 30423 10047
rect 30423 10013 30432 10047
rect 30380 10004 30432 10013
rect 36912 10047 36964 10056
rect 36912 10013 36921 10047
rect 36921 10013 36955 10047
rect 36955 10013 36964 10047
rect 36912 10004 36964 10013
rect 37832 10004 37884 10056
rect 27712 9868 27764 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 12440 9707 12492 9716
rect 12440 9673 12449 9707
rect 12449 9673 12483 9707
rect 12483 9673 12492 9707
rect 12440 9664 12492 9673
rect 12624 9664 12676 9716
rect 15752 9707 15804 9716
rect 15752 9673 15761 9707
rect 15761 9673 15795 9707
rect 15795 9673 15804 9707
rect 15752 9664 15804 9673
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 15844 9596 15896 9648
rect 17040 9639 17092 9648
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 20996 9639 21048 9648
rect 20996 9605 21005 9639
rect 21005 9605 21039 9639
rect 21039 9605 21048 9639
rect 20996 9596 21048 9605
rect 20076 9528 20128 9580
rect 15936 9392 15988 9444
rect 1584 9324 1636 9376
rect 9128 9324 9180 9376
rect 17868 9460 17920 9512
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 22744 9596 22796 9648
rect 23480 9639 23532 9648
rect 23480 9605 23489 9639
rect 23489 9605 23523 9639
rect 23523 9605 23532 9639
rect 23480 9596 23532 9605
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 29092 9664 29144 9716
rect 27988 9596 28040 9648
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 24860 9571 24912 9580
rect 24860 9537 24869 9571
rect 24869 9537 24903 9571
rect 24903 9537 24912 9571
rect 24860 9528 24912 9537
rect 28908 9528 28960 9580
rect 37924 9571 37976 9580
rect 37924 9537 37933 9571
rect 37933 9537 37967 9571
rect 37967 9537 37976 9571
rect 37924 9528 37976 9537
rect 25964 9460 26016 9512
rect 25872 9392 25924 9444
rect 37280 9392 37332 9444
rect 20352 9324 20404 9376
rect 26884 9324 26936 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 20536 9120 20588 9172
rect 22468 9120 22520 9172
rect 14648 8984 14700 9036
rect 28356 8984 28408 9036
rect 30564 9027 30616 9036
rect 30564 8993 30573 9027
rect 30573 8993 30607 9027
rect 30607 8993 30616 9027
rect 30564 8984 30616 8993
rect 37556 9027 37608 9036
rect 37556 8993 37565 9027
rect 37565 8993 37599 9027
rect 37599 8993 37608 9027
rect 37556 8984 37608 8993
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 12440 8916 12492 8968
rect 20352 8959 20404 8968
rect 20352 8925 20361 8959
rect 20361 8925 20395 8959
rect 20395 8925 20404 8959
rect 20352 8916 20404 8925
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 25504 8916 25556 8968
rect 32404 8916 32456 8968
rect 24768 8891 24820 8900
rect 24768 8857 24777 8891
rect 24777 8857 24811 8891
rect 24811 8857 24820 8891
rect 30104 8891 30156 8900
rect 24768 8848 24820 8857
rect 30104 8857 30113 8891
rect 30113 8857 30147 8891
rect 30147 8857 30156 8891
rect 30104 8848 30156 8857
rect 30288 8848 30340 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 27712 8780 27764 8832
rect 33600 8780 33652 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 17408 8576 17460 8628
rect 28908 8619 28960 8628
rect 28908 8585 28917 8619
rect 28917 8585 28951 8619
rect 28951 8585 28960 8619
rect 28908 8576 28960 8585
rect 30104 8619 30156 8628
rect 30104 8585 30113 8619
rect 30113 8585 30147 8619
rect 30147 8585 30156 8619
rect 30104 8576 30156 8585
rect 38108 8619 38160 8628
rect 38108 8585 38117 8619
rect 38117 8585 38151 8619
rect 38151 8585 38160 8619
rect 38108 8576 38160 8585
rect 22192 8551 22244 8560
rect 22192 8517 22201 8551
rect 22201 8517 22235 8551
rect 22235 8517 22244 8551
rect 22192 8508 22244 8517
rect 22744 8551 22796 8560
rect 22744 8517 22753 8551
rect 22753 8517 22787 8551
rect 22787 8517 22796 8551
rect 22744 8508 22796 8517
rect 27712 8551 27764 8560
rect 27712 8517 27721 8551
rect 27721 8517 27755 8551
rect 27755 8517 27764 8551
rect 27712 8508 27764 8517
rect 28356 8508 28408 8560
rect 4620 8440 4672 8492
rect 24860 8440 24912 8492
rect 27712 8372 27764 8424
rect 29368 8440 29420 8492
rect 38292 8483 38344 8492
rect 38292 8449 38301 8483
rect 38301 8449 38335 8483
rect 38335 8449 38344 8483
rect 38292 8440 38344 8449
rect 26516 8279 26568 8288
rect 26516 8245 26525 8279
rect 26525 8245 26559 8279
rect 26559 8245 26568 8279
rect 26516 8236 26568 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8024 8032 8076 8084
rect 9128 8032 9180 8084
rect 11520 8032 11572 8084
rect 32404 8032 32456 8084
rect 27712 8007 27764 8016
rect 27712 7973 27721 8007
rect 27721 7973 27755 8007
rect 27755 7973 27764 8007
rect 27712 7964 27764 7973
rect 38384 7964 38436 8016
rect 23204 7896 23256 7948
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 20996 7828 21048 7880
rect 27160 7828 27212 7880
rect 32404 7871 32456 7880
rect 32404 7837 32413 7871
rect 32413 7837 32447 7871
rect 32447 7837 32456 7871
rect 32404 7828 32456 7837
rect 37464 7871 37516 7880
rect 37464 7837 37473 7871
rect 37473 7837 37507 7871
rect 37507 7837 37516 7871
rect 37464 7828 37516 7837
rect 31392 7803 31444 7812
rect 31392 7769 31401 7803
rect 31401 7769 31435 7803
rect 31435 7769 31444 7803
rect 31392 7760 31444 7769
rect 27804 7692 27856 7744
rect 34336 7692 34388 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 26608 7531 26660 7540
rect 26608 7497 26617 7531
rect 26617 7497 26651 7531
rect 26651 7497 26660 7531
rect 26608 7488 26660 7497
rect 37740 7488 37792 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 22284 7352 22336 7404
rect 23204 7352 23256 7404
rect 24860 7352 24912 7404
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 26516 7352 26568 7404
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 6552 7216 6604 7268
rect 9128 7148 9180 7200
rect 24768 7148 24820 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12440 6808 12492 6860
rect 26608 6808 26660 6860
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 24768 6783 24820 6792
rect 24768 6749 24777 6783
rect 24777 6749 24811 6783
rect 24811 6749 24820 6783
rect 24768 6740 24820 6749
rect 30564 6808 30616 6860
rect 31668 6808 31720 6860
rect 30472 6715 30524 6724
rect 30472 6681 30481 6715
rect 30481 6681 30515 6715
rect 30515 6681 30524 6715
rect 30472 6672 30524 6681
rect 30840 6672 30892 6724
rect 29828 6647 29880 6656
rect 29828 6613 29837 6647
rect 29837 6613 29871 6647
rect 29871 6613 29880 6647
rect 29828 6604 29880 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 12440 6264 12492 6316
rect 23296 6264 23348 6316
rect 29828 6264 29880 6316
rect 23388 6060 23440 6112
rect 26332 6060 26384 6112
rect 31668 6060 31720 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1492 5856 1544 5908
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 26332 5695 26384 5704
rect 26332 5661 26341 5695
rect 26341 5661 26375 5695
rect 26375 5661 26384 5695
rect 26332 5652 26384 5661
rect 14004 5584 14056 5636
rect 28908 5516 28960 5568
rect 38200 5559 38252 5568
rect 38200 5525 38209 5559
rect 38209 5525 38243 5559
rect 38243 5525 38252 5559
rect 38200 5516 38252 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 18696 5312 18748 5364
rect 25964 5312 26016 5364
rect 30472 5312 30524 5364
rect 27620 5176 27672 5228
rect 37740 5108 37792 5160
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 37740 4675 37792 4684
rect 37740 4641 37749 4675
rect 37749 4641 37783 4675
rect 37783 4641 37792 4675
rect 37740 4632 37792 4641
rect 36728 4564 36780 4616
rect 37464 4607 37516 4616
rect 37464 4573 37473 4607
rect 37473 4573 37507 4607
rect 37507 4573 37516 4607
rect 37464 4564 37516 4573
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 36728 4088 36780 4140
rect 35900 3884 35952 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 36728 3723 36780 3732
rect 36728 3689 36737 3723
rect 36737 3689 36771 3723
rect 36771 3689 36780 3723
rect 36728 3680 36780 3689
rect 1860 3476 1912 3528
rect 37740 3544 37792 3596
rect 35992 3408 36044 3460
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 38200 3383 38252 3392
rect 38200 3349 38209 3383
rect 38209 3349 38243 3383
rect 38243 3349 38252 3383
rect 38200 3340 38252 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3424 3136 3476 3188
rect 4620 3136 4672 3188
rect 22928 3136 22980 3188
rect 36452 3136 36504 3188
rect 21640 3068 21692 3120
rect 2780 3000 2832 3052
rect 2872 3000 2924 3052
rect 3884 3000 3936 3052
rect 8208 3000 8260 3052
rect 12992 3000 13044 3052
rect 16764 3000 16816 3052
rect 22560 3000 22612 3052
rect 28908 3000 28960 3052
rect 35440 3043 35492 3052
rect 35440 3009 35449 3043
rect 35449 3009 35483 3043
rect 35483 3009 35492 3043
rect 35440 3000 35492 3009
rect 9036 2864 9088 2916
rect 31392 2932 31444 2984
rect 31576 2932 31628 2984
rect 35992 3043 36044 3052
rect 35992 3009 36001 3043
rect 36001 3009 36035 3043
rect 36035 3009 36044 3043
rect 35992 3000 36044 3009
rect 37372 3000 37424 3052
rect 30380 2864 30432 2916
rect 664 2796 716 2848
rect 5356 2839 5408 2848
rect 5356 2805 5365 2839
rect 5365 2805 5399 2839
rect 5399 2805 5408 2839
rect 5356 2796 5408 2805
rect 30288 2796 30340 2848
rect 38660 2796 38712 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8208 2592 8260 2644
rect 12532 2592 12584 2644
rect 20 2524 72 2576
rect 13176 2592 13228 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20260 2592 20312 2644
rect 22100 2592 22152 2644
rect 24676 2592 24728 2644
rect 27160 2635 27212 2644
rect 27160 2601 27169 2635
rect 27169 2601 27203 2635
rect 27203 2601 27212 2635
rect 27160 2592 27212 2601
rect 1952 2388 2004 2440
rect 5356 2456 5408 2508
rect 12164 2456 12216 2508
rect 22652 2524 22704 2576
rect 16672 2456 16724 2508
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 31208 2499 31260 2508
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4068 2388 4120 2440
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 7104 2388 7156 2440
rect 8392 2388 8444 2440
rect 9680 2388 9732 2440
rect 10324 2388 10376 2440
rect 11612 2388 11664 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13544 2388 13596 2440
rect 14832 2388 14884 2440
rect 16120 2388 16172 2440
rect 18052 2388 18104 2440
rect 19340 2388 19392 2440
rect 19984 2388 20036 2440
rect 13360 2320 13412 2372
rect 31208 2465 31217 2499
rect 31217 2465 31251 2499
rect 31251 2465 31260 2499
rect 31208 2456 31260 2465
rect 32036 2456 32088 2508
rect 34336 2456 34388 2508
rect 21272 2388 21324 2440
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 1952 2252 2004 2304
rect 3240 2252 3292 2304
rect 5172 2252 5224 2304
rect 6460 2252 6512 2304
rect 12440 2252 12492 2304
rect 12992 2252 13044 2304
rect 24492 2388 24544 2440
rect 25780 2388 25832 2440
rect 27068 2388 27120 2440
rect 27804 2431 27856 2440
rect 27804 2397 27813 2431
rect 27813 2397 27847 2431
rect 27847 2397 27856 2431
rect 27804 2388 27856 2397
rect 29736 2431 29788 2440
rect 29736 2397 29745 2431
rect 29745 2397 29779 2431
rect 29779 2397 29788 2431
rect 29736 2388 29788 2397
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 32220 2388 32272 2440
rect 33600 2431 33652 2440
rect 33600 2397 33609 2431
rect 33609 2397 33643 2431
rect 33643 2397 33652 2431
rect 33600 2388 33652 2397
rect 31668 2320 31720 2372
rect 35900 2431 35952 2440
rect 35900 2397 35909 2431
rect 35909 2397 35943 2431
rect 35943 2397 35952 2431
rect 35900 2388 35952 2397
rect 27620 2252 27672 2304
rect 27712 2252 27764 2304
rect 29000 2252 29052 2304
rect 33508 2252 33560 2304
rect 34152 2252 34204 2304
rect 37188 2320 37240 2372
rect 36820 2295 36872 2304
rect 36820 2261 36829 2295
rect 36829 2261 36863 2295
rect 36863 2261 36872 2295
rect 36820 2252 36872 2261
rect 37096 2252 37148 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 1950 39200 2006 39800
rect 2594 39200 2650 39800
rect 3422 39536 3478 39545
rect 3422 39471 3478 39480
rect 676 35154 704 39200
rect 1964 37330 1992 39200
rect 1952 37324 2004 37330
rect 1952 37266 2004 37272
rect 2136 37256 2188 37262
rect 2136 37198 2188 37204
rect 1584 36644 1636 36650
rect 1584 36586 1636 36592
rect 1596 36281 1624 36586
rect 1582 36272 1638 36281
rect 1582 36207 1584 36216
rect 1636 36207 1638 36216
rect 1584 36178 1636 36184
rect 1398 36136 1454 36145
rect 1398 36071 1454 36080
rect 1768 36100 1820 36106
rect 664 35148 716 35154
rect 664 35090 716 35096
rect 1412 35086 1440 36071
rect 1768 36042 1820 36048
rect 1780 35834 1808 36042
rect 1768 35828 1820 35834
rect 1768 35770 1820 35776
rect 1492 35692 1544 35698
rect 1492 35634 1544 35640
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1504 19786 1532 35634
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34105 1808 34342
rect 1766 34096 1822 34105
rect 1766 34031 1822 34040
rect 2148 33998 2176 37198
rect 2228 36848 2280 36854
rect 2228 36790 2280 36796
rect 2240 34746 2268 36790
rect 2608 36768 2636 39200
rect 2870 38856 2926 38865
rect 2870 38791 2926 38800
rect 2884 38350 2912 38791
rect 2872 38344 2924 38350
rect 2872 38286 2924 38292
rect 2870 37496 2926 37505
rect 2870 37431 2926 37440
rect 2780 36780 2832 36786
rect 2608 36740 2780 36768
rect 2780 36722 2832 36728
rect 2780 36576 2832 36582
rect 2780 36518 2832 36524
rect 2320 35692 2372 35698
rect 2320 35634 2372 35640
rect 2332 35601 2360 35634
rect 2318 35592 2374 35601
rect 2318 35527 2374 35536
rect 2228 34740 2280 34746
rect 2228 34682 2280 34688
rect 2320 34604 2372 34610
rect 2320 34546 2372 34552
rect 2136 33992 2188 33998
rect 2332 33969 2360 34546
rect 2792 33998 2820 36518
rect 2884 35562 2912 37431
rect 3436 37262 3464 39471
rect 3882 39200 3938 39800
rect 5170 39200 5226 39800
rect 5814 39200 5870 39800
rect 7102 39200 7158 39800
rect 8390 39200 8446 39800
rect 9034 39200 9090 39800
rect 10322 39200 10378 39800
rect 11610 39200 11666 39800
rect 12254 39200 12310 39800
rect 13542 39200 13598 39800
rect 14830 39200 14886 39800
rect 14936 39222 15148 39250
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3896 36768 3924 39200
rect 4620 38344 4672 38350
rect 4620 38286 4672 38292
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4160 36780 4212 36786
rect 3896 36740 4160 36768
rect 4160 36722 4212 36728
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 38286
rect 4896 37324 4948 37330
rect 4896 37266 4948 37272
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 3056 35760 3108 35766
rect 3054 35728 3056 35737
rect 3976 35760 4028 35766
rect 3108 35728 3110 35737
rect 3976 35702 4028 35708
rect 3054 35663 3110 35672
rect 2872 35556 2924 35562
rect 2872 35498 2924 35504
rect 3988 34678 4016 35702
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 3884 34604 3936 34610
rect 3884 34546 3936 34552
rect 2780 33992 2832 33998
rect 2136 33934 2188 33940
rect 2318 33960 2374 33969
rect 1584 33856 1636 33862
rect 1584 33798 1636 33804
rect 1596 32910 1624 33798
rect 1584 32904 1636 32910
rect 1584 32846 1636 32852
rect 1768 32768 1820 32774
rect 1766 32736 1768 32745
rect 1820 32736 1822 32745
rect 1766 32671 1822 32680
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 1768 32224 1820 32230
rect 1768 32166 1820 32172
rect 1780 32065 1808 32166
rect 1766 32056 1822 32065
rect 1766 31991 1822 32000
rect 1766 30696 1822 30705
rect 1766 30631 1822 30640
rect 1780 30598 1808 30631
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1860 29640 1912 29646
rect 1860 29582 1912 29588
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1780 29345 1808 29446
rect 1766 29336 1822 29345
rect 1766 29271 1822 29280
rect 1584 29096 1636 29102
rect 1584 29038 1636 29044
rect 1596 28665 1624 29038
rect 1582 28656 1638 28665
rect 1582 28591 1638 28600
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 1688 27305 1716 27338
rect 1674 27296 1730 27305
rect 1674 27231 1730 27240
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1780 25945 1808 26318
rect 1766 25936 1822 25945
rect 1766 25871 1822 25880
rect 1768 24608 1820 24614
rect 1766 24576 1768 24585
rect 1820 24576 1822 24585
rect 1766 24511 1822 24520
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 1596 23905 1624 24142
rect 1582 23896 1638 23905
rect 1582 23831 1638 23840
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22545 1808 22578
rect 1766 22536 1822 22545
rect 1766 22471 1822 22480
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1688 21185 1716 21490
rect 1674 21176 1730 21185
rect 1674 21111 1730 21120
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1688 20505 1716 20810
rect 1872 20602 1900 29582
rect 1952 29096 2004 29102
rect 1952 29038 2004 29044
rect 1964 23730 1992 29038
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1964 21554 1992 23666
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1674 20496 1730 20505
rect 1674 20431 1730 20440
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1872 19922 1900 20402
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1492 19780 1544 19786
rect 1492 19722 1544 19728
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1780 19145 1808 19314
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 1596 17785 1624 18158
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 17105 1808 17138
rect 1766 17096 1822 17105
rect 1766 17031 1822 17040
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1780 15745 1808 15846
rect 1766 15736 1822 15745
rect 1766 15671 1822 15680
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 14498 1808 15302
rect 1872 14618 1900 19858
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1780 14470 1900 14498
rect 1768 14408 1820 14414
rect 1766 14376 1768 14385
rect 1820 14376 1822 14385
rect 1766 14311 1822 14320
rect 1584 13932 1636 13938
rect 1584 13874 1636 13880
rect 1596 12986 1624 13874
rect 1768 13728 1820 13734
rect 1766 13696 1768 13705
rect 1820 13696 1822 13705
rect 1766 13631 1822 13640
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12345 1808 12582
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 5914 1532 12174
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1688 10985 1716 11018
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1780 10305 1808 10610
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8974 1624 9318
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1766 8936 1822 8945
rect 1766 8871 1822 8880
rect 1780 8838 1808 8871
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7585 1808 7822
rect 1766 7576 1822 7585
rect 1766 7511 1822 7520
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1780 6905 1808 7346
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1780 5545 1808 5646
rect 1766 5536 1822 5545
rect 1766 5471 1822 5480
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 4185 1808 4422
rect 1766 4176 1822 4185
rect 1766 4111 1822 4120
rect 1872 3534 1900 14470
rect 1860 3528 1912 3534
rect 1766 3496 1822 3505
rect 1860 3470 1912 3476
rect 1766 3431 1822 3440
rect 1780 3398 1808 3431
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 20 2576 72 2582
rect 20 2518 72 2524
rect 32 800 60 2518
rect 676 800 704 2790
rect 1964 2446 1992 21286
rect 2056 15094 2084 32370
rect 2148 29782 2176 33934
rect 2780 33934 2832 33940
rect 2318 33895 2374 33904
rect 2872 33856 2924 33862
rect 2872 33798 2924 33804
rect 2136 29776 2188 29782
rect 2136 29718 2188 29724
rect 2884 25362 2912 33798
rect 3896 33114 3924 34546
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3884 33108 3936 33114
rect 3884 33050 3936 33056
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 31482 4660 33526
rect 4620 31476 4672 31482
rect 4620 31418 4672 31424
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4724 29306 4752 30670
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27674 4660 28494
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 4632 24818 4660 27610
rect 4908 26874 4936 37266
rect 5184 37262 5212 39200
rect 5828 37262 5856 39200
rect 7116 37262 7144 39200
rect 8404 37330 8432 39200
rect 8392 37324 8444 37330
rect 8392 37266 8444 37272
rect 9048 37262 9076 39200
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 9496 37256 9548 37262
rect 9496 37198 9548 37204
rect 8116 37188 8168 37194
rect 8116 37130 8168 37136
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 6644 37120 6696 37126
rect 6644 37062 6696 37068
rect 7196 37120 7248 37126
rect 7196 37062 7248 37068
rect 5448 36100 5500 36106
rect 5448 36042 5500 36048
rect 4988 34944 5040 34950
rect 4988 34886 5040 34892
rect 5000 34610 5028 34886
rect 5460 34746 5488 36042
rect 5448 34740 5500 34746
rect 5448 34682 5500 34688
rect 4988 34604 5040 34610
rect 4988 34546 5040 34552
rect 5080 33448 5132 33454
rect 5080 33390 5132 33396
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5092 32978 5120 33390
rect 5080 32972 5132 32978
rect 5080 32914 5132 32920
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 5000 28014 5028 28358
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 4908 26846 5028 26874
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 3988 23594 4016 24754
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3976 23588 4028 23594
rect 3976 23530 4028 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22166 4660 22510
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 2044 15088 2096 15094
rect 2044 15030 2096 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9586 2084 9862
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 3436 3194 3464 11086
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1964 800 1992 2246
rect 2792 2145 2820 2994
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 18 200 74 800
rect 662 200 718 800
rect 1950 200 2006 800
rect 2884 785 2912 2994
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 800 3280 2246
rect 3896 800 3924 2994
rect 3988 2446 4016 11018
rect 4080 2446 4108 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 10810 4660 18226
rect 4724 12850 4752 26318
rect 4896 24132 4948 24138
rect 4896 24074 4948 24080
rect 4804 22024 4856 22030
rect 4804 21966 4856 21972
rect 4816 21690 4844 21966
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4908 12442 4936 24074
rect 5000 22094 5028 26846
rect 5276 26042 5304 31282
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 5092 24954 5120 25230
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 5000 22066 5120 22094
rect 5092 20262 5120 22066
rect 5368 20602 5396 33390
rect 6380 31278 6408 37062
rect 6552 35692 6604 35698
rect 6552 35634 6604 35640
rect 6564 35290 6592 35634
rect 6552 35284 6604 35290
rect 6552 35226 6604 35232
rect 6458 35184 6514 35193
rect 6458 35119 6514 35128
rect 6472 35086 6500 35119
rect 6460 35080 6512 35086
rect 6460 35022 6512 35028
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6564 34678 6592 34886
rect 6552 34672 6604 34678
rect 6552 34614 6604 34620
rect 6656 31346 6684 37062
rect 7208 36786 7236 37062
rect 8128 36786 8156 37130
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 7196 36780 7248 36786
rect 7196 36722 7248 36728
rect 8116 36780 8168 36786
rect 8116 36722 8168 36728
rect 8484 36780 8536 36786
rect 8484 36722 8536 36728
rect 8668 36780 8720 36786
rect 8668 36722 8720 36728
rect 8022 36680 8078 36689
rect 8022 36615 8024 36624
rect 8076 36615 8078 36624
rect 8024 36586 8076 36592
rect 8496 36378 8524 36722
rect 8680 36378 8708 36722
rect 8484 36372 8536 36378
rect 8484 36314 8536 36320
rect 8668 36372 8720 36378
rect 8668 36314 8720 36320
rect 6736 36168 6788 36174
rect 6734 36136 6736 36145
rect 6788 36136 6790 36145
rect 6734 36071 6790 36080
rect 6736 36032 6788 36038
rect 6736 35974 6788 35980
rect 8024 36032 8076 36038
rect 8024 35974 8076 35980
rect 9036 36032 9088 36038
rect 9036 35974 9088 35980
rect 6748 33454 6776 35974
rect 6920 35216 6972 35222
rect 6920 35158 6972 35164
rect 6932 33998 6960 35158
rect 6920 33992 6972 33998
rect 6920 33934 6972 33940
rect 8036 33590 8064 35974
rect 8300 35828 8352 35834
rect 8300 35770 8352 35776
rect 8312 34610 8340 35770
rect 8576 35692 8628 35698
rect 8576 35634 8628 35640
rect 8588 35562 8616 35634
rect 8668 35624 8720 35630
rect 8668 35566 8720 35572
rect 8576 35556 8628 35562
rect 8576 35498 8628 35504
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 8300 34604 8352 34610
rect 8300 34546 8352 34552
rect 8220 33833 8248 34546
rect 8206 33824 8262 33833
rect 8128 33782 8206 33810
rect 8024 33584 8076 33590
rect 8024 33526 8076 33532
rect 6736 33448 6788 33454
rect 6736 33390 6788 33396
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 7300 32502 7328 32710
rect 7288 32496 7340 32502
rect 7288 32438 7340 32444
rect 7196 32360 7248 32366
rect 7196 32302 7248 32308
rect 7208 31482 7236 32302
rect 7196 31476 7248 31482
rect 7196 31418 7248 31424
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 6368 31272 6420 31278
rect 6368 31214 6420 31220
rect 7748 29572 7800 29578
rect 7748 29514 7800 29520
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6840 28762 6868 29106
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7564 28552 7616 28558
rect 7564 28494 7616 28500
rect 7208 27674 7236 28494
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7104 27668 7156 27674
rect 7104 27610 7156 27616
rect 7196 27668 7248 27674
rect 7196 27610 7248 27616
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 5460 26382 5488 27338
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6000 26920 6052 26926
rect 6000 26862 6052 26868
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 5448 26240 5500 26246
rect 5448 26182 5500 26188
rect 5460 25906 5488 26182
rect 5448 25900 5500 25906
rect 5448 25842 5500 25848
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 5552 24682 5580 25774
rect 6012 25702 6040 26862
rect 6840 26450 6868 26998
rect 7024 26994 7052 27270
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7116 26790 7144 27610
rect 7208 26858 7236 27610
rect 7484 27470 7512 28018
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7196 26852 7248 26858
rect 7196 26794 7248 26800
rect 7104 26784 7156 26790
rect 7104 26726 7156 26732
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5540 24676 5592 24682
rect 5540 24618 5592 24624
rect 5644 21894 5672 25094
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 5828 24274 5856 24754
rect 6012 24682 6040 25638
rect 6840 24818 6868 26386
rect 7116 25906 7144 26726
rect 7576 26586 7604 28494
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 7576 24818 7604 25638
rect 7760 24818 7788 29514
rect 8036 29238 8064 33526
rect 8024 29232 8076 29238
rect 8024 29174 8076 29180
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7852 27538 7880 27814
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7944 27470 7972 27814
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 6000 24676 6052 24682
rect 6000 24618 6052 24624
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 5816 24268 5868 24274
rect 5816 24210 5868 24216
rect 6276 24132 6328 24138
rect 6276 24074 6328 24080
rect 6288 23866 6316 24074
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6748 23730 6776 24550
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 7300 22778 7328 24142
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5644 20398 5672 21830
rect 7576 20874 7604 21830
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 6656 20058 6684 20470
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5460 12918 5488 19926
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6840 19514 6868 19790
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 7300 17746 7328 20334
rect 7484 18426 7512 20810
rect 7668 19514 7696 21490
rect 7852 20466 7880 25638
rect 7944 25498 7972 27406
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7748 20324 7800 20330
rect 7748 20266 7800 20272
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7760 19378 7788 20266
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 7760 18766 7788 19314
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7944 18222 7972 24754
rect 8036 24614 8064 25298
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 8036 21962 8064 24550
rect 8128 23118 8156 33782
rect 8206 33759 8262 33768
rect 8680 33522 8708 35566
rect 9048 33658 9076 35974
rect 9036 33652 9088 33658
rect 9036 33594 9088 33600
rect 8668 33516 8720 33522
rect 8496 33476 8668 33504
rect 8208 33108 8260 33114
rect 8208 33050 8260 33056
rect 8220 30258 8248 33050
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8404 30938 8432 32846
rect 8392 30932 8444 30938
rect 8392 30874 8444 30880
rect 8404 30394 8432 30874
rect 8392 30388 8444 30394
rect 8392 30330 8444 30336
rect 8208 30252 8260 30258
rect 8208 30194 8260 30200
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 8312 25294 8340 26250
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8404 24342 8432 28426
rect 8392 24336 8444 24342
rect 8392 24278 8444 24284
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8312 23798 8340 24006
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 8404 23254 8432 24278
rect 8392 23248 8444 23254
rect 8392 23190 8444 23196
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8404 22030 8432 22714
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 8496 21010 8524 33476
rect 8668 33458 8720 33464
rect 9140 31822 9168 37062
rect 9312 36576 9364 36582
rect 9312 36518 9364 36524
rect 9404 36576 9456 36582
rect 9404 36518 9456 36524
rect 9324 35154 9352 36518
rect 9416 36038 9444 36518
rect 9404 36032 9456 36038
rect 9404 35974 9456 35980
rect 9404 35760 9456 35766
rect 9404 35702 9456 35708
rect 9416 35630 9444 35702
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 9416 35034 9444 35566
rect 9324 35018 9444 35034
rect 9312 35012 9444 35018
rect 9364 35006 9444 35012
rect 9312 34954 9364 34960
rect 9220 33584 9272 33590
rect 9220 33526 9272 33532
rect 9232 33114 9260 33526
rect 9220 33108 9272 33114
rect 9220 33050 9272 33056
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 8668 30388 8720 30394
rect 8668 30330 8720 30336
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8588 24410 8616 24686
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8588 21622 8616 24346
rect 8680 22778 8708 30330
rect 9128 30252 9180 30258
rect 9128 30194 9180 30200
rect 9140 29578 9168 30194
rect 9128 29572 9180 29578
rect 9128 29514 9180 29520
rect 9324 28150 9352 34954
rect 9402 33960 9458 33969
rect 9402 33895 9458 33904
rect 9416 31686 9444 33895
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9312 28144 9364 28150
rect 9312 28086 9364 28092
rect 9416 27962 9444 31622
rect 9140 27934 9444 27962
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8576 21616 8628 21622
rect 8628 21576 8708 21604
rect 8576 21558 8628 21564
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8036 19922 8064 20198
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 16114 7972 17682
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8128 15162 8156 19314
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7576 14618 7604 15030
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11150 7604 11494
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3194 4660 8434
rect 8036 8090 8064 14962
rect 8588 11218 8616 17070
rect 8680 14414 8708 21576
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8772 19446 8800 20198
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8864 19292 8892 26318
rect 9140 24818 9168 27934
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9232 25362 9260 25774
rect 9416 25498 9444 25842
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9508 25378 9536 37198
rect 10048 37188 10100 37194
rect 10048 37130 10100 37136
rect 9772 37120 9824 37126
rect 9772 37062 9824 37068
rect 9784 36854 9812 37062
rect 9772 36848 9824 36854
rect 9678 36816 9734 36825
rect 9772 36790 9824 36796
rect 9864 36848 9916 36854
rect 9864 36790 9916 36796
rect 9678 36751 9680 36760
rect 9732 36751 9734 36760
rect 9680 36722 9732 36728
rect 9876 36378 9904 36790
rect 10060 36417 10088 37130
rect 10336 37126 10364 39200
rect 11060 37188 11112 37194
rect 11060 37130 11112 37136
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10598 36816 10654 36825
rect 10654 36760 10732 36768
rect 10598 36751 10600 36760
rect 10652 36740 10732 36760
rect 10600 36722 10652 36728
rect 10508 36576 10560 36582
rect 10508 36518 10560 36524
rect 10046 36408 10102 36417
rect 9864 36372 9916 36378
rect 10046 36343 10102 36352
rect 9864 36314 9916 36320
rect 9588 36168 9640 36174
rect 9588 36110 9640 36116
rect 9600 34202 9628 36110
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9692 35018 9720 35974
rect 10060 35578 10088 36343
rect 10416 36032 10468 36038
rect 10416 35974 10468 35980
rect 9968 35550 10088 35578
rect 10324 35624 10376 35630
rect 10324 35566 10376 35572
rect 9680 35012 9732 35018
rect 9680 34954 9732 34960
rect 9588 34196 9640 34202
rect 9588 34138 9640 34144
rect 9588 33312 9640 33318
rect 9588 33254 9640 33260
rect 9600 30802 9628 33254
rect 9770 32736 9826 32745
rect 9770 32671 9826 32680
rect 9784 31822 9812 32671
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9588 30796 9640 30802
rect 9588 30738 9640 30744
rect 9588 30660 9640 30666
rect 9588 30602 9640 30608
rect 9600 30394 9628 30602
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9692 25838 9720 31078
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 9784 29782 9812 30194
rect 9876 30138 9904 31758
rect 9968 31754 9996 35550
rect 10048 35488 10100 35494
rect 10140 35488 10192 35494
rect 10048 35430 10100 35436
rect 10138 35456 10140 35465
rect 10192 35456 10194 35465
rect 10060 35154 10088 35430
rect 10138 35391 10194 35400
rect 10048 35148 10100 35154
rect 10048 35090 10100 35096
rect 10048 34536 10100 34542
rect 10152 34524 10180 35391
rect 10100 34496 10180 34524
rect 10048 34478 10100 34484
rect 10140 33448 10192 33454
rect 10140 33390 10192 33396
rect 10152 32502 10180 33390
rect 10336 33114 10364 35566
rect 10428 34678 10456 35974
rect 10520 35329 10548 36518
rect 10600 36372 10652 36378
rect 10600 36314 10652 36320
rect 10612 36174 10640 36314
rect 10704 36174 10732 36740
rect 11072 36718 11100 37130
rect 11336 37120 11388 37126
rect 11336 37062 11388 37068
rect 11060 36712 11112 36718
rect 11060 36654 11112 36660
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 10692 36168 10744 36174
rect 10692 36110 10744 36116
rect 10506 35320 10562 35329
rect 10506 35255 10562 35264
rect 10508 35216 10560 35222
rect 10508 35158 10560 35164
rect 10416 34672 10468 34678
rect 10416 34614 10468 34620
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 10324 33108 10376 33114
rect 10324 33050 10376 33056
rect 10230 33008 10286 33017
rect 10230 32943 10286 32952
rect 10244 32910 10272 32943
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10428 32570 10456 33526
rect 10520 33454 10548 35158
rect 10612 34610 10640 36110
rect 10704 35698 10732 36110
rect 11060 36032 11112 36038
rect 11060 35974 11112 35980
rect 10782 35864 10838 35873
rect 10782 35799 10784 35808
rect 10836 35799 10838 35808
rect 10784 35770 10836 35776
rect 10692 35692 10744 35698
rect 10692 35634 10744 35640
rect 10600 34604 10652 34610
rect 10600 34546 10652 34552
rect 10704 33454 10732 35634
rect 10876 35148 10928 35154
rect 10876 35090 10928 35096
rect 10784 35012 10836 35018
rect 10784 34954 10836 34960
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10692 33448 10744 33454
rect 10692 33390 10744 33396
rect 10416 32564 10468 32570
rect 10416 32506 10468 32512
rect 10140 32496 10192 32502
rect 10140 32438 10192 32444
rect 10152 32230 10180 32438
rect 10232 32292 10284 32298
rect 10232 32234 10284 32240
rect 10140 32224 10192 32230
rect 10140 32166 10192 32172
rect 9968 31726 10180 31754
rect 9876 30110 10088 30138
rect 9772 29776 9824 29782
rect 9772 29718 9824 29724
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 9864 29504 9916 29510
rect 9864 29446 9916 29452
rect 9876 29238 9904 29446
rect 9864 29232 9916 29238
rect 9864 29174 9916 29180
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9324 25350 9536 25378
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9140 22574 9168 23598
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 9140 22094 9168 22510
rect 8772 19264 8892 19292
rect 8956 22066 9168 22094
rect 9220 22092 9272 22098
rect 8772 15502 8800 19264
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17270 8892 17478
rect 8852 17264 8904 17270
rect 8852 17206 8904 17212
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 13938 8892 14214
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8956 10810 8984 22066
rect 9324 22094 9352 25350
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 9876 24682 9904 25162
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9876 24274 9904 24618
rect 9864 24268 9916 24274
rect 9864 24210 9916 24216
rect 9968 24154 9996 29650
rect 10060 28490 10088 30110
rect 10048 28484 10100 28490
rect 10048 28426 10100 28432
rect 10048 26920 10100 26926
rect 10048 26862 10100 26868
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9876 24126 9996 24154
rect 9508 23186 9536 24074
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9784 23050 9812 23258
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 22710 9444 22918
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9324 22066 9444 22094
rect 9220 22034 9272 22040
rect 9036 21956 9088 21962
rect 9036 21898 9088 21904
rect 9048 17134 9076 21898
rect 9232 21486 9260 22034
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9128 20868 9180 20874
rect 9128 20810 9180 20816
rect 9140 19310 9168 20810
rect 9416 19854 9444 22066
rect 9692 21962 9720 22374
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9784 20913 9812 21422
rect 9770 20904 9826 20913
rect 9770 20839 9826 20848
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 17134 9168 19246
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9324 17610 9352 18566
rect 9416 18290 9444 19790
rect 9600 18834 9628 19790
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9784 18426 9812 19790
rect 9876 19718 9904 24126
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9968 20534 9996 23462
rect 10060 22094 10088 26862
rect 10152 24206 10180 31726
rect 10244 30870 10272 32234
rect 10600 32224 10652 32230
rect 10600 32166 10652 32172
rect 10416 31204 10468 31210
rect 10416 31146 10468 31152
rect 10232 30864 10284 30870
rect 10232 30806 10284 30812
rect 10244 30326 10272 30806
rect 10232 30320 10284 30326
rect 10232 30262 10284 30268
rect 10428 30122 10456 31146
rect 10612 30598 10640 32166
rect 10796 31754 10824 34954
rect 10888 34746 10916 35090
rect 10966 34776 11022 34785
rect 10876 34740 10928 34746
rect 10966 34711 10968 34720
rect 10876 34682 10928 34688
rect 11020 34711 11022 34720
rect 10968 34682 11020 34688
rect 10876 34604 10928 34610
rect 10876 34546 10928 34552
rect 10888 32910 10916 34546
rect 10968 34536 11020 34542
rect 10968 34478 11020 34484
rect 10980 33561 11008 34478
rect 11072 34406 11100 35974
rect 11348 35698 11376 37062
rect 11624 36854 11652 39200
rect 12268 37262 12296 39200
rect 13556 37754 13584 39200
rect 14844 39114 14872 39200
rect 14936 39114 14964 39222
rect 14844 39086 14964 39114
rect 13556 37726 13768 37754
rect 12256 37256 12308 37262
rect 12256 37198 12308 37204
rect 13636 37256 13688 37262
rect 13740 37244 13768 37726
rect 14740 37460 14792 37466
rect 14740 37402 14792 37408
rect 13820 37256 13872 37262
rect 13740 37216 13820 37244
rect 13636 37198 13688 37204
rect 13820 37198 13872 37204
rect 11612 36848 11664 36854
rect 11612 36790 11664 36796
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12164 36712 12216 36718
rect 12164 36654 12216 36660
rect 11980 36644 12032 36650
rect 11980 36586 12032 36592
rect 11428 36576 11480 36582
rect 11428 36518 11480 36524
rect 11612 36576 11664 36582
rect 11612 36518 11664 36524
rect 11336 35692 11388 35698
rect 11336 35634 11388 35640
rect 11336 35216 11388 35222
rect 11336 35158 11388 35164
rect 11060 34400 11112 34406
rect 11060 34342 11112 34348
rect 11348 33946 11376 35158
rect 11440 34134 11468 36518
rect 11520 36236 11572 36242
rect 11520 36178 11572 36184
rect 11532 36009 11560 36178
rect 11518 36000 11574 36009
rect 11518 35935 11574 35944
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11532 35222 11560 35702
rect 11520 35216 11572 35222
rect 11520 35158 11572 35164
rect 11428 34128 11480 34134
rect 11428 34070 11480 34076
rect 11348 33918 11468 33946
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 10966 33552 11022 33561
rect 10966 33487 11022 33496
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10888 32434 10916 32846
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 11164 31890 11192 33798
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 10704 31726 10824 31754
rect 11244 31748 11296 31754
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 10704 30546 10732 31726
rect 11244 31690 11296 31696
rect 11060 31408 11112 31414
rect 11060 31350 11112 31356
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10796 30666 10824 31078
rect 10784 30660 10836 30666
rect 10784 30602 10836 30608
rect 10416 30116 10468 30122
rect 10416 30058 10468 30064
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10232 27396 10284 27402
rect 10232 27338 10284 27344
rect 10244 26518 10272 27338
rect 10336 27062 10364 27814
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10232 26512 10284 26518
rect 10232 26454 10284 26460
rect 10244 24750 10272 26454
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10428 24562 10456 30058
rect 10244 24534 10456 24562
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10060 22066 10180 22094
rect 10152 21486 10180 22066
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9876 17746 9904 19654
rect 10060 18834 10088 20334
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9048 11762 9076 14350
rect 9232 14074 9260 17546
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 15026 9812 16934
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9232 12434 9260 14010
rect 9140 12406 9260 12434
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11354 9076 11494
rect 9140 11354 9168 12406
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5368 2514 5396 2790
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 6564 2446 6592 7210
rect 8220 3058 8248 7822
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8220 2650 8248 2994
rect 9048 2922 9076 10610
rect 9140 9382 9168 11086
rect 10152 10062 10180 21422
rect 10244 21010 10272 24534
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10336 21010 10364 23122
rect 10612 22098 10640 30534
rect 10704 30518 10824 30546
rect 10796 28490 10824 30518
rect 10876 30048 10928 30054
rect 10876 29990 10928 29996
rect 10888 29646 10916 29990
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 11072 29170 11100 31350
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11256 28762 11284 31690
rect 11244 28756 11296 28762
rect 11244 28698 11296 28704
rect 10784 28484 10836 28490
rect 10784 28426 10836 28432
rect 10692 26920 10744 26926
rect 10692 26862 10744 26868
rect 10704 26450 10732 26862
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 10796 24274 10824 28426
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10888 26382 10916 26726
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 10876 25764 10928 25770
rect 10876 25706 10928 25712
rect 10784 24268 10836 24274
rect 10784 24210 10836 24216
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10600 22092 10652 22098
rect 10600 22034 10652 22040
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10336 19990 10364 20946
rect 10324 19984 10376 19990
rect 10324 19926 10376 19932
rect 10428 18170 10456 21898
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10520 18358 10548 21490
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10612 18698 10640 20946
rect 10704 20466 10732 21286
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10796 18290 10824 24006
rect 10888 23610 10916 25706
rect 10980 25362 11008 25978
rect 11348 25514 11376 32710
rect 11440 30433 11468 33918
rect 11520 33108 11572 33114
rect 11520 33050 11572 33056
rect 11532 32910 11560 33050
rect 11520 32904 11572 32910
rect 11520 32846 11572 32852
rect 11426 30424 11482 30433
rect 11426 30359 11482 30368
rect 11520 30320 11572 30326
rect 11520 30262 11572 30268
rect 11532 29850 11560 30262
rect 11520 29844 11572 29850
rect 11520 29786 11572 29792
rect 11428 29640 11480 29646
rect 11428 29582 11480 29588
rect 11440 28966 11468 29582
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11072 25486 11376 25514
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 10968 23792 11020 23798
rect 10966 23760 10968 23769
rect 11020 23760 11022 23769
rect 10966 23695 11022 23704
rect 10888 23582 11008 23610
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 10888 21146 10916 22034
rect 10980 21962 11008 23582
rect 11072 22642 11100 25486
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10966 21040 11022 21049
rect 10966 20975 11022 20984
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 10888 20058 10916 20266
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10980 19446 11008 20975
rect 11072 20942 11100 22578
rect 11164 22574 11192 24686
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11164 20058 11192 22510
rect 11256 21321 11284 22918
rect 11242 21312 11298 21321
rect 11242 21247 11298 21256
rect 11440 20942 11468 28902
rect 11520 27872 11572 27878
rect 11520 27814 11572 27820
rect 11532 27402 11560 27814
rect 11520 27396 11572 27402
rect 11520 27338 11572 27344
rect 11520 27056 11572 27062
rect 11520 26998 11572 27004
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11164 19446 11192 19654
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11532 18426 11560 26998
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10428 18142 10548 18170
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10428 15434 10456 18022
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10336 13870 10364 15370
rect 10520 13938 10548 18142
rect 10796 17542 10824 18226
rect 11532 17882 11560 18362
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 11164 17338 11192 17546
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10796 13870 10824 14758
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10336 11354 10364 13806
rect 10796 13394 10824 13806
rect 11072 13394 11100 13874
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12918 10916 13194
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 11624 12434 11652 36518
rect 11992 36378 12020 36586
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 11980 36372 12032 36378
rect 11980 36314 12032 36320
rect 11900 36106 11928 36314
rect 11888 36100 11940 36106
rect 11888 36042 11940 36048
rect 12072 36032 12124 36038
rect 12072 35974 12124 35980
rect 11794 35864 11850 35873
rect 11978 35864 12034 35873
rect 11850 35822 11928 35850
rect 11794 35799 11850 35808
rect 11900 35766 11928 35822
rect 11978 35799 12034 35808
rect 11888 35760 11940 35766
rect 11888 35702 11940 35708
rect 11888 35216 11940 35222
rect 11888 35158 11940 35164
rect 11900 34678 11928 35158
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11704 34604 11756 34610
rect 11704 34546 11756 34552
rect 11716 33998 11744 34546
rect 11704 33992 11756 33998
rect 11704 33934 11756 33940
rect 11992 33658 12020 35799
rect 12084 35766 12112 35974
rect 12072 35760 12124 35766
rect 12072 35702 12124 35708
rect 12176 35018 12204 36654
rect 12256 36644 12308 36650
rect 12256 36586 12308 36592
rect 12268 35018 12296 36586
rect 12348 35828 12400 35834
rect 12348 35770 12400 35776
rect 12164 35012 12216 35018
rect 12164 34954 12216 34960
rect 12256 35012 12308 35018
rect 12256 34954 12308 34960
rect 12256 34128 12308 34134
rect 12256 34070 12308 34076
rect 12268 33998 12296 34070
rect 12164 33992 12216 33998
rect 12164 33934 12216 33940
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 12072 33856 12124 33862
rect 12072 33798 12124 33804
rect 12084 33697 12112 33798
rect 12070 33688 12126 33697
rect 11980 33652 12032 33658
rect 12070 33623 12126 33632
rect 11980 33594 12032 33600
rect 12176 33522 12204 33934
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 11704 32428 11756 32434
rect 11704 32370 11756 32376
rect 11716 32337 11744 32370
rect 11702 32328 11758 32337
rect 11702 32263 11758 32272
rect 12072 32020 12124 32026
rect 12072 31962 12124 31968
rect 12084 31736 12112 31962
rect 11900 31708 12112 31736
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11716 30938 11744 31282
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11796 30184 11848 30190
rect 11796 30126 11848 30132
rect 11808 29714 11836 30126
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11716 26042 11744 29242
rect 11900 28626 11928 31708
rect 12176 30954 12204 33458
rect 12256 33448 12308 33454
rect 12256 33390 12308 33396
rect 12268 32434 12296 33390
rect 12360 32910 12388 35770
rect 12636 35630 12664 36722
rect 13648 36718 13676 37198
rect 13636 36712 13688 36718
rect 13636 36654 13688 36660
rect 12992 36644 13044 36650
rect 12992 36586 13044 36592
rect 14372 36644 14424 36650
rect 14372 36586 14424 36592
rect 13004 36174 13032 36586
rect 13176 36576 13228 36582
rect 13176 36518 13228 36524
rect 13188 36242 13216 36518
rect 13176 36236 13228 36242
rect 13176 36178 13228 36184
rect 13820 36236 13872 36242
rect 13820 36178 13872 36184
rect 12992 36168 13044 36174
rect 12992 36110 13044 36116
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 13096 35834 13124 36110
rect 13084 35828 13136 35834
rect 13084 35770 13136 35776
rect 12716 35692 12768 35698
rect 12716 35634 12768 35640
rect 12624 35624 12676 35630
rect 12624 35566 12676 35572
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 12532 32836 12584 32842
rect 12532 32778 12584 32784
rect 12348 32768 12400 32774
rect 12348 32710 12400 32716
rect 12360 32473 12388 32710
rect 12346 32464 12402 32473
rect 12256 32428 12308 32434
rect 12346 32399 12402 32408
rect 12256 32370 12308 32376
rect 11992 30926 12204 30954
rect 11888 28620 11940 28626
rect 11888 28562 11940 28568
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11808 26790 11836 28494
rect 11888 28212 11940 28218
rect 11888 28154 11940 28160
rect 11900 27878 11928 28154
rect 11888 27872 11940 27878
rect 11888 27814 11940 27820
rect 11992 27010 12020 30926
rect 12164 30728 12216 30734
rect 12268 30716 12296 32370
rect 12544 31890 12572 32778
rect 12532 31884 12584 31890
rect 12532 31826 12584 31832
rect 12544 31754 12572 31826
rect 12544 31726 12664 31754
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12216 30688 12296 30716
rect 12164 30670 12216 30676
rect 12176 30054 12204 30670
rect 12256 30116 12308 30122
rect 12256 30058 12308 30064
rect 12164 30048 12216 30054
rect 12164 29990 12216 29996
rect 12268 29714 12296 30058
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12268 29594 12296 29650
rect 12176 29566 12296 29594
rect 12348 29572 12400 29578
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12084 27130 12112 27270
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 11992 26982 12112 27010
rect 11796 26784 11848 26790
rect 11796 26726 11848 26732
rect 11704 26036 11756 26042
rect 11704 25978 11756 25984
rect 11808 23118 11836 26726
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 22574 11836 22918
rect 11900 22710 11928 22986
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 11716 15706 11744 22442
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11808 21321 11836 21490
rect 11794 21312 11850 21321
rect 11794 21247 11850 21256
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11808 20534 11836 20946
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11900 16454 11928 19722
rect 11992 18834 12020 24074
rect 12084 22166 12112 26982
rect 12176 22982 12204 29566
rect 12348 29514 12400 29520
rect 12360 29306 12388 29514
rect 12348 29300 12400 29306
rect 12348 29242 12400 29248
rect 12256 29164 12308 29170
rect 12256 29106 12308 29112
rect 12268 28490 12296 29106
rect 12452 28626 12480 31214
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12256 28484 12308 28490
rect 12256 28426 12308 28432
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 23866 12296 24074
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12360 22506 12388 27406
rect 12348 22500 12400 22506
rect 12348 22442 12400 22448
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12256 21888 12308 21894
rect 12254 21856 12256 21865
rect 12308 21856 12310 21865
rect 12254 21791 12310 21800
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12164 21616 12216 21622
rect 12268 21593 12296 21626
rect 12164 21558 12216 21564
rect 12254 21584 12310 21593
rect 12176 20602 12204 21558
rect 12254 21519 12310 21528
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12268 21146 12296 21354
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12164 20596 12216 20602
rect 12164 20538 12216 20544
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12084 19718 12112 19858
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12084 19378 12112 19654
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12268 18698 12296 20742
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12360 18034 12388 21898
rect 12452 19242 12480 28562
rect 12544 28218 12572 28630
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12544 22710 12572 22918
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12532 22092 12584 22098
rect 12636 22094 12664 31726
rect 12728 29186 12756 35634
rect 12900 35624 12952 35630
rect 12900 35566 12952 35572
rect 13084 35624 13136 35630
rect 13084 35566 13136 35572
rect 12808 34944 12860 34950
rect 12808 34886 12860 34892
rect 12820 34678 12848 34886
rect 12808 34672 12860 34678
rect 12808 34614 12860 34620
rect 12912 33289 12940 35566
rect 13096 34542 13124 35566
rect 13188 35154 13216 36178
rect 13544 36032 13596 36038
rect 13832 36009 13860 36178
rect 13544 35974 13596 35980
rect 13818 36000 13874 36009
rect 13556 35465 13584 35974
rect 13818 35935 13874 35944
rect 14278 36000 14334 36009
rect 14278 35935 14334 35944
rect 13542 35456 13598 35465
rect 13542 35391 13598 35400
rect 13176 35148 13228 35154
rect 13176 35090 13228 35096
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 13268 35012 13320 35018
rect 13268 34954 13320 34960
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 13188 34202 13216 34954
rect 13176 34196 13228 34202
rect 13176 34138 13228 34144
rect 13084 33992 13136 33998
rect 13084 33934 13136 33940
rect 13096 33658 13124 33934
rect 13084 33652 13136 33658
rect 13084 33594 13136 33600
rect 13280 33504 13308 34954
rect 13360 34196 13412 34202
rect 13360 34138 13412 34144
rect 13188 33476 13308 33504
rect 13188 33386 13216 33476
rect 13372 33402 13400 34138
rect 13636 33856 13688 33862
rect 13636 33798 13688 33804
rect 13176 33380 13228 33386
rect 13176 33322 13228 33328
rect 13280 33374 13400 33402
rect 12898 33280 12954 33289
rect 12898 33215 12954 33224
rect 12806 32464 12862 32473
rect 12806 32399 12862 32408
rect 12820 31958 12848 32399
rect 12808 31952 12860 31958
rect 12808 31894 12860 31900
rect 12808 31748 12860 31754
rect 12808 31690 12860 31696
rect 12820 31482 12848 31690
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12820 30394 12848 30534
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12728 29158 12848 29186
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12728 27062 12756 29038
rect 12820 27470 12848 29158
rect 12912 27606 12940 33215
rect 13188 32858 13216 33322
rect 13280 33318 13308 33374
rect 13268 33312 13320 33318
rect 13268 33254 13320 33260
rect 13360 33312 13412 33318
rect 13360 33254 13412 33260
rect 13188 32830 13308 32858
rect 13372 32842 13400 33254
rect 13084 32768 13136 32774
rect 13084 32710 13136 32716
rect 13176 32768 13228 32774
rect 13176 32710 13228 32716
rect 13280 32722 13308 32830
rect 13360 32836 13412 32842
rect 13360 32778 13412 32784
rect 12990 32600 13046 32609
rect 12990 32535 13046 32544
rect 13004 32502 13032 32535
rect 13096 32502 13124 32710
rect 12992 32496 13044 32502
rect 12992 32438 13044 32444
rect 13084 32496 13136 32502
rect 13084 32438 13136 32444
rect 12992 30592 13044 30598
rect 12992 30534 13044 30540
rect 12900 27600 12952 27606
rect 12900 27542 12952 27548
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12716 26512 12768 26518
rect 12716 26454 12768 26460
rect 12728 26314 12756 26454
rect 12716 26308 12768 26314
rect 12716 26250 12768 26256
rect 12820 22642 12848 26930
rect 13004 26330 13032 30534
rect 13188 29238 13216 32710
rect 13280 32694 13492 32722
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13372 31754 13400 31826
rect 13280 31726 13400 31754
rect 13280 30802 13308 31726
rect 13464 30802 13492 32694
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 13176 29232 13228 29238
rect 13176 29174 13228 29180
rect 13084 28008 13136 28014
rect 13082 27976 13084 27985
rect 13136 27976 13138 27985
rect 13082 27911 13138 27920
rect 13176 27532 13228 27538
rect 13176 27474 13228 27480
rect 13084 27396 13136 27402
rect 13084 27338 13136 27344
rect 13096 27130 13124 27338
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 12912 26302 13032 26330
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12820 22098 12848 22442
rect 12636 22066 12756 22094
rect 12532 22034 12584 22040
rect 12544 21978 12572 22034
rect 12544 21950 12664 21978
rect 12532 21888 12584 21894
rect 12530 21856 12532 21865
rect 12584 21856 12586 21865
rect 12530 21791 12586 21800
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12544 21457 12572 21490
rect 12530 21448 12586 21457
rect 12530 21383 12586 21392
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12544 19922 12572 21286
rect 12636 21078 12664 21950
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12636 19854 12664 20742
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18222 12664 19110
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12268 18006 12388 18034
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 12084 14550 12112 17546
rect 12268 16046 12296 18006
rect 12360 17882 12480 17898
rect 12348 17876 12480 17882
rect 12400 17870 12480 17876
rect 12348 17818 12400 17824
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14006 11928 14214
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 12084 13870 12112 14486
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12268 12918 12296 15982
rect 12452 15910 12480 17870
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 11532 12406 11652 12434
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9140 8090 9168 9318
rect 11532 8090 11560 12406
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9140 6798 9168 7142
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 12176 2514 12204 12786
rect 12636 11898 12664 18158
rect 12728 15434 12756 22066
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 12820 20534 12848 22034
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12820 19310 12848 20334
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12912 18902 12940 26302
rect 13188 24682 13216 27474
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13280 24562 13308 30738
rect 13452 29572 13504 29578
rect 13452 29514 13504 29520
rect 13464 29034 13492 29514
rect 13648 29510 13676 33798
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 13372 26450 13400 27950
rect 13360 26444 13412 26450
rect 13360 26386 13412 26392
rect 13096 24534 13308 24562
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13004 21350 13032 22578
rect 13096 21536 13124 24534
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13372 23322 13400 24006
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13464 22094 13492 28970
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13556 27674 13584 28494
rect 13544 27668 13596 27674
rect 13544 27610 13596 27616
rect 13636 22432 13688 22438
rect 13636 22374 13688 22380
rect 13464 22066 13584 22094
rect 13096 21508 13308 21536
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13004 20806 13032 21286
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13188 19922 13216 20470
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13096 19786 13124 19858
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 13004 15162 13032 19722
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13096 17746 13124 19450
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13188 18698 13216 19382
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13188 15570 13216 18634
rect 13280 18222 13308 21508
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13464 20942 13492 21354
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 19514 13492 20334
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13556 19446 13584 22066
rect 13648 21622 13676 22374
rect 13636 21616 13688 21622
rect 13740 21593 13768 33458
rect 13832 33046 13860 35935
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 13912 34672 13964 34678
rect 13912 34614 13964 34620
rect 13820 33040 13872 33046
rect 13820 32982 13872 32988
rect 13924 30190 13952 34614
rect 13912 30184 13964 30190
rect 13912 30126 13964 30132
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13832 26042 13860 26182
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13636 21558 13688 21564
rect 13726 21584 13782 21593
rect 13726 21519 13782 21528
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13280 17785 13308 18158
rect 13266 17776 13322 17785
rect 13266 17711 13322 17720
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13556 15026 13584 16594
rect 13740 16250 13768 18838
rect 13924 18358 13952 19654
rect 14016 19242 14044 35022
rect 14186 34640 14242 34649
rect 14186 34575 14188 34584
rect 14240 34575 14242 34584
rect 14188 34546 14240 34552
rect 14292 34202 14320 35935
rect 14384 35086 14412 36586
rect 14464 36100 14516 36106
rect 14464 36042 14516 36048
rect 14476 35834 14504 36042
rect 14464 35828 14516 35834
rect 14464 35770 14516 35776
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14384 34678 14412 35022
rect 14660 34950 14688 35022
rect 14556 34944 14608 34950
rect 14556 34886 14608 34892
rect 14648 34944 14700 34950
rect 14648 34886 14700 34892
rect 14372 34672 14424 34678
rect 14372 34614 14424 34620
rect 14464 34468 14516 34474
rect 14464 34410 14516 34416
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14476 33930 14504 34410
rect 14568 33998 14596 34886
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 14464 33924 14516 33930
rect 14464 33866 14516 33872
rect 14648 33448 14700 33454
rect 14648 33390 14700 33396
rect 14096 33040 14148 33046
rect 14096 32982 14148 32988
rect 14108 31278 14136 32982
rect 14556 32360 14608 32366
rect 14556 32302 14608 32308
rect 14096 31272 14148 31278
rect 14096 31214 14148 31220
rect 14108 29238 14136 31214
rect 14568 31210 14596 32302
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14370 30288 14426 30297
rect 14370 30223 14372 30232
rect 14424 30223 14426 30232
rect 14372 30194 14424 30200
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 14096 29232 14148 29238
rect 14096 29174 14148 29180
rect 14096 27532 14148 27538
rect 14096 27474 14148 27480
rect 14108 26926 14136 27474
rect 14188 27056 14240 27062
rect 14188 26998 14240 27004
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 19854 14136 20742
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14108 19378 14136 19790
rect 14200 19514 14228 26998
rect 14292 25906 14320 30058
rect 14372 28144 14424 28150
rect 14372 28086 14424 28092
rect 14384 27606 14412 28086
rect 14372 27600 14424 27606
rect 14372 27542 14424 27548
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14372 25696 14424 25702
rect 14372 25638 14424 25644
rect 14384 25294 14412 25638
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14384 23730 14412 24074
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 14384 20942 14412 23462
rect 14372 20936 14424 20942
rect 14278 20904 14334 20913
rect 14372 20878 14424 20884
rect 14278 20839 14334 20848
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14004 19236 14056 19242
rect 14004 19178 14056 19184
rect 13912 18352 13964 18358
rect 13912 18294 13964 18300
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12782 13124 13126
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9722 12480 9998
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12452 6866 12480 8910
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5184 800 5212 2246
rect 6472 800 6500 2246
rect 7116 800 7144 2382
rect 8404 800 8432 2382
rect 9692 800 9720 2382
rect 10336 800 10364 2382
rect 11624 800 11652 2382
rect 12452 2310 12480 6258
rect 12544 2650 12572 11698
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 13004 3058 13032 11086
rect 13096 9586 13124 12718
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12912 800 12940 2382
rect 13004 2310 13032 2994
rect 13188 2650 13216 12174
rect 13556 11558 13584 14962
rect 13648 13938 13676 15098
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13372 2378 13400 11018
rect 14016 5642 14044 18022
rect 14108 17542 14136 18022
rect 14292 17678 14320 20839
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 19990 14412 20334
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 15094 14412 17478
rect 14476 16658 14504 30670
rect 14660 29170 14688 33390
rect 14752 31754 14780 37402
rect 15120 37244 15148 39222
rect 16118 39200 16174 39800
rect 16762 39200 16818 39800
rect 18050 39200 18106 39800
rect 18156 39222 18368 39250
rect 15200 37256 15252 37262
rect 15120 37216 15200 37244
rect 15200 37198 15252 37204
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 15934 37224 15990 37233
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 14936 36922 14964 37062
rect 14924 36916 14976 36922
rect 14924 36858 14976 36864
rect 14924 33040 14976 33046
rect 14924 32982 14976 32988
rect 14936 32570 14964 32982
rect 14924 32564 14976 32570
rect 14924 32506 14976 32512
rect 14924 32428 14976 32434
rect 15028 32416 15056 37062
rect 15304 34898 15332 37198
rect 15934 37159 15936 37168
rect 15988 37159 15990 37168
rect 15936 37130 15988 37136
rect 16132 37126 16160 39200
rect 16776 37126 16804 39200
rect 18064 39114 18092 39200
rect 18156 39114 18184 39222
rect 18064 39086 18184 39114
rect 17776 37460 17828 37466
rect 17776 37402 17828 37408
rect 16856 37256 16908 37262
rect 16856 37198 16908 37204
rect 16120 37120 16172 37126
rect 16120 37062 16172 37068
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 15660 36848 15712 36854
rect 16868 36825 16896 37198
rect 17788 36922 17816 37402
rect 17868 37392 17920 37398
rect 18144 37392 18196 37398
rect 17920 37340 18144 37346
rect 17868 37334 18196 37340
rect 17880 37318 18184 37334
rect 18236 37256 18288 37262
rect 17880 37216 18236 37244
rect 17776 36916 17828 36922
rect 17776 36858 17828 36864
rect 17880 36854 17908 37216
rect 18236 37198 18288 37204
rect 18340 37194 18368 39222
rect 19338 39200 19394 39800
rect 19982 39200 20038 39800
rect 21270 39200 21326 39800
rect 22558 39200 22614 39800
rect 23202 39200 23258 39800
rect 24490 39200 24546 39800
rect 25778 39200 25834 39800
rect 26422 39200 26478 39800
rect 27710 39200 27766 39800
rect 28998 39200 29054 39800
rect 29642 39200 29698 39800
rect 30930 39200 30986 39800
rect 32218 39200 32274 39800
rect 32862 39200 32918 39800
rect 34150 39200 34206 39800
rect 34256 39222 34468 39250
rect 18972 37392 19024 37398
rect 18972 37334 19024 37340
rect 18878 37224 18934 37233
rect 18328 37188 18380 37194
rect 18878 37159 18880 37168
rect 18328 37130 18380 37136
rect 18932 37159 18934 37168
rect 18880 37130 18932 37136
rect 18052 36916 18104 36922
rect 18052 36858 18104 36864
rect 17868 36848 17920 36854
rect 15660 36790 15712 36796
rect 16854 36816 16910 36825
rect 15384 35284 15436 35290
rect 15384 35226 15436 35232
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15212 34870 15332 34898
rect 15212 34202 15240 34870
rect 15290 34776 15346 34785
rect 15290 34711 15346 34720
rect 15304 34678 15332 34711
rect 15292 34672 15344 34678
rect 15292 34614 15344 34620
rect 15200 34196 15252 34202
rect 15200 34138 15252 34144
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 14976 32388 15056 32416
rect 14924 32370 14976 32376
rect 15108 32360 15160 32366
rect 15212 32337 15240 32506
rect 15108 32302 15160 32308
rect 15198 32328 15254 32337
rect 15016 32224 15068 32230
rect 15016 32166 15068 32172
rect 15028 31958 15056 32166
rect 15016 31952 15068 31958
rect 15016 31894 15068 31900
rect 15120 31822 15148 32302
rect 15396 32298 15424 35226
rect 15580 33862 15608 35226
rect 15568 33856 15620 33862
rect 15568 33798 15620 33804
rect 15474 33144 15530 33153
rect 15474 33079 15530 33088
rect 15198 32263 15254 32272
rect 15384 32292 15436 32298
rect 15384 32234 15436 32240
rect 15384 31884 15436 31890
rect 15384 31826 15436 31832
rect 15108 31816 15160 31822
rect 15108 31758 15160 31764
rect 14752 31726 14964 31754
rect 14832 30660 14884 30666
rect 14832 30602 14884 30608
rect 14844 29850 14872 30602
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14568 26994 14596 28018
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14568 26450 14596 26930
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14556 24676 14608 24682
rect 14556 24618 14608 24624
rect 14568 23594 14596 24618
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 14660 22094 14688 28970
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 14844 27606 14872 27950
rect 14832 27600 14884 27606
rect 14832 27542 14884 27548
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14568 22066 14688 22094
rect 14568 20534 14596 22066
rect 14752 21962 14780 25094
rect 14740 21956 14792 21962
rect 14740 21898 14792 21904
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14646 21040 14702 21049
rect 14646 20975 14702 20984
rect 14660 20942 14688 20975
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14752 20534 14780 21082
rect 14556 20528 14608 20534
rect 14556 20470 14608 20476
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 14844 20058 14872 26250
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14568 15502 14596 18226
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14936 14414 14964 31726
rect 15120 30802 15148 31758
rect 15108 30796 15160 30802
rect 15108 30738 15160 30744
rect 15108 30320 15160 30326
rect 15108 30262 15160 30268
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 15120 29646 15148 30262
rect 15108 29640 15160 29646
rect 15108 29582 15160 29588
rect 15120 28626 15148 29582
rect 15108 28620 15160 28626
rect 15108 28562 15160 28568
rect 15120 28150 15148 28562
rect 15108 28144 15160 28150
rect 15108 28086 15160 28092
rect 15304 25922 15332 30262
rect 15396 29782 15424 31826
rect 15488 30297 15516 33079
rect 15672 31754 15700 36790
rect 15752 36780 15804 36786
rect 17868 36790 17920 36796
rect 16854 36751 16910 36760
rect 15752 36722 15804 36728
rect 15764 34649 15792 36722
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 16210 36408 16266 36417
rect 16210 36343 16266 36352
rect 16224 36106 16252 36343
rect 16868 36242 16896 36654
rect 17682 36408 17738 36417
rect 17682 36343 17738 36352
rect 17960 36372 18012 36378
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 16948 36236 17000 36242
rect 16948 36178 17000 36184
rect 16212 36100 16264 36106
rect 16212 36042 16264 36048
rect 16672 36100 16724 36106
rect 16672 36042 16724 36048
rect 16684 35562 16712 36042
rect 16868 35698 16896 36178
rect 16960 36009 16988 36178
rect 16946 36000 17002 36009
rect 16946 35935 17002 35944
rect 17592 35760 17644 35766
rect 17592 35702 17644 35708
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16672 35556 16724 35562
rect 16672 35498 16724 35504
rect 16396 35488 16448 35494
rect 16396 35430 16448 35436
rect 15750 34640 15806 34649
rect 15750 34575 15806 34584
rect 15764 33862 15792 34575
rect 16304 34400 16356 34406
rect 16304 34342 16356 34348
rect 15934 33960 15990 33969
rect 15934 33895 15936 33904
rect 15988 33895 15990 33904
rect 16120 33924 16172 33930
rect 15936 33866 15988 33872
rect 16120 33866 16172 33872
rect 15752 33856 15804 33862
rect 15752 33798 15804 33804
rect 15948 33454 15976 33866
rect 16132 33590 16160 33866
rect 16120 33584 16172 33590
rect 16120 33526 16172 33532
rect 15936 33448 15988 33454
rect 15936 33390 15988 33396
rect 15752 33380 15804 33386
rect 15752 33322 15804 33328
rect 15580 31726 15700 31754
rect 15580 30802 15608 31726
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 15764 30666 15792 33322
rect 16316 33153 16344 34342
rect 16408 33454 16436 35430
rect 16868 35154 16896 35634
rect 17132 35624 17184 35630
rect 17130 35592 17132 35601
rect 17500 35624 17552 35630
rect 17184 35592 17186 35601
rect 17052 35550 17130 35578
rect 16856 35148 16908 35154
rect 16856 35090 16908 35096
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16684 33522 16712 34342
rect 16868 34066 16896 35090
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16868 33522 16896 34002
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16396 33448 16448 33454
rect 16396 33390 16448 33396
rect 16302 33144 16358 33153
rect 16302 33079 16358 33088
rect 16948 32904 17000 32910
rect 16946 32872 16948 32881
rect 17000 32872 17002 32881
rect 16946 32807 17002 32816
rect 15844 32496 15896 32502
rect 15844 32438 15896 32444
rect 15856 31754 15884 32438
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16868 32230 16896 32370
rect 16764 32224 16816 32230
rect 16764 32166 16816 32172
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16672 31952 16724 31958
rect 16672 31894 16724 31900
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 16120 31204 16172 31210
rect 16120 31146 16172 31152
rect 15752 30660 15804 30666
rect 15752 30602 15804 30608
rect 16132 30326 16160 31146
rect 16580 30388 16632 30394
rect 16580 30330 16632 30336
rect 16120 30320 16172 30326
rect 15474 30288 15530 30297
rect 16120 30262 16172 30268
rect 15474 30223 15530 30232
rect 16028 30116 16080 30122
rect 16028 30058 16080 30064
rect 15384 29776 15436 29782
rect 15384 29718 15436 29724
rect 16040 29714 16068 30058
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16132 29714 16160 29990
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15672 29578 15700 29650
rect 15660 29572 15712 29578
rect 15488 29532 15660 29560
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15212 25894 15332 25922
rect 15212 22778 15240 25894
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15304 23633 15332 25774
rect 15290 23624 15346 23633
rect 15290 23559 15346 23568
rect 15304 23050 15332 23559
rect 15396 23322 15424 27542
rect 15488 26330 15516 29532
rect 15660 29514 15712 29520
rect 16120 29028 16172 29034
rect 16120 28970 16172 28976
rect 16132 28694 16160 28970
rect 16120 28688 16172 28694
rect 16120 28630 16172 28636
rect 16316 28218 16344 29990
rect 16592 29238 16620 30330
rect 16684 29594 16712 31894
rect 16776 31822 16804 32166
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16776 30802 16804 31758
rect 16764 30796 16816 30802
rect 16764 30738 16816 30744
rect 16856 30728 16908 30734
rect 16856 30670 16908 30676
rect 16764 30116 16816 30122
rect 16764 30058 16816 30064
rect 16776 29782 16804 30058
rect 16764 29776 16816 29782
rect 16764 29718 16816 29724
rect 16684 29566 16804 29594
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16684 29306 16712 29446
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 16396 29096 16448 29102
rect 16396 29038 16448 29044
rect 16304 28212 16356 28218
rect 16304 28154 16356 28160
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15580 27470 15608 27950
rect 15568 27464 15620 27470
rect 15568 27406 15620 27412
rect 16316 26926 16344 28154
rect 16304 26920 16356 26926
rect 16304 26862 16356 26868
rect 15844 26852 15896 26858
rect 15844 26794 15896 26800
rect 15856 26602 15884 26794
rect 16408 26790 16436 29038
rect 16776 28966 16804 29566
rect 16868 29306 16896 30670
rect 16948 29572 17000 29578
rect 16948 29514 17000 29520
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16868 29170 16896 29242
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 16764 28960 16816 28966
rect 16764 28902 16816 28908
rect 16500 28490 16528 28902
rect 16488 28484 16540 28490
rect 16488 28426 16540 28432
rect 16500 28218 16528 28426
rect 16488 28212 16540 28218
rect 16488 28154 16540 28160
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 16396 26784 16448 26790
rect 16396 26726 16448 26732
rect 15580 26574 15884 26602
rect 15580 26518 15608 26574
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15948 26450 15976 26726
rect 15936 26444 15988 26450
rect 15936 26386 15988 26392
rect 15488 26302 15700 26330
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15580 24206 15608 24686
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15384 23316 15436 23322
rect 15384 23258 15436 23264
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15212 18766 15240 21082
rect 15382 21040 15438 21049
rect 15382 20975 15384 20984
rect 15436 20975 15438 20984
rect 15384 20946 15436 20952
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15028 15094 15056 16186
rect 15120 15978 15148 17546
rect 15108 15972 15160 15978
rect 15108 15914 15160 15920
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15212 14414 15240 14894
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 13530 14504 13806
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 12714 14872 13262
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14936 11150 14964 14350
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 14292 2650 14320 10542
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14660 9042 14688 10406
rect 14936 9926 14964 10678
rect 15212 10674 15240 14350
rect 15304 14346 15332 19654
rect 15396 19446 15424 19654
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15580 18970 15608 22170
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15672 17678 15700 26302
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15764 24206 15792 25094
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 24410 15884 24550
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15764 23866 15792 24142
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15764 23186 15792 23802
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15844 21480 15896 21486
rect 15842 21448 15844 21457
rect 15896 21448 15898 21457
rect 15842 21383 15898 21392
rect 15948 19854 15976 25978
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15856 12850 15884 13738
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 11150 15884 12786
rect 16040 11830 16068 24346
rect 16316 24138 16344 24890
rect 16304 24132 16356 24138
rect 16304 24074 16356 24080
rect 16212 23792 16264 23798
rect 16212 23734 16264 23740
rect 16224 21622 16252 23734
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16408 20602 16436 26726
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 25106 16804 26182
rect 16868 25294 16896 29106
rect 16960 29102 16988 29514
rect 16948 29096 17000 29102
rect 16948 29038 17000 29044
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16948 25220 17000 25226
rect 16948 25162 17000 25168
rect 16856 25152 16908 25158
rect 16776 25100 16856 25106
rect 16776 25094 16908 25100
rect 16776 25078 16896 25094
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16684 23526 16712 24006
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16776 23322 16804 23598
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16776 22094 16804 23258
rect 16592 22066 16804 22094
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16316 19446 16344 19858
rect 16592 19854 16620 22066
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16776 21690 16804 21898
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16684 17610 16712 20266
rect 16776 20058 16804 20470
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16776 19378 16804 19722
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16868 16674 16896 25078
rect 16960 21962 16988 25162
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16960 19786 16988 21490
rect 17052 21146 17080 35550
rect 17500 35566 17552 35572
rect 17130 35527 17186 35536
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17132 33856 17184 33862
rect 17130 33824 17132 33833
rect 17184 33824 17186 33833
rect 17130 33759 17186 33768
rect 17144 33658 17172 33759
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 17236 32502 17264 35430
rect 17406 35320 17462 35329
rect 17406 35255 17462 35264
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17224 32496 17276 32502
rect 17224 32438 17276 32444
rect 17236 28014 17264 32438
rect 17224 28008 17276 28014
rect 17224 27950 17276 27956
rect 17328 26858 17356 35022
rect 17420 33862 17448 35255
rect 17512 35086 17540 35566
rect 17500 35080 17552 35086
rect 17500 35022 17552 35028
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17500 32972 17552 32978
rect 17500 32914 17552 32920
rect 17512 32881 17540 32914
rect 17498 32872 17554 32881
rect 17408 32836 17460 32842
rect 17498 32807 17554 32816
rect 17408 32778 17460 32784
rect 17420 31822 17448 32778
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17420 29646 17448 30534
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17500 29028 17552 29034
rect 17500 28970 17552 28976
rect 17512 28150 17540 28970
rect 17500 28144 17552 28150
rect 17500 28086 17552 28092
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17316 26852 17368 26858
rect 17316 26794 17368 26800
rect 17420 26450 17448 27270
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17512 23662 17540 24006
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 17144 21350 17172 21898
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17222 21312 17278 21321
rect 17222 21247 17278 21256
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17236 20874 17264 21247
rect 17040 20868 17092 20874
rect 17040 20810 17092 20816
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16960 18902 16988 19722
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16776 16646 16896 16674
rect 16776 15502 16804 16646
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 15026 16344 15302
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9178 14964 9862
rect 15764 9722 15792 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15856 9654 15884 11086
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10674 15976 10950
rect 16040 10810 16068 11766
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16132 10266 16160 10406
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15948 9450 15976 9998
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 16684 2514 16712 15030
rect 16776 11762 16804 15438
rect 16960 15094 16988 18702
rect 17052 18630 17080 20810
rect 17420 20058 17448 22986
rect 17604 22094 17632 35702
rect 17696 33998 17724 36343
rect 17960 36314 18012 36320
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 17776 36100 17828 36106
rect 17776 36042 17828 36048
rect 17788 35601 17816 36042
rect 17774 35592 17830 35601
rect 17774 35527 17830 35536
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17776 33448 17828 33454
rect 17774 33416 17776 33425
rect 17828 33416 17830 33425
rect 17774 33351 17830 33360
rect 17880 31890 17908 36110
rect 17972 35193 18000 36314
rect 18064 35748 18092 36858
rect 18420 36848 18472 36854
rect 18420 36790 18472 36796
rect 18432 35873 18460 36790
rect 18418 35864 18474 35873
rect 18418 35799 18474 35808
rect 18420 35760 18472 35766
rect 18064 35720 18420 35748
rect 17958 35184 18014 35193
rect 17958 35119 18014 35128
rect 18064 32609 18092 35720
rect 18420 35702 18472 35708
rect 18788 35012 18840 35018
rect 18788 34954 18840 34960
rect 18800 34678 18828 34954
rect 18788 34672 18840 34678
rect 18788 34614 18840 34620
rect 18236 34468 18288 34474
rect 18236 34410 18288 34416
rect 18248 34202 18276 34410
rect 18236 34196 18288 34202
rect 18236 34138 18288 34144
rect 18604 33992 18656 33998
rect 18604 33934 18656 33940
rect 18616 33658 18644 33934
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 18418 33144 18474 33153
rect 18418 33079 18474 33088
rect 18050 32600 18106 32609
rect 18050 32535 18106 32544
rect 18432 32502 18460 33079
rect 18420 32496 18472 32502
rect 18420 32438 18472 32444
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 17868 31884 17920 31890
rect 17868 31826 17920 31832
rect 17868 30592 17920 30598
rect 17868 30534 17920 30540
rect 17776 29096 17828 29102
rect 17776 29038 17828 29044
rect 17788 28626 17816 29038
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 28014 17816 28562
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17788 27538 17816 27950
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17880 26330 17908 30534
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 17960 28960 18012 28966
rect 17960 28902 18012 28908
rect 17972 26994 18000 28902
rect 18156 28558 18184 29038
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18156 26994 18184 28494
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 17788 26302 17908 26330
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17696 23050 17724 24074
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17512 22066 17632 22094
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17512 19514 17540 22066
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17604 19378 17632 20470
rect 17696 20466 17724 21490
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17696 19854 17724 20402
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17696 19378 17724 19790
rect 17788 19514 17816 26302
rect 18064 24614 18092 26862
rect 18144 25220 18196 25226
rect 18144 25162 18196 25168
rect 18156 24818 18184 25162
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18052 24608 18104 24614
rect 18052 24550 18104 24556
rect 18156 23866 18184 24754
rect 18248 24290 18276 32370
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18524 31890 18552 32166
rect 18512 31884 18564 31890
rect 18512 31826 18564 31832
rect 18524 31346 18552 31826
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18524 30802 18552 31282
rect 18512 30796 18564 30802
rect 18512 30738 18564 30744
rect 18524 30258 18552 30738
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18616 30190 18644 32166
rect 18800 31754 18828 34614
rect 18708 31726 18828 31754
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18328 30116 18380 30122
rect 18328 30058 18380 30064
rect 18340 24886 18368 30058
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 18432 26926 18460 27950
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18328 24880 18380 24886
rect 18328 24822 18380 24828
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18432 24410 18460 24686
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18248 24262 18460 24290
rect 18328 24132 18380 24138
rect 18328 24074 18380 24080
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18156 23662 18184 23802
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 18156 23474 18184 23598
rect 17880 23446 18184 23474
rect 17880 22710 17908 23446
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18064 22094 18092 22510
rect 18064 22066 18184 22094
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17696 18766 17724 19314
rect 17880 18902 17908 20742
rect 18064 20466 18092 20878
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17052 15162 17080 16118
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17512 15434 17540 15914
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16868 10538 16896 14214
rect 16960 13394 16988 14418
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16960 12442 16988 13330
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17052 11898 17080 13194
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 17052 9654 17080 9862
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13556 800 13584 2382
rect 14844 800 14872 2382
rect 16132 800 16160 2382
rect 16776 800 16804 2994
rect 17144 2514 17172 14282
rect 17236 13394 17264 15370
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17604 14346 17632 14962
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17788 13870 17816 15982
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 17880 14006 17908 14486
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 18156 13258 18184 22066
rect 18248 20602 18276 23666
rect 18340 22574 18368 24074
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18432 22234 18460 24262
rect 18420 22228 18472 22234
rect 18420 22170 18472 22176
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18524 18970 18552 28426
rect 18708 24954 18736 31726
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18708 23866 18736 24278
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18616 23633 18644 23802
rect 18602 23624 18658 23633
rect 18602 23559 18658 23568
rect 18602 23488 18658 23497
rect 18602 23423 18658 23432
rect 18616 19156 18644 23423
rect 18696 23044 18748 23050
rect 18696 22986 18748 22992
rect 18708 22234 18736 22986
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18694 21584 18750 21593
rect 18694 21519 18750 21528
rect 18708 20942 18736 21519
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18800 20262 18828 26726
rect 18892 20602 18920 26998
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18616 19128 18736 19156
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 16182 18552 17478
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18432 12782 18460 13806
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 17420 8634 17448 12718
rect 18616 12374 18644 13398
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18616 11830 18644 12310
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17788 10062 17816 10474
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17880 9518 17908 10202
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 18156 2650 18184 11086
rect 18708 5370 18736 19128
rect 18984 16250 19012 37334
rect 19352 37126 19380 39200
rect 19996 37126 20024 39200
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19984 37120 20036 37126
rect 19984 37062 20036 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 20260 36576 20312 36582
rect 20260 36518 20312 36524
rect 19444 36174 19472 36518
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19708 35760 19760 35766
rect 19708 35702 19760 35708
rect 20076 35760 20128 35766
rect 20076 35702 20128 35708
rect 19720 35630 19748 35702
rect 19340 35624 19392 35630
rect 19340 35566 19392 35572
rect 19616 35624 19668 35630
rect 19616 35566 19668 35572
rect 19708 35624 19760 35630
rect 19708 35566 19760 35572
rect 19352 35154 19380 35566
rect 19628 35290 19656 35566
rect 19616 35284 19668 35290
rect 19616 35226 19668 35232
rect 20088 35222 20116 35702
rect 20076 35216 20128 35222
rect 20076 35158 20128 35164
rect 19340 35148 19392 35154
rect 19340 35090 19392 35096
rect 19352 34762 19380 35090
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19352 34746 19472 34762
rect 19352 34740 19484 34746
rect 19352 34734 19432 34740
rect 19352 34066 19380 34734
rect 19432 34682 19484 34688
rect 19524 34740 19576 34746
rect 19524 34682 19576 34688
rect 19536 34626 19564 34682
rect 19444 34598 19564 34626
rect 19340 34060 19392 34066
rect 19340 34002 19392 34008
rect 19444 33946 19472 34598
rect 19996 34542 20024 34954
rect 19984 34536 20036 34542
rect 19984 34478 20036 34484
rect 19984 34196 20036 34202
rect 19984 34138 20036 34144
rect 19260 33918 19472 33946
rect 19628 33930 19932 33946
rect 19616 33924 19932 33930
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 19076 30190 19104 33594
rect 19260 32745 19288 33918
rect 19668 33918 19932 33924
rect 19616 33866 19668 33872
rect 19904 33862 19932 33918
rect 19892 33856 19944 33862
rect 19892 33798 19944 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19430 33688 19486 33697
rect 19574 33691 19882 33700
rect 19430 33623 19486 33632
rect 19444 33153 19472 33623
rect 19996 33590 20024 34138
rect 19984 33584 20036 33590
rect 19984 33526 20036 33532
rect 19430 33144 19486 33153
rect 19430 33079 19486 33088
rect 20168 33040 20220 33046
rect 20168 32982 20220 32988
rect 19246 32736 19302 32745
rect 19246 32671 19302 32680
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19260 31890 19288 32302
rect 19248 31884 19300 31890
rect 19248 31826 19300 31832
rect 20076 31884 20128 31890
rect 20076 31826 20128 31832
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 19156 30048 19208 30054
rect 19156 29990 19208 29996
rect 19168 28966 19196 29990
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 19260 27946 19288 31214
rect 20088 30682 20116 31826
rect 20180 31754 20208 32982
rect 20272 32978 20300 36518
rect 20548 36242 20576 37198
rect 21284 37126 21312 39200
rect 22572 37262 22600 39200
rect 22744 37324 22796 37330
rect 22744 37266 22796 37272
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 21272 37120 21324 37126
rect 21272 37062 21324 37068
rect 22560 36712 22612 36718
rect 22560 36654 22612 36660
rect 20628 36304 20680 36310
rect 20680 36252 20852 36258
rect 20628 36246 20852 36252
rect 20536 36236 20588 36242
rect 20640 36230 20852 36246
rect 22572 36242 22600 36654
rect 20536 36178 20588 36184
rect 20352 35080 20404 35086
rect 20350 35048 20352 35057
rect 20404 35048 20406 35057
rect 20824 35018 20852 36230
rect 22284 36236 22336 36242
rect 22284 36178 22336 36184
rect 22560 36236 22612 36242
rect 22560 36178 22612 36184
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 20996 36100 21048 36106
rect 20996 36042 21048 36048
rect 20902 35728 20958 35737
rect 20902 35663 20958 35672
rect 20350 34983 20406 34992
rect 20720 35012 20772 35018
rect 20720 34954 20772 34960
rect 20812 35012 20864 35018
rect 20812 34954 20864 34960
rect 20732 34746 20760 34954
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20916 34678 20944 35663
rect 20904 34672 20956 34678
rect 20904 34614 20956 34620
rect 20902 33416 20958 33425
rect 20902 33351 20958 33360
rect 20916 33318 20944 33351
rect 20812 33312 20864 33318
rect 20812 33254 20864 33260
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 20824 32978 20852 33254
rect 20260 32972 20312 32978
rect 20260 32914 20312 32920
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 21008 31754 21036 36042
rect 22112 36009 22140 36110
rect 22098 36000 22154 36009
rect 22098 35935 22154 35944
rect 22296 35698 22324 36178
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 21824 35284 21876 35290
rect 21824 35226 21876 35232
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 21178 33960 21234 33969
rect 21178 33895 21180 33904
rect 21232 33895 21234 33904
rect 21180 33866 21232 33872
rect 21732 33448 21784 33454
rect 21732 33390 21784 33396
rect 21546 33144 21602 33153
rect 21546 33079 21602 33088
rect 21560 32842 21588 33079
rect 21548 32836 21600 32842
rect 21548 32778 21600 32784
rect 21456 32564 21508 32570
rect 21456 32506 21508 32512
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 21100 32026 21128 32370
rect 21468 32230 21496 32506
rect 21744 32366 21772 33390
rect 21836 33266 21864 35226
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 22112 34066 22140 34886
rect 22204 34746 22232 35226
rect 22296 35154 22324 35634
rect 22284 35148 22336 35154
rect 22284 35090 22336 35096
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22296 34610 22324 35090
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22020 33454 22048 33934
rect 22100 33924 22152 33930
rect 22100 33866 22152 33872
rect 22468 33924 22520 33930
rect 22468 33866 22520 33872
rect 22112 33658 22140 33866
rect 22100 33652 22152 33658
rect 22100 33594 22152 33600
rect 22008 33448 22060 33454
rect 22008 33390 22060 33396
rect 21836 33238 21956 33266
rect 21928 33130 21956 33238
rect 21928 33102 22140 33130
rect 22112 33046 22140 33102
rect 22100 33040 22152 33046
rect 22100 32982 22152 32988
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 22008 32360 22060 32366
rect 22008 32302 22060 32308
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21640 31884 21692 31890
rect 21640 31826 21692 31832
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 20916 31726 21036 31754
rect 20536 31408 20588 31414
rect 20536 31350 20588 31356
rect 20168 31136 20220 31142
rect 20168 31078 20220 31084
rect 19996 30666 20116 30682
rect 19984 30660 20116 30666
rect 20036 30654 20116 30660
rect 19984 30602 20036 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19352 28422 19380 29786
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19064 25968 19116 25974
rect 19064 25910 19116 25916
rect 19076 19514 19104 25910
rect 19260 25702 19288 27882
rect 19444 25922 19472 28426
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19444 25894 19564 25922
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19444 24750 19472 25774
rect 19536 25770 19564 25894
rect 19524 25764 19576 25770
rect 19524 25706 19576 25712
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19444 24274 19472 24686
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19168 19922 19196 21354
rect 19260 20942 19288 21966
rect 19352 21146 19380 24006
rect 19444 23186 19472 24210
rect 19536 24070 19564 24754
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 19444 21146 19472 22646
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21486 20024 30602
rect 20076 28960 20128 28966
rect 20076 28902 20128 28908
rect 20088 28490 20116 28902
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 20088 24682 20116 28426
rect 20180 28014 20208 31078
rect 20548 28234 20576 31350
rect 20916 30598 20944 31726
rect 20904 30592 20956 30598
rect 20904 30534 20956 30540
rect 20628 29640 20680 29646
rect 20680 29588 20760 29594
rect 20628 29582 20760 29588
rect 20640 29566 20760 29582
rect 20732 29102 20760 29566
rect 20720 29096 20772 29102
rect 20720 29038 20772 29044
rect 20732 28626 20760 29038
rect 20720 28620 20772 28626
rect 21100 28608 21128 31758
rect 21456 30660 21508 30666
rect 21456 30602 21508 30608
rect 21272 30592 21324 30598
rect 21272 30534 21324 30540
rect 21180 29572 21232 29578
rect 21180 29514 21232 29520
rect 20720 28562 20772 28568
rect 20916 28580 21128 28608
rect 20548 28206 20668 28234
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 20180 26042 20208 27950
rect 20548 27130 20576 28086
rect 20536 27124 20588 27130
rect 20536 27066 20588 27072
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20168 26036 20220 26042
rect 20168 25978 20220 25984
rect 20260 25424 20312 25430
rect 20260 25366 20312 25372
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20180 23662 20208 24550
rect 20272 23662 20300 25366
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 20088 22506 20116 22986
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19260 17338 19288 18362
rect 19444 18290 19472 19314
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19628 17678 19656 18022
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19260 16794 19288 17138
rect 19996 17134 20024 18770
rect 20088 17882 20116 22170
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20088 17270 20116 17478
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15162 20024 17070
rect 20180 16658 20208 23598
rect 20272 22710 20300 23598
rect 20260 22704 20312 22710
rect 20260 22646 20312 22652
rect 20272 22234 20300 22646
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20272 19514 20300 19654
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 20180 15026 20208 16390
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 12918 19012 13670
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18800 11286 18828 11630
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 19444 2650 19472 14418
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 19996 13394 20024 13806
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19904 12442 19932 12786
rect 20180 12714 20208 13806
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 19892 12436 19944 12442
rect 20364 12434 20392 26250
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20456 21010 20484 21966
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 20456 17338 20484 19926
rect 20548 19378 20576 26726
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20640 17746 20668 28206
rect 20732 28082 20760 28562
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20732 26450 20760 28018
rect 20824 27946 20852 28358
rect 20812 27940 20864 27946
rect 20812 27882 20864 27888
rect 20720 26444 20772 26450
rect 20720 26386 20772 26392
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20732 22098 20760 23734
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20824 20330 20852 24142
rect 20812 20324 20864 20330
rect 20812 20266 20864 20272
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20628 15496 20680 15502
rect 20548 15444 20628 15450
rect 20548 15438 20680 15444
rect 20548 15422 20668 15438
rect 20548 15366 20576 15422
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20732 14482 20760 19382
rect 20824 19378 20852 19722
rect 20916 19514 20944 28580
rect 21192 25820 21220 29514
rect 21100 25792 21220 25820
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 23526 21036 25638
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21008 20534 21036 22714
rect 21100 21078 21128 25792
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 21192 21298 21220 25094
rect 21284 21894 21312 30534
rect 21364 28144 21416 28150
rect 21364 28086 21416 28092
rect 21376 25158 21404 28086
rect 21468 26858 21496 30602
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21560 27130 21588 27270
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21456 26852 21508 26858
rect 21456 26794 21508 26800
rect 21454 26344 21510 26353
rect 21454 26279 21510 26288
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 21376 22778 21404 22986
rect 21468 22982 21496 26279
rect 21560 24857 21588 27066
rect 21652 25498 21680 31826
rect 22020 31822 22048 32302
rect 22008 31816 22060 31822
rect 21836 31764 22008 31770
rect 21836 31758 22060 31764
rect 21836 31742 22048 31758
rect 21836 30802 21864 31742
rect 22480 31686 22508 33866
rect 22652 32292 22704 32298
rect 22652 32234 22704 32240
rect 22664 31890 22692 32234
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 21824 30796 21876 30802
rect 21824 30738 21876 30744
rect 21916 30592 21968 30598
rect 21916 30534 21968 30540
rect 21640 25492 21692 25498
rect 21640 25434 21692 25440
rect 21546 24848 21602 24857
rect 21546 24783 21602 24792
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21272 21888 21324 21894
rect 21272 21830 21324 21836
rect 21192 21270 21496 21298
rect 21178 21176 21234 21185
rect 21178 21111 21180 21120
rect 21232 21111 21234 21120
rect 21180 21082 21232 21088
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 21270 21040 21326 21049
rect 21270 20975 21326 20984
rect 21284 20874 21312 20975
rect 21364 20936 21416 20942
rect 21362 20904 21364 20913
rect 21416 20904 21418 20913
rect 21272 20868 21324 20874
rect 21192 20828 21272 20856
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 21008 19922 21036 20470
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20904 18896 20956 18902
rect 20904 18838 20956 18844
rect 20812 14612 20864 14618
rect 20916 14600 20944 18838
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21008 16046 21036 16934
rect 21192 16590 21220 20828
rect 21362 20839 21418 20848
rect 21272 20810 21324 20816
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 21270 19136 21326 19145
rect 21270 19071 21326 19080
rect 21284 18834 21312 19071
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21376 17814 21404 19926
rect 21468 18086 21496 21270
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21560 18834 21588 20742
rect 21652 19378 21680 25434
rect 21824 23044 21876 23050
rect 21824 22986 21876 22992
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21376 17270 21404 17750
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21180 16584 21232 16590
rect 21100 16532 21180 16538
rect 21100 16526 21232 16532
rect 21100 16510 21220 16526
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20864 14572 20944 14600
rect 20812 14554 20864 14560
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 19892 12378 19944 12384
rect 20272 12406 20392 12434
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20088 11830 20116 12038
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 20088 9586 20116 11630
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20272 2650 20300 12406
rect 20916 11830 20944 14572
rect 21100 13530 21128 16510
rect 21272 15972 21324 15978
rect 21272 15914 21324 15920
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21192 14006 21220 15846
rect 21284 14550 21312 15914
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 21192 13734 21220 13942
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21468 11898 21496 17002
rect 21560 16590 21588 18770
rect 21652 18222 21680 19314
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21560 14482 21588 14894
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21652 14346 21680 15302
rect 21836 14498 21864 22986
rect 21928 18358 21956 30534
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22020 26994 22048 29106
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22020 22642 22048 26930
rect 22284 25220 22336 25226
rect 22284 25162 22336 25168
rect 22296 24682 22324 25162
rect 22284 24676 22336 24682
rect 22284 24618 22336 24624
rect 22296 23730 22324 24618
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22296 23186 22324 23666
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22296 22642 22324 23122
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22020 21010 22048 22578
rect 22388 22506 22416 22714
rect 22376 22500 22428 22506
rect 22376 22442 22428 22448
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22204 21554 22232 21898
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22020 20466 22048 20946
rect 22204 20942 22232 21490
rect 22376 21344 22428 21350
rect 22376 21286 22428 21292
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22112 18698 22140 19110
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 21916 18352 21968 18358
rect 21916 18294 21968 18300
rect 22388 18290 22416 21286
rect 22480 18834 22508 27338
rect 22560 26308 22612 26314
rect 22560 26250 22612 26256
rect 22572 20058 22600 26250
rect 22664 21486 22692 31826
rect 22756 26586 22784 37266
rect 23216 37126 23244 39200
rect 24504 37262 24532 39200
rect 25792 37330 25820 39200
rect 25780 37324 25832 37330
rect 25780 37266 25832 37272
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 24492 37256 24544 37262
rect 24492 37198 24544 37204
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 23492 36689 23520 37198
rect 24676 36848 24728 36854
rect 24676 36790 24728 36796
rect 25504 36848 25556 36854
rect 25504 36790 25556 36796
rect 23478 36680 23534 36689
rect 23478 36615 23534 36624
rect 23940 36644 23992 36650
rect 23940 36586 23992 36592
rect 24584 36644 24636 36650
rect 24584 36586 24636 36592
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23112 36100 23164 36106
rect 23112 36042 23164 36048
rect 22928 35080 22980 35086
rect 22926 35048 22928 35057
rect 22980 35048 22982 35057
rect 23124 35018 23152 36042
rect 23296 35760 23348 35766
rect 23296 35702 23348 35708
rect 22926 34983 22982 34992
rect 23112 35012 23164 35018
rect 23112 34954 23164 34960
rect 22836 34060 22888 34066
rect 22836 34002 22888 34008
rect 22744 26580 22796 26586
rect 22744 26522 22796 26528
rect 22848 26450 22876 34002
rect 23124 32434 23152 34954
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23124 30258 23152 32370
rect 23308 31754 23336 35702
rect 23492 35154 23520 36314
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23480 35148 23532 35154
rect 23480 35090 23532 35096
rect 23584 34406 23612 35566
rect 23952 35494 23980 36586
rect 24596 36310 24624 36586
rect 24584 36304 24636 36310
rect 24584 36246 24636 36252
rect 24584 36100 24636 36106
rect 24584 36042 24636 36048
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23308 31726 23428 31754
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 23020 29708 23072 29714
rect 23020 29650 23072 29656
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22848 26330 22876 26386
rect 22756 26302 22876 26330
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22664 19378 22692 20878
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22468 17264 22520 17270
rect 22468 17206 22520 17212
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 21836 14482 21956 14498
rect 21824 14476 21956 14482
rect 21876 14470 21956 14476
rect 21824 14418 21876 14424
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21836 13938 21864 14282
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21928 13802 21956 14470
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 22020 13569 22048 17138
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22006 13560 22062 13569
rect 22006 13495 22062 13504
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 21008 9654 21036 11222
rect 21284 11218 21312 11494
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 21468 10062 21496 11834
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 8974 20392 9318
rect 20548 9178 20576 9454
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 21008 7886 21036 9590
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21652 3126 21680 13126
rect 22020 12306 22048 13495
rect 22112 13326 22140 16186
rect 22204 14006 22232 16458
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22296 15502 22324 15982
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22388 15348 22416 16050
rect 22480 15502 22508 17206
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22388 15320 22508 15348
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22388 12714 22416 14282
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22284 12164 22336 12170
rect 22284 12106 22336 12112
rect 22296 11354 22324 12106
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22388 11218 22416 12650
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21640 3120 21692 3126
rect 21640 3062 21692 3068
rect 22112 2650 22140 11086
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22192 9920 22244 9926
rect 22296 9897 22324 10610
rect 22480 10198 22508 15320
rect 22572 11082 22600 17614
rect 22664 16538 22692 19314
rect 22756 16658 22784 26302
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22848 22094 22876 25434
rect 22940 24886 22968 25774
rect 22928 24880 22980 24886
rect 22928 24822 22980 24828
rect 22940 24682 22968 24822
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 23032 22098 23060 29650
rect 23124 29306 23152 30194
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23296 28212 23348 28218
rect 23296 28154 23348 28160
rect 23308 27538 23336 28154
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23216 25838 23244 27474
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 22848 22066 22968 22094
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22848 20602 22876 21422
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 22848 18698 22876 19178
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22664 16510 22784 16538
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 15502 22692 16390
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22756 14618 22784 16510
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 22848 14346 22876 18634
rect 22940 18034 22968 22066
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 23032 20330 23060 22034
rect 23216 21350 23244 25774
rect 23400 22438 23428 31726
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23860 30802 23888 31622
rect 23952 31482 23980 35430
rect 24596 34474 24624 36042
rect 24584 34468 24636 34474
rect 24584 34410 24636 34416
rect 24032 34400 24084 34406
rect 24032 34342 24084 34348
rect 24044 31958 24072 34342
rect 24400 33924 24452 33930
rect 24400 33866 24452 33872
rect 24216 33856 24268 33862
rect 24216 33798 24268 33804
rect 24228 33454 24256 33798
rect 24216 33448 24268 33454
rect 24216 33390 24268 33396
rect 24032 31952 24084 31958
rect 24032 31894 24084 31900
rect 23940 31476 23992 31482
rect 23940 31418 23992 31424
rect 23848 30796 23900 30802
rect 23848 30738 23900 30744
rect 23940 29572 23992 29578
rect 23940 29514 23992 29520
rect 23848 24948 23900 24954
rect 23848 24890 23900 24896
rect 23860 23497 23888 24890
rect 23952 23798 23980 29514
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23846 23488 23902 23497
rect 23846 23423 23902 23432
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 23308 20942 23336 21966
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23308 20398 23336 20878
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23204 20392 23256 20398
rect 23204 20334 23256 20340
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 23216 20058 23244 20334
rect 23400 20262 23428 20538
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23032 19310 23060 19858
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23400 19334 23428 19722
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23308 19306 23428 19334
rect 23308 18068 23336 19306
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23400 18222 23428 18838
rect 23492 18426 23520 19722
rect 23584 18970 23612 20470
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23308 18040 23428 18068
rect 22940 18006 23244 18034
rect 23018 17912 23074 17921
rect 23018 17847 23074 17856
rect 23032 17678 23060 17847
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22940 17270 22968 17478
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 23216 16590 23244 18006
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23216 15450 23244 16526
rect 23032 15422 23244 15450
rect 23294 15464 23350 15473
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 14006 22968 14214
rect 23032 14074 23060 15422
rect 23294 15399 23296 15408
rect 23348 15399 23350 15408
rect 23296 15370 23348 15376
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23124 15162 23152 15302
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23124 14482 23152 15098
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22756 12918 22784 13126
rect 22744 12912 22796 12918
rect 22744 12854 22796 12860
rect 23124 12850 23152 14214
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 23216 12170 23244 15302
rect 23400 15162 23428 18040
rect 23676 16726 23704 18566
rect 23664 16720 23716 16726
rect 23664 16662 23716 16668
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23308 13870 23336 14486
rect 23492 13938 23520 16594
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23584 15026 23612 16390
rect 23662 15192 23718 15201
rect 23662 15127 23718 15136
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23676 14414 23704 15127
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23204 12164 23256 12170
rect 23204 12106 23256 12112
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22192 9862 22244 9868
rect 22282 9888 22338 9897
rect 22204 8566 22232 9862
rect 22282 9823 22338 9832
rect 22480 9178 22508 10134
rect 22572 10130 22600 10678
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22664 9994 22692 10406
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22296 7410 22324 8910
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 18064 800 18092 2382
rect 19352 800 19380 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2382
rect 21284 800 21312 2382
rect 22572 800 22600 2994
rect 22664 2582 22692 9522
rect 22756 8566 22784 9590
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22940 3194 22968 8910
rect 23204 7948 23256 7954
rect 23204 7890 23256 7896
rect 23216 7410 23244 7890
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23308 6322 23336 13806
rect 23584 12782 23612 14214
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23676 12102 23704 13806
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23768 11830 23796 23122
rect 23952 22094 23980 23734
rect 23952 22066 24072 22094
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23952 21010 23980 21626
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23952 20534 23980 20946
rect 23940 20528 23992 20534
rect 23940 20470 23992 20476
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 17270 23888 18634
rect 23952 18290 23980 19246
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23952 17678 23980 18226
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 23952 12306 23980 15914
rect 24044 15706 24072 22066
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24136 19378 24164 20402
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24228 18970 24256 33390
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 24320 22642 24348 24006
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24214 18456 24270 18465
rect 24214 18391 24270 18400
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 24228 15502 24256 18391
rect 24320 17066 24348 22578
rect 24412 18426 24440 33866
rect 24492 33584 24544 33590
rect 24492 33526 24544 33532
rect 24504 24857 24532 33526
rect 24596 32910 24624 34410
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 24688 31754 24716 36790
rect 24768 36712 24820 36718
rect 24768 36654 24820 36660
rect 24780 36242 24808 36654
rect 25136 36576 25188 36582
rect 25136 36518 25188 36524
rect 25228 36576 25280 36582
rect 25228 36518 25280 36524
rect 25148 36242 25176 36518
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 25136 36236 25188 36242
rect 25136 36178 25188 36184
rect 25240 36038 25268 36518
rect 25228 36032 25280 36038
rect 25228 35974 25280 35980
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24596 31726 24716 31754
rect 24490 24848 24546 24857
rect 24490 24783 24546 24792
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24504 22166 24532 22646
rect 24492 22160 24544 22166
rect 24492 22102 24544 22108
rect 24492 20868 24544 20874
rect 24492 20810 24544 20816
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24308 17060 24360 17066
rect 24308 17002 24360 17008
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24504 12374 24532 20810
rect 24596 19514 24624 31726
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24688 30394 24716 30874
rect 24676 30388 24728 30394
rect 24676 30330 24728 30336
rect 24676 25968 24728 25974
rect 24676 25910 24728 25916
rect 24688 20534 24716 25910
rect 24780 22250 24808 34614
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 24952 33652 25004 33658
rect 24952 33594 25004 33600
rect 24964 31822 24992 33594
rect 25044 33584 25096 33590
rect 25044 33526 25096 33532
rect 25056 33046 25084 33526
rect 25424 33318 25452 33934
rect 25412 33312 25464 33318
rect 25412 33254 25464 33260
rect 25044 33040 25096 33046
rect 25044 32982 25096 32988
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 25516 31754 25544 36790
rect 26068 36145 26096 37198
rect 26436 37126 26464 39200
rect 27724 37262 27752 39200
rect 28172 37392 28224 37398
rect 28172 37334 28224 37340
rect 27712 37256 27764 37262
rect 28080 37256 28132 37262
rect 27712 37198 27764 37204
rect 28078 37224 28080 37233
rect 28132 37224 28134 37233
rect 27528 37188 27580 37194
rect 28078 37159 28134 37168
rect 27528 37130 27580 37136
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 26146 36544 26202 36553
rect 26146 36479 26202 36488
rect 26054 36136 26110 36145
rect 26054 36071 26110 36080
rect 26160 33998 26188 36479
rect 26620 36378 26648 36858
rect 27540 36718 27568 37130
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27804 36712 27856 36718
rect 27804 36654 27856 36660
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 27068 36372 27120 36378
rect 27068 36314 27120 36320
rect 26422 36272 26478 36281
rect 26422 36207 26478 36216
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 26252 36009 26280 36110
rect 26436 36106 26464 36207
rect 27080 36174 27108 36314
rect 27068 36168 27120 36174
rect 27068 36110 27120 36116
rect 26424 36100 26476 36106
rect 26424 36042 26476 36048
rect 26238 36000 26294 36009
rect 26238 35935 26294 35944
rect 27172 34610 27200 36654
rect 27712 36168 27764 36174
rect 27710 36136 27712 36145
rect 27764 36136 27766 36145
rect 27710 36071 27766 36080
rect 27344 35624 27396 35630
rect 27344 35566 27396 35572
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 26238 34504 26294 34513
rect 26238 34439 26294 34448
rect 26148 33992 26200 33998
rect 26148 33934 26200 33940
rect 26252 33561 26280 34439
rect 26238 33552 26294 33561
rect 27172 33522 27200 34546
rect 27356 34202 27384 35566
rect 27436 35556 27488 35562
rect 27436 35498 27488 35504
rect 27344 34196 27396 34202
rect 27344 34138 27396 34144
rect 27448 33930 27476 35498
rect 27436 33924 27488 33930
rect 27436 33866 27488 33872
rect 27528 33924 27580 33930
rect 27528 33866 27580 33872
rect 27448 33658 27476 33866
rect 27436 33652 27488 33658
rect 27436 33594 27488 33600
rect 26238 33487 26294 33496
rect 27160 33516 27212 33522
rect 26252 33454 26280 33487
rect 27160 33458 27212 33464
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 26240 33448 26292 33454
rect 26240 33390 26292 33396
rect 25608 32978 25636 33390
rect 25596 32972 25648 32978
rect 25596 32914 25648 32920
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 26160 31754 26188 32370
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 25332 31726 25544 31754
rect 26068 31726 26188 31754
rect 25228 30592 25280 30598
rect 25228 30534 25280 30540
rect 25044 26240 25096 26246
rect 25044 26182 25096 26188
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24872 23866 24900 25774
rect 25056 25362 25084 26182
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 24952 25220 25004 25226
rect 24952 25162 25004 25168
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24780 22222 24900 22250
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 24780 21690 24808 22102
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24872 21570 24900 22222
rect 24780 21542 24900 21570
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24780 19378 24808 21542
rect 24860 19712 24912 19718
rect 24860 19654 24912 19660
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24872 19310 24900 19654
rect 24964 19514 24992 25162
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24596 18766 24624 19110
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24780 18766 24808 18906
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24780 18358 24808 18702
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24596 15502 24624 17818
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24688 13870 24716 15846
rect 25056 15026 25084 25162
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25148 20874 25176 21286
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 20058 25176 20334
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25148 17678 25176 19994
rect 25240 17882 25268 30534
rect 25332 20641 25360 31726
rect 25412 31408 25464 31414
rect 25412 31350 25464 31356
rect 25424 25226 25452 31350
rect 25872 30592 25924 30598
rect 25872 30534 25924 30540
rect 25884 26246 25912 30534
rect 25962 27704 26018 27713
rect 25962 27639 25964 27648
rect 26016 27639 26018 27648
rect 25964 27610 26016 27616
rect 25872 26240 25924 26246
rect 25872 26182 25924 26188
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25596 25152 25648 25158
rect 25596 25094 25648 25100
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25516 22506 25544 23598
rect 25504 22500 25556 22506
rect 25504 22442 25556 22448
rect 25318 20632 25374 20641
rect 25318 20567 25374 20576
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25424 20398 25452 20538
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25332 19446 25360 19858
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25320 19440 25372 19446
rect 25320 19382 25372 19388
rect 25424 19378 25452 19722
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25332 16182 25360 18022
rect 25320 16176 25372 16182
rect 25320 16118 25372 16124
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25056 14906 25084 14962
rect 25056 14878 25176 14906
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24780 14006 24808 14214
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 12782 24716 13806
rect 24768 12912 24820 12918
rect 24872 12900 24900 14282
rect 24964 14278 24992 14758
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 25056 12918 25084 14758
rect 25148 14618 25176 14878
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 24820 12872 24900 12900
rect 24768 12854 24820 12860
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 24492 12368 24544 12374
rect 24492 12310 24544 12316
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23492 9654 23520 11494
rect 24688 10810 24716 12106
rect 24872 11626 24900 12872
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 25240 12306 25268 15642
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 25240 10674 25268 12242
rect 25424 11830 25452 15302
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25516 10538 25544 22442
rect 25608 22234 25636 25094
rect 25688 23792 25740 23798
rect 25688 23734 25740 23740
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25608 16250 25636 22170
rect 25700 20602 25728 23734
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25792 22642 25820 23054
rect 25964 23044 26016 23050
rect 25964 22986 26016 22992
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25792 22098 25820 22578
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25778 20904 25834 20913
rect 25778 20839 25780 20848
rect 25832 20839 25834 20848
rect 25872 20868 25924 20874
rect 25780 20810 25832 20816
rect 25872 20810 25924 20816
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25700 20369 25728 20402
rect 25686 20360 25742 20369
rect 25686 20295 25742 20304
rect 25884 19854 25912 20810
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 25976 19514 26004 22986
rect 26068 22094 26096 31726
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 26160 29714 26188 30738
rect 26252 30598 26280 32302
rect 26332 32224 26384 32230
rect 26332 32166 26384 32172
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26344 29782 26372 32166
rect 27540 32026 27568 33866
rect 27620 33312 27672 33318
rect 27620 33254 27672 33260
rect 27632 32978 27660 33254
rect 27620 32972 27672 32978
rect 27620 32914 27672 32920
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 27436 31136 27488 31142
rect 27436 31078 27488 31084
rect 26700 30932 26752 30938
rect 26700 30874 26752 30880
rect 26332 29776 26384 29782
rect 26332 29718 26384 29724
rect 26148 29708 26200 29714
rect 26148 29650 26200 29656
rect 26160 29170 26188 29650
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26344 28098 26372 29718
rect 26252 28070 26372 28098
rect 26068 22066 26188 22094
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26068 20398 26096 20878
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 25964 19236 26016 19242
rect 25964 19178 26016 19184
rect 25976 18698 26004 19178
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25976 18290 26004 18634
rect 26054 18456 26110 18465
rect 26054 18391 26056 18400
rect 26108 18391 26110 18400
rect 26056 18362 26108 18368
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25700 17202 25728 17614
rect 26160 17338 26188 22066
rect 26252 21418 26280 28070
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26424 28008 26476 28014
rect 26424 27950 26476 27956
rect 26344 26314 26372 27950
rect 26436 27470 26464 27950
rect 26424 27464 26476 27470
rect 26424 27406 26476 27412
rect 26436 26926 26464 27406
rect 26424 26920 26476 26926
rect 26424 26862 26476 26868
rect 26436 26450 26464 26862
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26436 25906 26464 26386
rect 26608 26036 26660 26042
rect 26608 25978 26660 25984
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26436 25362 26464 25842
rect 26424 25356 26476 25362
rect 26424 25298 26476 25304
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26528 22778 26556 24346
rect 26516 22772 26568 22778
rect 26516 22714 26568 22720
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 26252 20924 26280 21354
rect 26424 21072 26476 21078
rect 26424 21014 26476 21020
rect 26332 20936 26384 20942
rect 26252 20896 26332 20924
rect 26332 20878 26384 20884
rect 26436 20448 26464 21014
rect 26528 20602 26556 22714
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26516 20460 26568 20466
rect 26436 20420 26516 20448
rect 26516 20402 26568 20408
rect 26240 20392 26292 20398
rect 26240 20334 26292 20340
rect 26252 19854 26280 20334
rect 26528 20262 26556 20402
rect 26424 20256 26476 20262
rect 26424 20198 26476 20204
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26252 18630 26280 19314
rect 26332 19168 26384 19174
rect 26330 19136 26332 19145
rect 26384 19136 26386 19145
rect 26330 19071 26386 19080
rect 26330 19000 26386 19009
rect 26330 18935 26332 18944
rect 26384 18935 26386 18944
rect 26332 18906 26384 18912
rect 26436 18834 26464 20198
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 26344 16658 26372 17478
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25976 15502 26004 15846
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26160 15502 26188 15642
rect 26344 15586 26372 16594
rect 26252 15558 26372 15586
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25700 11286 25728 12106
rect 25872 11620 25924 11626
rect 25872 11562 25924 11568
rect 25688 11280 25740 11286
rect 25688 11222 25740 11228
rect 25504 10532 25556 10538
rect 25504 10474 25556 10480
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 9988 24728 9994
rect 24676 9930 24728 9936
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23400 6118 23428 6734
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 24688 2650 24716 9930
rect 24780 8906 24808 10406
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24964 9654 24992 9998
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24860 9580 24912 9586
rect 24860 9522 24912 9528
rect 24768 8900 24820 8906
rect 24768 8842 24820 8848
rect 24872 8498 24900 9522
rect 25516 8974 25544 10474
rect 25884 9450 25912 11562
rect 26252 10266 26280 15558
rect 26620 15026 26648 25978
rect 26712 24342 26740 30874
rect 26884 30048 26936 30054
rect 26884 29990 26936 29996
rect 26896 29510 26924 29990
rect 26884 29504 26936 29510
rect 26884 29446 26936 29452
rect 27344 28960 27396 28966
rect 27344 28902 27396 28908
rect 26884 28144 26936 28150
rect 26884 28086 26936 28092
rect 26700 24336 26752 24342
rect 26700 24278 26752 24284
rect 26712 19378 26740 24278
rect 26792 21888 26844 21894
rect 26792 21830 26844 21836
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26804 15910 26832 21830
rect 26792 15904 26844 15910
rect 26792 15846 26844 15852
rect 26896 15042 26924 28086
rect 27160 27668 27212 27674
rect 27160 27610 27212 27616
rect 26976 27396 27028 27402
rect 26976 27338 27028 27344
rect 26988 23866 27016 27338
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 26988 18698 27016 19382
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26804 15026 26924 15042
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26804 15020 26936 15026
rect 26804 15014 26884 15020
rect 26620 14550 26648 14962
rect 26608 14544 26660 14550
rect 26608 14486 26660 14492
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26332 13728 26384 13734
rect 26332 13670 26384 13676
rect 26344 13394 26372 13670
rect 26712 13462 26740 14418
rect 26804 14414 26832 15014
rect 26884 14962 26936 14968
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26896 14482 26924 14826
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26792 14408 26844 14414
rect 26988 14362 27016 18634
rect 27080 18358 27108 22986
rect 27172 21894 27200 27610
rect 27356 23361 27384 28902
rect 27448 28150 27476 31078
rect 27620 30252 27672 30258
rect 27620 30194 27672 30200
rect 27632 29646 27660 30194
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27436 28144 27488 28150
rect 27436 28086 27488 28092
rect 27632 26994 27660 29582
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27436 26512 27488 26518
rect 27436 26454 27488 26460
rect 27448 26353 27476 26454
rect 27434 26344 27490 26353
rect 27434 26279 27490 26288
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 27342 23352 27398 23361
rect 27342 23287 27398 23296
rect 27448 22710 27476 25638
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27448 22094 27476 22646
rect 27264 22066 27476 22094
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 26792 14350 26844 14356
rect 26896 14334 27016 14362
rect 26700 13456 26752 13462
rect 26700 13398 26752 13404
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25872 9444 25924 9450
rect 25872 9386 25924 9392
rect 25504 8968 25556 8974
rect 25504 8910 25556 8916
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24872 7410 24900 8434
rect 25976 7410 26004 9454
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 26528 7410 26556 8230
rect 26620 7546 26648 12038
rect 26896 9382 26924 14334
rect 27172 13326 27200 20538
rect 27264 19530 27292 22066
rect 27436 21956 27488 21962
rect 27436 21898 27488 21904
rect 27448 19990 27476 21898
rect 27540 20058 27568 25162
rect 27632 24750 27660 26930
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27632 24274 27660 24686
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 27264 19502 27384 19530
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27264 17610 27292 19314
rect 27252 17604 27304 17610
rect 27252 17546 27304 17552
rect 27356 16658 27384 19502
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27448 18834 27476 19314
rect 27436 18828 27488 18834
rect 27436 18770 27488 18776
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27448 18426 27476 18634
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27264 15502 27292 16390
rect 27448 15910 27476 16730
rect 27436 15904 27488 15910
rect 27436 15846 27488 15852
rect 27252 15496 27304 15502
rect 27252 15438 27304 15444
rect 27540 15026 27568 17478
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27632 14346 27660 16390
rect 27724 15026 27752 31758
rect 27816 18970 27844 36654
rect 27986 36272 28042 36281
rect 27986 36207 27988 36216
rect 28040 36207 28042 36216
rect 27988 36178 28040 36184
rect 28092 31890 28120 37159
rect 28184 36174 28212 37334
rect 28264 36848 28316 36854
rect 28264 36790 28316 36796
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 28080 31884 28132 31890
rect 28080 31826 28132 31832
rect 28276 31754 28304 36790
rect 28816 36644 28868 36650
rect 28816 36586 28868 36592
rect 28828 36553 28856 36586
rect 28814 36544 28870 36553
rect 28814 36479 28870 36488
rect 28446 36272 28502 36281
rect 28446 36207 28448 36216
rect 28500 36207 28502 36216
rect 28448 36178 28500 36184
rect 29012 36174 29040 39200
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 29104 36582 29132 37266
rect 29656 36922 29684 39200
rect 30944 37466 30972 39200
rect 30932 37460 30984 37466
rect 30932 37402 30984 37408
rect 31300 37256 31352 37262
rect 31298 37224 31300 37233
rect 31576 37256 31628 37262
rect 31352 37224 31354 37233
rect 30380 37188 30432 37194
rect 30380 37130 30432 37136
rect 30748 37188 30800 37194
rect 31576 37198 31628 37204
rect 31298 37159 31354 37168
rect 30748 37130 30800 37136
rect 29644 36916 29696 36922
rect 29644 36858 29696 36864
rect 30392 36854 30420 37130
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 30380 36848 30432 36854
rect 30380 36790 30432 36796
rect 29828 36712 29880 36718
rect 29828 36654 29880 36660
rect 29840 36582 29868 36654
rect 29092 36576 29144 36582
rect 29092 36518 29144 36524
rect 29828 36576 29880 36582
rect 29828 36518 29880 36524
rect 29092 36236 29144 36242
rect 29092 36178 29144 36184
rect 29000 36168 29052 36174
rect 28630 36136 28686 36145
rect 29000 36110 29052 36116
rect 28630 36071 28686 36080
rect 28644 36038 28672 36071
rect 28356 36032 28408 36038
rect 28354 36000 28356 36009
rect 28448 36032 28500 36038
rect 28408 36000 28410 36009
rect 28448 35974 28500 35980
rect 28632 36032 28684 36038
rect 28632 35974 28684 35980
rect 28354 35935 28410 35944
rect 28460 34048 28488 35974
rect 28724 35488 28776 35494
rect 28724 35430 28776 35436
rect 28736 34785 28764 35430
rect 29104 35154 29132 36178
rect 30484 36174 30512 37062
rect 30564 36848 30616 36854
rect 30564 36790 30616 36796
rect 30472 36168 30524 36174
rect 30472 36110 30524 36116
rect 29184 36032 29236 36038
rect 29182 36000 29184 36009
rect 29236 36000 29238 36009
rect 29182 35935 29238 35944
rect 29276 35828 29328 35834
rect 29276 35770 29328 35776
rect 29092 35148 29144 35154
rect 29092 35090 29144 35096
rect 28722 34776 28778 34785
rect 28722 34711 28778 34720
rect 28538 34640 28594 34649
rect 28538 34575 28540 34584
rect 28592 34575 28594 34584
rect 28540 34546 28592 34552
rect 29288 34542 29316 35770
rect 30288 35012 30340 35018
rect 30288 34954 30340 34960
rect 30012 34604 30064 34610
rect 30012 34546 30064 34552
rect 29184 34536 29236 34542
rect 29184 34478 29236 34484
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 29000 34400 29052 34406
rect 29000 34342 29052 34348
rect 28368 34020 28488 34048
rect 28368 32842 28396 34020
rect 28448 33924 28500 33930
rect 28448 33866 28500 33872
rect 28460 33289 28488 33866
rect 28724 33448 28776 33454
rect 28724 33390 28776 33396
rect 28446 33280 28502 33289
rect 28446 33215 28502 33224
rect 28448 32972 28500 32978
rect 28448 32914 28500 32920
rect 28460 32881 28488 32914
rect 28446 32872 28502 32881
rect 28356 32836 28408 32842
rect 28446 32807 28448 32816
rect 28356 32778 28408 32784
rect 28500 32807 28502 32816
rect 28448 32778 28500 32784
rect 28460 32747 28488 32778
rect 28736 32570 28764 33390
rect 28724 32564 28776 32570
rect 28724 32506 28776 32512
rect 28184 31726 28304 31754
rect 28080 25968 28132 25974
rect 28080 25910 28132 25916
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 27908 18766 27936 20810
rect 27986 19272 28042 19281
rect 27986 19207 28042 19216
rect 28000 18834 28028 19207
rect 27988 18828 28040 18834
rect 27988 18770 28040 18776
rect 27896 18760 27948 18766
rect 27896 18702 27948 18708
rect 27908 17678 27936 18702
rect 28092 17882 28120 25910
rect 28184 20602 28212 31726
rect 28632 30660 28684 30666
rect 28632 30602 28684 30608
rect 28264 29232 28316 29238
rect 28264 29174 28316 29180
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28172 20392 28224 20398
rect 28172 20334 28224 20340
rect 28184 19242 28212 20334
rect 28276 19972 28304 29174
rect 28540 25764 28592 25770
rect 28540 25706 28592 25712
rect 28552 24750 28580 25706
rect 28540 24744 28592 24750
rect 28368 24704 28540 24732
rect 28368 20074 28396 24704
rect 28540 24686 28592 24692
rect 28448 22704 28500 22710
rect 28448 22646 28500 22652
rect 28460 20346 28488 22646
rect 28538 20632 28594 20641
rect 28538 20567 28594 20576
rect 28552 20534 28580 20567
rect 28644 20534 28672 30602
rect 29012 29034 29040 34342
rect 29196 29850 29224 34478
rect 30024 33590 30052 34546
rect 30300 34202 30328 34954
rect 30484 34678 30512 36110
rect 30576 36009 30604 36790
rect 30562 36000 30618 36009
rect 30562 35935 30618 35944
rect 30472 34672 30524 34678
rect 30472 34614 30524 34620
rect 30288 34196 30340 34202
rect 30288 34138 30340 34144
rect 30484 34066 30512 34614
rect 30472 34060 30524 34066
rect 30472 34002 30524 34008
rect 30012 33584 30064 33590
rect 30012 33526 30064 33532
rect 29828 33516 29880 33522
rect 29828 33458 29880 33464
rect 29840 33289 29868 33458
rect 29920 33448 29972 33454
rect 29920 33390 29972 33396
rect 29826 33280 29882 33289
rect 29826 33215 29882 33224
rect 29644 30388 29696 30394
rect 29644 30330 29696 30336
rect 29184 29844 29236 29850
rect 29184 29786 29236 29792
rect 29656 29578 29684 30330
rect 29736 30184 29788 30190
rect 29736 30126 29788 30132
rect 29748 29714 29776 30126
rect 29736 29708 29788 29714
rect 29736 29650 29788 29656
rect 29644 29572 29696 29578
rect 29644 29514 29696 29520
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 29276 29028 29328 29034
rect 29276 28970 29328 28976
rect 28724 28144 28776 28150
rect 28724 28086 28776 28092
rect 29184 28144 29236 28150
rect 29184 28086 29236 28092
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28632 20528 28684 20534
rect 28632 20470 28684 20476
rect 28460 20318 28672 20346
rect 28368 20046 28580 20074
rect 28356 19984 28408 19990
rect 28276 19944 28356 19972
rect 28356 19926 28408 19932
rect 28172 19236 28224 19242
rect 28172 19178 28224 19184
rect 28184 18290 28212 19178
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 28184 17678 28212 18226
rect 28448 18080 28500 18086
rect 28448 18022 28500 18028
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28262 16824 28318 16833
rect 28262 16759 28264 16768
rect 28316 16759 28318 16768
rect 28264 16730 28316 16736
rect 28356 16720 28408 16726
rect 28356 16662 28408 16668
rect 27804 16176 27856 16182
rect 27804 16118 27856 16124
rect 27988 16176 28040 16182
rect 27988 16118 28040 16124
rect 27816 15706 27844 16118
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27710 14376 27766 14385
rect 27620 14340 27672 14346
rect 27710 14311 27766 14320
rect 27620 14282 27672 14288
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26988 12646 27016 13126
rect 27632 12850 27660 13806
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 27252 11688 27304 11694
rect 27252 11630 27304 11636
rect 27264 10606 27292 11630
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 27356 10742 27384 11494
rect 27344 10736 27396 10742
rect 27344 10678 27396 10684
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27724 9926 27752 14311
rect 27816 14006 27844 15302
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27712 9920 27764 9926
rect 27712 9862 27764 9868
rect 28000 9654 28028 16118
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28184 15366 28212 15438
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 28276 12850 28304 13466
rect 28264 12844 28316 12850
rect 28264 12786 28316 12792
rect 28368 10742 28396 16662
rect 28460 16182 28488 18022
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28552 15892 28580 20046
rect 28644 19718 28672 20318
rect 28632 19712 28684 19718
rect 28632 19654 28684 19660
rect 28736 18426 28764 28086
rect 29092 27396 29144 27402
rect 29092 27338 29144 27344
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29012 24138 29040 24550
rect 29000 24132 29052 24138
rect 29000 24074 29052 24080
rect 28908 23656 28960 23662
rect 28908 23598 28960 23604
rect 28920 22574 28948 23598
rect 29012 23526 29040 24074
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 29012 23186 29040 23462
rect 29000 23180 29052 23186
rect 29000 23122 29052 23128
rect 29012 22778 29040 23122
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 28908 22568 28960 22574
rect 28908 22510 28960 22516
rect 28920 21622 28948 22510
rect 28908 21616 28960 21622
rect 28908 21558 28960 21564
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28920 20942 28948 21422
rect 29104 21146 29132 27338
rect 29092 21140 29144 21146
rect 29092 21082 29144 21088
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 28816 20460 28868 20466
rect 28816 20402 28868 20408
rect 28828 19854 28856 20402
rect 28908 20392 28960 20398
rect 28906 20360 28908 20369
rect 28960 20360 28962 20369
rect 28906 20295 28962 20304
rect 28906 20088 28962 20097
rect 28906 20023 28908 20032
rect 28960 20023 28962 20032
rect 28908 19994 28960 20000
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 29012 19514 29040 19722
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 29196 19360 29224 28086
rect 29288 19446 29316 28970
rect 29656 28150 29684 29514
rect 29644 28144 29696 28150
rect 29644 28086 29696 28092
rect 29368 26920 29420 26926
rect 29368 26862 29420 26868
rect 29380 25906 29408 26862
rect 29552 26308 29604 26314
rect 29552 26250 29604 26256
rect 29368 25900 29420 25906
rect 29368 25842 29420 25848
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29276 19440 29328 19446
rect 29276 19382 29328 19388
rect 29104 19332 29224 19360
rect 28908 19304 28960 19310
rect 29000 19304 29052 19310
rect 28908 19246 28960 19252
rect 28998 19272 29000 19281
rect 29052 19272 29054 19281
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 28828 18290 28856 18906
rect 28920 18426 28948 19246
rect 28998 19207 29054 19216
rect 29012 19174 29040 19207
rect 29000 19168 29052 19174
rect 29000 19110 29052 19116
rect 28908 18420 28960 18426
rect 28908 18362 28960 18368
rect 28816 18284 28868 18290
rect 28816 18226 28868 18232
rect 28630 17912 28686 17921
rect 28630 17847 28632 17856
rect 28684 17847 28686 17856
rect 28632 17818 28684 17824
rect 29000 17604 29052 17610
rect 29000 17546 29052 17552
rect 29012 16425 29040 17546
rect 29104 16658 29132 19332
rect 29182 17368 29238 17377
rect 29182 17303 29184 17312
rect 29236 17303 29238 17312
rect 29184 17274 29236 17280
rect 29092 16652 29144 16658
rect 29092 16594 29144 16600
rect 28998 16416 29054 16425
rect 28998 16351 29054 16360
rect 28552 15864 28672 15892
rect 28446 15464 28502 15473
rect 28446 15399 28448 15408
rect 28500 15399 28502 15408
rect 28448 15370 28500 15376
rect 28540 14952 28592 14958
rect 28540 14894 28592 14900
rect 28552 14618 28580 14894
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28540 14612 28592 14618
rect 28540 14554 28592 14560
rect 28460 14414 28488 14554
rect 28448 14408 28500 14414
rect 28448 14350 28500 14356
rect 28538 14376 28594 14385
rect 28538 14311 28540 14320
rect 28592 14311 28594 14320
rect 28540 14282 28592 14288
rect 28446 13560 28502 13569
rect 28644 13530 28672 15864
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 28828 15558 29224 15586
rect 28828 15162 28856 15558
rect 29196 15502 29224 15558
rect 29184 15496 29236 15502
rect 29184 15438 29236 15444
rect 28908 15428 28960 15434
rect 28908 15370 28960 15376
rect 28920 15314 28948 15370
rect 28920 15286 29040 15314
rect 29012 15162 29040 15286
rect 28816 15156 28868 15162
rect 28816 15098 28868 15104
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 29288 15026 29316 15642
rect 29276 15020 29328 15026
rect 29276 14962 29328 14968
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 28446 13495 28448 13504
rect 28500 13495 28502 13504
rect 28632 13524 28684 13530
rect 28448 13466 28500 13472
rect 28632 13466 28684 13472
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 29012 12850 29040 13126
rect 29104 12986 29132 13874
rect 29288 13818 29316 14962
rect 29196 13790 29316 13818
rect 29092 12980 29144 12986
rect 29092 12922 29144 12928
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 29196 12714 29224 13790
rect 29276 13728 29328 13734
rect 29276 13670 29328 13676
rect 29288 13394 29316 13670
rect 29276 13388 29328 13394
rect 29276 13330 29328 13336
rect 29184 12708 29236 12714
rect 29184 12650 29236 12656
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 28356 10736 28408 10742
rect 28356 10678 28408 10684
rect 27988 9648 28040 9654
rect 27988 9590 28040 9596
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 28368 9042 28396 10678
rect 28920 10674 28948 10950
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29104 9722 29132 10542
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28356 9036 28408 9042
rect 28356 8978 28408 8984
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 27724 8566 27752 8774
rect 28368 8566 28396 8978
rect 28920 8634 28948 9522
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 27712 8560 27764 8566
rect 27712 8502 27764 8508
rect 28356 8560 28408 8566
rect 28356 8502 28408 8508
rect 29380 8498 29408 22986
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29472 19922 29500 20402
rect 29460 19916 29512 19922
rect 29460 19858 29512 19864
rect 29564 18970 29592 26250
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29644 24676 29696 24682
rect 29644 24618 29696 24624
rect 29656 24342 29684 24618
rect 29644 24336 29696 24342
rect 29644 24278 29696 24284
rect 29840 21146 29868 24754
rect 29932 23050 29960 33390
rect 30024 30258 30052 33526
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 30392 30190 30420 31758
rect 30760 31754 30788 37130
rect 31300 36576 31352 36582
rect 31300 36518 31352 36524
rect 31116 36100 31168 36106
rect 31116 36042 31168 36048
rect 31022 34640 31078 34649
rect 31022 34575 31024 34584
rect 31076 34575 31078 34584
rect 31024 34546 31076 34552
rect 31128 33998 31156 36042
rect 31312 36038 31340 36518
rect 31300 36032 31352 36038
rect 31300 35974 31352 35980
rect 31588 35834 31616 37198
rect 31668 37120 31720 37126
rect 31668 37062 31720 37068
rect 31680 36922 31708 37062
rect 31668 36916 31720 36922
rect 31668 36858 31720 36864
rect 32232 36854 32260 39200
rect 32876 37346 32904 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 32876 37318 33088 37346
rect 32956 37256 33008 37262
rect 32956 37198 33008 37204
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 32220 36848 32272 36854
rect 32220 36790 32272 36796
rect 32312 36576 32364 36582
rect 32312 36518 32364 36524
rect 32404 36576 32456 36582
rect 32404 36518 32456 36524
rect 31576 35828 31628 35834
rect 31576 35770 31628 35776
rect 31484 35692 31536 35698
rect 31484 35634 31536 35640
rect 31208 35012 31260 35018
rect 31208 34954 31260 34960
rect 31220 34649 31248 34954
rect 31496 34746 31524 35634
rect 32324 35290 32352 36518
rect 32416 36378 32444 36518
rect 32508 36378 32536 36858
rect 32404 36372 32456 36378
rect 32404 36314 32456 36320
rect 32496 36372 32548 36378
rect 32496 36314 32548 36320
rect 32588 36032 32640 36038
rect 32588 35974 32640 35980
rect 32312 35284 32364 35290
rect 32312 35226 32364 35232
rect 32600 35018 32628 35974
rect 32968 35894 32996 37198
rect 33060 37108 33088 37318
rect 33692 37256 33744 37262
rect 33692 37198 33744 37204
rect 33508 37188 33560 37194
rect 33508 37130 33560 37136
rect 33140 37120 33192 37126
rect 33060 37080 33140 37108
rect 33140 37062 33192 37068
rect 33140 36644 33192 36650
rect 33140 36586 33192 36592
rect 32876 35866 32996 35894
rect 33152 35894 33180 36586
rect 33520 36174 33548 37130
rect 33704 36242 33732 37198
rect 34440 37108 34468 39222
rect 35438 39200 35494 39800
rect 36082 39200 36138 39800
rect 37370 39200 37426 39800
rect 38658 39200 38714 39800
rect 39302 39200 39358 39800
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 34520 37062 34572 37068
rect 34060 36848 34112 36854
rect 34060 36790 34112 36796
rect 33692 36236 33744 36242
rect 33692 36178 33744 36184
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33152 35866 33272 35894
rect 32588 35012 32640 35018
rect 32588 34954 32640 34960
rect 31484 34740 31536 34746
rect 31484 34682 31536 34688
rect 31206 34640 31262 34649
rect 31206 34575 31262 34584
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 31128 33862 31156 33934
rect 32128 33924 32180 33930
rect 32128 33866 32180 33872
rect 31116 33856 31168 33862
rect 31116 33798 31168 33804
rect 31128 33522 31156 33798
rect 31116 33516 31168 33522
rect 31116 33458 31168 33464
rect 30668 31726 30788 31754
rect 30380 30184 30432 30190
rect 30380 30126 30432 30132
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30484 27878 30512 29650
rect 30472 27872 30524 27878
rect 30472 27814 30524 27820
rect 30472 27396 30524 27402
rect 30472 27338 30524 27344
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 30196 26784 30248 26790
rect 30196 26726 30248 26732
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 30024 24410 30052 24550
rect 30012 24404 30064 24410
rect 30012 24346 30064 24352
rect 29920 23044 29972 23050
rect 29920 22986 29972 22992
rect 30208 22094 30236 26726
rect 30392 25498 30420 26862
rect 30380 25492 30432 25498
rect 30380 25434 30432 25440
rect 30288 23792 30340 23798
rect 30288 23734 30340 23740
rect 30116 22066 30236 22094
rect 29828 21140 29880 21146
rect 29828 21082 29880 21088
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29748 20602 29776 20878
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29748 20262 29776 20538
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29736 19984 29788 19990
rect 29734 19952 29736 19961
rect 29788 19952 29790 19961
rect 29734 19887 29790 19896
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 29840 19689 29868 19858
rect 29932 19786 29960 20742
rect 29920 19780 29972 19786
rect 29920 19722 29972 19728
rect 29826 19680 29882 19689
rect 29826 19615 29882 19624
rect 29734 19272 29790 19281
rect 29734 19207 29790 19216
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29748 18766 29776 19207
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 30024 18630 30052 20742
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29840 16454 29868 17546
rect 29920 16992 29972 16998
rect 29920 16934 29972 16940
rect 29460 16448 29512 16454
rect 29460 16390 29512 16396
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 29472 16182 29500 16390
rect 29840 16250 29868 16390
rect 29828 16244 29880 16250
rect 29828 16186 29880 16192
rect 29460 16176 29512 16182
rect 29460 16118 29512 16124
rect 29932 16046 29960 16934
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29472 14822 29500 15982
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29748 14414 29776 14486
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29460 14272 29512 14278
rect 29460 14214 29512 14220
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 29472 13394 29500 14214
rect 30024 14006 30052 14214
rect 30012 14000 30064 14006
rect 30012 13942 30064 13948
rect 30116 13938 30144 22066
rect 30300 19514 30328 23734
rect 30380 23520 30432 23526
rect 30378 23488 30380 23497
rect 30432 23488 30434 23497
rect 30378 23423 30434 23432
rect 30484 23186 30512 27338
rect 30564 26444 30616 26450
rect 30564 26386 30616 26392
rect 30576 25362 30604 26386
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30564 24132 30616 24138
rect 30564 24074 30616 24080
rect 30472 23180 30524 23186
rect 30472 23122 30524 23128
rect 30576 21690 30604 24074
rect 30668 23526 30696 31726
rect 31208 29844 31260 29850
rect 31208 29786 31260 29792
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30852 26518 30880 26794
rect 30840 26512 30892 26518
rect 30840 26454 30892 26460
rect 30748 25900 30800 25906
rect 30748 25842 30800 25848
rect 30656 23520 30708 23526
rect 30656 23462 30708 23468
rect 30656 23180 30708 23186
rect 30656 23122 30708 23128
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 30472 21412 30524 21418
rect 30472 21354 30524 21360
rect 30484 21010 30512 21354
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30378 20632 30434 20641
rect 30378 20567 30434 20576
rect 30392 20466 30420 20567
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30484 19922 30512 20946
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 30288 19508 30340 19514
rect 30288 19450 30340 19456
rect 30208 18714 30236 19450
rect 30564 19304 30616 19310
rect 30564 19246 30616 19252
rect 30576 18834 30604 19246
rect 30564 18828 30616 18834
rect 30564 18770 30616 18776
rect 30286 18728 30342 18737
rect 30208 18686 30286 18714
rect 30286 18663 30342 18672
rect 30196 17264 30248 17270
rect 30196 17206 30248 17212
rect 30208 14074 30236 17206
rect 30300 17134 30328 18663
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 30484 17882 30512 18226
rect 30472 17876 30524 17882
rect 30472 17818 30524 17824
rect 30564 17808 30616 17814
rect 30378 17776 30434 17785
rect 30564 17750 30616 17756
rect 30378 17711 30380 17720
rect 30432 17711 30434 17720
rect 30380 17682 30432 17688
rect 30576 17134 30604 17750
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30564 17128 30616 17134
rect 30564 17070 30616 17076
rect 30380 17060 30432 17066
rect 30380 17002 30432 17008
rect 30288 16516 30340 16522
rect 30288 16458 30340 16464
rect 30300 16250 30328 16458
rect 30288 16244 30340 16250
rect 30288 16186 30340 16192
rect 30392 16046 30420 17002
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30288 15020 30340 15026
rect 30288 14962 30340 14968
rect 30300 14890 30328 14962
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 29460 13388 29512 13394
rect 29460 13330 29512 13336
rect 30116 12434 30144 13874
rect 30116 12406 30236 12434
rect 29828 12300 29880 12306
rect 29828 12242 29880 12248
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29656 11354 29684 12174
rect 29644 11348 29696 11354
rect 29644 11290 29696 11296
rect 29840 10810 29868 12242
rect 30208 11626 30236 12406
rect 30196 11620 30248 11626
rect 30196 11562 30248 11568
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29840 10198 29868 10746
rect 29828 10192 29880 10198
rect 29828 10134 29880 10140
rect 29734 9888 29790 9897
rect 29734 9823 29790 9832
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 27724 8022 27752 8366
rect 27712 8016 27764 8022
rect 27712 7958 27764 7964
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24780 6798 24808 7142
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 25976 5370 26004 7346
rect 26620 6866 26648 7482
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26344 5710 26372 6054
rect 26332 5704 26384 5710
rect 26332 5646 26384 5652
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 27172 2650 27200 7822
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 24676 2644 24728 2650
rect 24676 2586 24728 2592
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 23216 800 23244 2382
rect 24504 800 24532 2382
rect 25792 800 25820 2382
rect 27080 800 27108 2382
rect 27632 2310 27660 5170
rect 27816 2446 27844 7686
rect 28908 5568 28960 5574
rect 28908 5510 28960 5516
rect 28920 3058 28948 5510
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 29748 2446 29776 9823
rect 30300 8906 30328 14554
rect 30392 14550 30420 15982
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30484 15094 30512 15302
rect 30472 15088 30524 15094
rect 30472 15030 30524 15036
rect 30564 14816 30616 14822
rect 30564 14758 30616 14764
rect 30380 14544 30432 14550
rect 30380 14486 30432 14492
rect 30392 13870 30420 14486
rect 30576 14346 30604 14758
rect 30472 14340 30524 14346
rect 30472 14282 30524 14288
rect 30564 14340 30616 14346
rect 30564 14282 30616 14288
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30484 13530 30512 14282
rect 30564 14000 30616 14006
rect 30564 13942 30616 13948
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 30392 11898 30420 12718
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30484 10266 30512 13194
rect 30472 10260 30524 10266
rect 30472 10202 30524 10208
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30104 8900 30156 8906
rect 30104 8842 30156 8848
rect 30288 8900 30340 8906
rect 30288 8842 30340 8848
rect 30116 8634 30144 8842
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 29840 6322 29868 6598
rect 29828 6316 29880 6322
rect 29828 6258 29880 6264
rect 30392 2922 30420 9998
rect 30576 9042 30604 13942
rect 30668 12374 30696 23122
rect 30760 21146 30788 25842
rect 30840 25696 30892 25702
rect 30840 25638 30892 25644
rect 30852 25226 30880 25638
rect 30840 25220 30892 25226
rect 30840 25162 30892 25168
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 30760 18766 30788 19790
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30760 18358 30788 18702
rect 30748 18352 30800 18358
rect 30748 18294 30800 18300
rect 30852 17218 30880 25162
rect 30760 17190 30880 17218
rect 30656 12368 30708 12374
rect 30656 12310 30708 12316
rect 30668 11150 30696 12310
rect 30760 11830 30788 17190
rect 30944 15910 30972 27814
rect 31116 27532 31168 27538
rect 31116 27474 31168 27480
rect 31024 26920 31076 26926
rect 31024 26862 31076 26868
rect 31036 22094 31064 26862
rect 31128 26450 31156 27474
rect 31116 26444 31168 26450
rect 31116 26386 31168 26392
rect 31036 22066 31156 22094
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 31036 19922 31064 21490
rect 31128 20602 31156 22066
rect 31220 21962 31248 29786
rect 31392 29572 31444 29578
rect 31392 29514 31444 29520
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 31312 26790 31340 29242
rect 31300 26784 31352 26790
rect 31300 26726 31352 26732
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31220 21554 31248 21898
rect 31208 21548 31260 21554
rect 31208 21490 31260 21496
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 31300 20324 31352 20330
rect 31300 20266 31352 20272
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 31116 19372 31168 19378
rect 31116 19314 31168 19320
rect 31128 18766 31156 19314
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31024 17808 31076 17814
rect 31024 17750 31076 17756
rect 31036 16794 31064 17750
rect 31128 16998 31156 18702
rect 31220 18358 31248 20198
rect 31312 19854 31340 20266
rect 31404 20058 31432 29514
rect 31668 27396 31720 27402
rect 31668 27338 31720 27344
rect 31680 27130 31708 27338
rect 31760 27328 31812 27334
rect 31760 27270 31812 27276
rect 31668 27124 31720 27130
rect 31668 27066 31720 27072
rect 31772 26314 31800 27270
rect 31760 26308 31812 26314
rect 31760 26250 31812 26256
rect 31852 25220 31904 25226
rect 31852 25162 31904 25168
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31496 22574 31524 24006
rect 31576 23112 31628 23118
rect 31576 23054 31628 23060
rect 31484 22568 31536 22574
rect 31484 22510 31536 22516
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31300 19848 31352 19854
rect 31300 19790 31352 19796
rect 31484 19848 31536 19854
rect 31484 19790 31536 19796
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 31312 18358 31340 19110
rect 31208 18352 31260 18358
rect 31208 18294 31260 18300
rect 31300 18352 31352 18358
rect 31300 18294 31352 18300
rect 31392 18216 31444 18222
rect 31392 18158 31444 18164
rect 31404 17746 31432 18158
rect 31392 17740 31444 17746
rect 31392 17682 31444 17688
rect 31116 16992 31168 16998
rect 31116 16934 31168 16940
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31404 16658 31432 17682
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31206 16280 31262 16289
rect 31206 16215 31262 16224
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 30932 15904 30984 15910
rect 30932 15846 30984 15852
rect 30944 15502 30972 15846
rect 31036 15706 31064 16050
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 31220 15502 31248 16215
rect 30932 15496 30984 15502
rect 30932 15438 30984 15444
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 30840 14952 30892 14958
rect 30838 14920 30840 14929
rect 31024 14952 31076 14958
rect 30892 14920 30894 14929
rect 31024 14894 31076 14900
rect 30838 14855 30894 14864
rect 31036 14550 31064 14894
rect 31024 14544 31076 14550
rect 31024 14486 31076 14492
rect 31128 14362 31156 15302
rect 31206 14920 31262 14929
rect 31206 14855 31262 14864
rect 30944 14334 31156 14362
rect 30840 14272 30892 14278
rect 30840 14214 30892 14220
rect 30748 11824 30800 11830
rect 30748 11766 30800 11772
rect 30760 11558 30788 11766
rect 30748 11552 30800 11558
rect 30748 11494 30800 11500
rect 30656 11144 30708 11150
rect 30656 11086 30708 11092
rect 30564 9036 30616 9042
rect 30564 8978 30616 8984
rect 30576 6866 30604 8978
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30852 6730 30880 14214
rect 30944 11830 30972 14334
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 31036 13326 31064 13806
rect 31220 13394 31248 14855
rect 31300 14816 31352 14822
rect 31300 14758 31352 14764
rect 31312 14618 31340 14758
rect 31300 14612 31352 14618
rect 31300 14554 31352 14560
rect 31300 13728 31352 13734
rect 31300 13670 31352 13676
rect 31208 13388 31260 13394
rect 31208 13330 31260 13336
rect 31024 13320 31076 13326
rect 31024 13262 31076 13268
rect 31036 12442 31064 13262
rect 31312 13190 31340 13670
rect 31300 13184 31352 13190
rect 31300 13126 31352 13132
rect 31312 12850 31340 13126
rect 31496 12850 31524 19790
rect 31588 19446 31616 23054
rect 31668 22568 31720 22574
rect 31668 22510 31720 22516
rect 31576 19440 31628 19446
rect 31576 19382 31628 19388
rect 31680 19122 31708 22510
rect 31864 21146 31892 25162
rect 31944 24744 31996 24750
rect 31944 24686 31996 24692
rect 31956 23662 31984 24686
rect 31944 23656 31996 23662
rect 31944 23598 31996 23604
rect 31956 23118 31984 23598
rect 31944 23112 31996 23118
rect 31944 23054 31996 23060
rect 31956 22642 31984 23054
rect 32036 22976 32088 22982
rect 32036 22918 32088 22924
rect 31944 22636 31996 22642
rect 31944 22578 31996 22584
rect 31956 22098 31984 22578
rect 31944 22092 31996 22098
rect 31944 22034 31996 22040
rect 31944 21344 31996 21350
rect 31944 21286 31996 21292
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 31956 20942 31984 21286
rect 31944 20936 31996 20942
rect 31944 20878 31996 20884
rect 31944 20528 31996 20534
rect 31942 20496 31944 20505
rect 31996 20496 31998 20505
rect 31942 20431 31998 20440
rect 31944 19984 31996 19990
rect 31944 19926 31996 19932
rect 31956 19378 31984 19926
rect 31944 19372 31996 19378
rect 31944 19314 31996 19320
rect 31588 19094 31708 19122
rect 31588 16182 31616 19094
rect 31668 18148 31720 18154
rect 31668 18090 31720 18096
rect 31680 17746 31708 18090
rect 31668 17740 31720 17746
rect 31668 17682 31720 17688
rect 32048 17354 32076 22918
rect 32140 18426 32168 33866
rect 32310 33008 32366 33017
rect 32310 32943 32366 32952
rect 32324 31890 32352 32943
rect 32312 31884 32364 31890
rect 32312 31826 32364 31832
rect 32600 31482 32628 34954
rect 32680 34400 32732 34406
rect 32678 34368 32680 34377
rect 32732 34368 32734 34377
rect 32678 34303 32734 34312
rect 32692 34134 32720 34303
rect 32680 34128 32732 34134
rect 32680 34070 32732 34076
rect 32588 31476 32640 31482
rect 32588 31418 32640 31424
rect 32220 31272 32272 31278
rect 32220 31214 32272 31220
rect 32232 30802 32260 31214
rect 32220 30796 32272 30802
rect 32220 30738 32272 30744
rect 32232 29714 32260 30738
rect 32772 30660 32824 30666
rect 32772 30602 32824 30608
rect 32784 30569 32812 30602
rect 32770 30560 32826 30569
rect 32770 30495 32826 30504
rect 32220 29708 32272 29714
rect 32220 29650 32272 29656
rect 32232 29170 32260 29650
rect 32220 29164 32272 29170
rect 32220 29106 32272 29112
rect 32232 28626 32260 29106
rect 32876 28762 32904 35866
rect 33244 35630 33272 35866
rect 33520 35766 33548 36110
rect 34072 35894 34100 36790
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35256 36100 35308 36106
rect 35256 36042 35308 36048
rect 33980 35866 34100 35894
rect 35268 35894 35296 36042
rect 35268 35866 35388 35894
rect 33508 35760 33560 35766
rect 33508 35702 33560 35708
rect 33232 35624 33284 35630
rect 33232 35566 33284 35572
rect 33244 35154 33272 35566
rect 33232 35148 33284 35154
rect 33232 35090 33284 35096
rect 33244 34746 33272 35090
rect 33324 35012 33376 35018
rect 33324 34954 33376 34960
rect 33232 34740 33284 34746
rect 33232 34682 33284 34688
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 32968 30734 32996 33458
rect 32956 30728 33008 30734
rect 32956 30670 33008 30676
rect 32956 29572 33008 29578
rect 32956 29514 33008 29520
rect 32864 28756 32916 28762
rect 32864 28698 32916 28704
rect 32220 28620 32272 28626
rect 32220 28562 32272 28568
rect 32772 28484 32824 28490
rect 32772 28426 32824 28432
rect 32496 28144 32548 28150
rect 32496 28086 32548 28092
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32312 27328 32364 27334
rect 32312 27270 32364 27276
rect 32324 25242 32352 27270
rect 32232 25214 32352 25242
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 31956 17326 32076 17354
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31576 16176 31628 16182
rect 31576 16118 31628 16124
rect 31666 15600 31722 15609
rect 31864 15570 31892 16458
rect 31666 15535 31722 15544
rect 31852 15564 31904 15570
rect 31680 15502 31708 15535
rect 31852 15506 31904 15512
rect 31956 15502 31984 17326
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31484 12844 31536 12850
rect 31484 12786 31536 12792
rect 31208 12776 31260 12782
rect 31208 12718 31260 12724
rect 31024 12436 31076 12442
rect 31024 12378 31076 12384
rect 31116 12164 31168 12170
rect 31116 12106 31168 12112
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 31128 11354 31156 12106
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 30472 6724 30524 6730
rect 30472 6666 30524 6672
rect 30840 6724 30892 6730
rect 30840 6666 30892 6672
rect 30484 5370 30512 6666
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 27620 2304 27672 2310
rect 27620 2246 27672 2252
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 27724 800 27752 2246
rect 29012 800 29040 2246
rect 30300 800 30328 2790
rect 31220 2514 31248 12718
rect 31576 12640 31628 12646
rect 31576 12582 31628 12588
rect 31392 12368 31444 12374
rect 31392 12310 31444 12316
rect 31404 12170 31432 12310
rect 31392 12164 31444 12170
rect 31392 12106 31444 12112
rect 31588 11830 31616 12582
rect 31576 11824 31628 11830
rect 31576 11766 31628 11772
rect 31668 11824 31720 11830
rect 31668 11766 31720 11772
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31312 11218 31340 11630
rect 31300 11212 31352 11218
rect 31300 11154 31352 11160
rect 31392 7812 31444 7818
rect 31392 7754 31444 7760
rect 31404 2990 31432 7754
rect 31680 6866 31708 11766
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 31680 6202 31708 6802
rect 31588 6174 31708 6202
rect 31588 2990 31616 6174
rect 31668 6112 31720 6118
rect 31668 6054 31720 6060
rect 31392 2984 31444 2990
rect 31392 2926 31444 2932
rect 31576 2984 31628 2990
rect 31576 2926 31628 2932
rect 31208 2508 31260 2514
rect 31208 2450 31260 2456
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 30944 800 30972 2382
rect 31680 2378 31708 6054
rect 32048 2514 32076 17138
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 32140 12918 32168 17070
rect 32232 15094 32260 25214
rect 32312 22092 32364 22098
rect 32312 22034 32364 22040
rect 32324 18970 32352 22034
rect 32312 18964 32364 18970
rect 32312 18906 32364 18912
rect 32416 18630 32444 27406
rect 32508 22982 32536 28086
rect 32680 23860 32732 23866
rect 32680 23802 32732 23808
rect 32692 23526 32720 23802
rect 32588 23520 32640 23526
rect 32588 23462 32640 23468
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32496 22976 32548 22982
rect 32496 22918 32548 22924
rect 32600 20602 32628 23462
rect 32680 21480 32732 21486
rect 32680 21422 32732 21428
rect 32692 20874 32720 21422
rect 32680 20868 32732 20874
rect 32680 20810 32732 20816
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32692 20058 32720 20810
rect 32680 20052 32732 20058
rect 32680 19994 32732 20000
rect 32678 19952 32734 19961
rect 32678 19887 32734 19896
rect 32692 19786 32720 19887
rect 32680 19780 32732 19786
rect 32680 19722 32732 19728
rect 32784 19156 32812 28426
rect 32864 22094 32916 22098
rect 32968 22094 32996 29514
rect 33140 29096 33192 29102
rect 33060 29056 33140 29084
rect 33060 28490 33088 29056
rect 33140 29038 33192 29044
rect 33048 28484 33100 28490
rect 33048 28426 33100 28432
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33152 27554 33180 27950
rect 33152 27538 33272 27554
rect 33152 27532 33284 27538
rect 33152 27526 33232 27532
rect 33048 27056 33100 27062
rect 33048 26998 33100 27004
rect 33060 26518 33088 26998
rect 33152 26926 33180 27526
rect 33232 27474 33284 27480
rect 33140 26920 33192 26926
rect 33140 26862 33192 26868
rect 33048 26512 33100 26518
rect 33048 26454 33100 26460
rect 33060 26217 33088 26454
rect 33336 26217 33364 34954
rect 33416 34944 33468 34950
rect 33416 34886 33468 34892
rect 33428 31414 33456 34886
rect 33980 34746 34008 35866
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 34704 35488 34756 35494
rect 34704 35430 34756 35436
rect 34428 35080 34480 35086
rect 34428 35022 34480 35028
rect 33968 34740 34020 34746
rect 33968 34682 34020 34688
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 33416 31408 33468 31414
rect 33416 31350 33468 31356
rect 33520 26908 33548 31894
rect 33600 31816 33652 31822
rect 33600 31758 33652 31764
rect 33428 26880 33548 26908
rect 33046 26208 33102 26217
rect 33046 26143 33102 26152
rect 33322 26208 33378 26217
rect 33322 26143 33378 26152
rect 33048 24744 33100 24750
rect 33048 24686 33100 24692
rect 33060 24274 33088 24686
rect 33048 24268 33100 24274
rect 33048 24210 33100 24216
rect 33232 24064 33284 24070
rect 33232 24006 33284 24012
rect 33244 23186 33272 24006
rect 33324 23656 33376 23662
rect 33324 23598 33376 23604
rect 33336 23254 33364 23598
rect 33324 23248 33376 23254
rect 33324 23190 33376 23196
rect 33232 23180 33284 23186
rect 33232 23122 33284 23128
rect 33140 22568 33192 22574
rect 32864 22092 32996 22094
rect 32916 22066 32996 22092
rect 33060 22528 33140 22556
rect 32864 22034 32916 22040
rect 33060 21978 33088 22528
rect 33140 22510 33192 22516
rect 33140 22432 33192 22438
rect 33140 22374 33192 22380
rect 33152 22273 33180 22374
rect 33138 22264 33194 22273
rect 33138 22199 33194 22208
rect 32876 21950 33088 21978
rect 32876 21894 32904 21950
rect 32864 21888 32916 21894
rect 32864 21830 32916 21836
rect 32692 19128 32812 19156
rect 32404 18624 32456 18630
rect 32404 18566 32456 18572
rect 32310 17912 32366 17921
rect 32310 17847 32366 17856
rect 32220 15088 32272 15094
rect 32220 15030 32272 15036
rect 32324 15026 32352 17847
rect 32692 16182 32720 19128
rect 32876 18834 32904 21830
rect 33140 21004 33192 21010
rect 33140 20946 33192 20952
rect 33152 20602 33180 20946
rect 33140 20596 33192 20602
rect 33140 20538 33192 20544
rect 33048 20460 33100 20466
rect 33048 20402 33100 20408
rect 32954 19408 33010 19417
rect 32954 19343 33010 19352
rect 32864 18828 32916 18834
rect 32864 18770 32916 18776
rect 32864 18692 32916 18698
rect 32864 18634 32916 18640
rect 32876 18222 32904 18634
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32864 17536 32916 17542
rect 32864 17478 32916 17484
rect 32770 16552 32826 16561
rect 32876 16522 32904 17478
rect 32770 16487 32772 16496
rect 32824 16487 32826 16496
rect 32864 16516 32916 16522
rect 32772 16458 32824 16464
rect 32864 16458 32916 16464
rect 32680 16176 32732 16182
rect 32680 16118 32732 16124
rect 32968 15502 32996 19343
rect 33060 18698 33088 20402
rect 33244 19802 33272 23122
rect 33324 21616 33376 21622
rect 33324 21558 33376 21564
rect 33336 20058 33364 21558
rect 33428 21078 33456 26880
rect 33612 26874 33640 31758
rect 33784 28484 33836 28490
rect 33784 28426 33836 28432
rect 33612 26846 33732 26874
rect 33600 26784 33652 26790
rect 33600 26726 33652 26732
rect 33612 26450 33640 26726
rect 33600 26444 33652 26450
rect 33600 26386 33652 26392
rect 33612 25906 33640 26386
rect 33600 25900 33652 25906
rect 33600 25842 33652 25848
rect 33704 25786 33732 26846
rect 33612 25758 33732 25786
rect 33508 23860 33560 23866
rect 33508 23802 33560 23808
rect 33416 21072 33468 21078
rect 33416 21014 33468 21020
rect 33324 20052 33376 20058
rect 33324 19994 33376 20000
rect 33416 19848 33468 19854
rect 33244 19774 33364 19802
rect 33520 19836 33548 23802
rect 33468 19808 33548 19836
rect 33416 19790 33468 19796
rect 33232 19712 33284 19718
rect 33232 19654 33284 19660
rect 33244 19514 33272 19654
rect 33232 19508 33284 19514
rect 33232 19450 33284 19456
rect 33232 19236 33284 19242
rect 33232 19178 33284 19184
rect 33140 18760 33192 18766
rect 33244 18748 33272 19178
rect 33192 18720 33272 18748
rect 33140 18702 33192 18708
rect 33048 18692 33100 18698
rect 33048 18634 33100 18640
rect 33152 18290 33180 18702
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 33048 18148 33100 18154
rect 33048 18090 33100 18096
rect 33060 16998 33088 18090
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 33048 16040 33100 16046
rect 33048 15982 33100 15988
rect 33060 15638 33088 15982
rect 33048 15632 33100 15638
rect 33048 15574 33100 15580
rect 32772 15496 32824 15502
rect 32772 15438 32824 15444
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32404 15360 32456 15366
rect 32404 15302 32456 15308
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32416 14482 32444 15302
rect 32404 14476 32456 14482
rect 32404 14418 32456 14424
rect 32784 13938 32812 15438
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32772 13932 32824 13938
rect 32772 13874 32824 13880
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32128 12912 32180 12918
rect 32128 12854 32180 12860
rect 32324 12850 32352 13262
rect 32600 12986 32628 13874
rect 32954 13696 33010 13705
rect 32954 13631 33010 13640
rect 32968 13326 32996 13631
rect 33336 13326 33364 19774
rect 33428 17610 33456 19790
rect 33508 18964 33560 18970
rect 33508 18906 33560 18912
rect 33520 17678 33548 18906
rect 33612 18426 33640 25758
rect 33692 23248 33744 23254
rect 33692 23190 33744 23196
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33508 17672 33560 17678
rect 33508 17614 33560 17620
rect 33416 17604 33468 17610
rect 33416 17546 33468 17552
rect 33508 17536 33560 17542
rect 33704 17490 33732 23190
rect 33796 21078 33824 28426
rect 33876 27872 33928 27878
rect 33876 27814 33928 27820
rect 33888 25974 33916 27814
rect 33980 27713 34008 34682
rect 34440 34066 34468 35022
rect 34716 35018 34744 35430
rect 34612 35012 34664 35018
rect 34612 34954 34664 34960
rect 34704 35012 34756 35018
rect 34704 34954 34756 34960
rect 34428 34060 34480 34066
rect 34428 34002 34480 34008
rect 34440 33590 34468 34002
rect 34520 33924 34572 33930
rect 34520 33866 34572 33872
rect 34428 33584 34480 33590
rect 34428 33526 34480 33532
rect 34532 33114 34560 33866
rect 34060 33108 34112 33114
rect 34060 33050 34112 33056
rect 34520 33108 34572 33114
rect 34520 33050 34572 33056
rect 34072 31958 34100 33050
rect 34060 31952 34112 31958
rect 34060 31894 34112 31900
rect 34072 31822 34100 31894
rect 34060 31816 34112 31822
rect 34060 31758 34112 31764
rect 34244 30932 34296 30938
rect 34244 30874 34296 30880
rect 34060 29232 34112 29238
rect 34060 29174 34112 29180
rect 33966 27704 34022 27713
rect 33966 27639 34022 27648
rect 33876 25968 33928 25974
rect 33876 25910 33928 25916
rect 33888 23746 33916 25910
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 33980 23866 34008 24686
rect 33968 23860 34020 23866
rect 33968 23802 34020 23808
rect 33888 23718 34008 23746
rect 33876 23044 33928 23050
rect 33876 22986 33928 22992
rect 33784 21072 33836 21078
rect 33784 21014 33836 21020
rect 33888 19718 33916 22986
rect 33876 19712 33928 19718
rect 33876 19654 33928 19660
rect 33508 17478 33560 17484
rect 33520 17270 33548 17478
rect 33612 17462 33732 17490
rect 33508 17264 33560 17270
rect 33508 17206 33560 17212
rect 32956 13320 33008 13326
rect 32956 13262 33008 13268
rect 33324 13320 33376 13326
rect 33324 13262 33376 13268
rect 32588 12980 32640 12986
rect 32588 12922 32640 12928
rect 33612 12850 33640 17462
rect 33692 15428 33744 15434
rect 33692 15370 33744 15376
rect 33704 14822 33732 15370
rect 33980 14958 34008 23718
rect 34072 21622 34100 29174
rect 34256 28422 34284 30874
rect 34624 30161 34652 34954
rect 34716 33998 34744 34954
rect 34704 33992 34756 33998
rect 34704 33934 34756 33940
rect 34808 31249 34836 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35256 35284 35308 35290
rect 35256 35226 35308 35232
rect 35268 34610 35296 35226
rect 35256 34604 35308 34610
rect 35256 34546 35308 34552
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34794 31240 34850 31249
rect 34794 31175 34850 31184
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30184 34848 30190
rect 34610 30152 34666 30161
rect 35256 30184 35308 30190
rect 34796 30126 34848 30132
rect 35254 30152 35256 30161
rect 35308 30152 35310 30161
rect 34610 30087 34666 30096
rect 34808 29714 34836 30126
rect 35254 30087 35310 30096
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29708 34848 29714
rect 34796 29650 34848 29656
rect 35164 29572 35216 29578
rect 35164 29514 35216 29520
rect 35176 29306 35204 29514
rect 35164 29300 35216 29306
rect 35164 29242 35216 29248
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34244 28416 34296 28422
rect 34244 28358 34296 28364
rect 34256 23497 34284 28358
rect 34796 28144 34848 28150
rect 34796 28086 34848 28092
rect 34612 27668 34664 27674
rect 34612 27610 34664 27616
rect 34428 27464 34480 27470
rect 34428 27406 34480 27412
rect 34440 26790 34468 27406
rect 34624 27130 34652 27610
rect 34612 27124 34664 27130
rect 34612 27066 34664 27072
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34440 26450 34468 26726
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34428 26444 34480 26450
rect 34428 26386 34480 26392
rect 34520 26308 34572 26314
rect 34520 26250 34572 26256
rect 34428 24404 34480 24410
rect 34428 24346 34480 24352
rect 34336 23792 34388 23798
rect 34336 23734 34388 23740
rect 34242 23488 34298 23497
rect 34242 23423 34298 23432
rect 34060 21616 34112 21622
rect 34060 21558 34112 21564
rect 34152 21548 34204 21554
rect 34152 21490 34204 21496
rect 34164 21146 34192 21490
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 34060 20868 34112 20874
rect 34060 20810 34112 20816
rect 34072 20058 34100 20810
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 34244 19712 34296 19718
rect 34244 19654 34296 19660
rect 34058 19544 34114 19553
rect 34058 19479 34114 19488
rect 34072 18970 34100 19479
rect 34256 19446 34284 19654
rect 34348 19514 34376 23734
rect 34440 23610 34468 24346
rect 34532 24206 34560 26250
rect 34716 25362 34744 26522
rect 34704 25356 34756 25362
rect 34704 25298 34756 25304
rect 34612 25288 34664 25294
rect 34612 25230 34664 25236
rect 34624 24274 34652 25230
rect 34612 24268 34664 24274
rect 34612 24210 34664 24216
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34624 23746 34652 24210
rect 34532 23730 34652 23746
rect 34520 23724 34652 23730
rect 34572 23718 34652 23724
rect 34520 23666 34572 23672
rect 34440 23582 34560 23610
rect 34532 22094 34560 23582
rect 34624 23186 34652 23718
rect 34612 23180 34664 23186
rect 34612 23122 34664 23128
rect 34624 22642 34652 23122
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 34716 22234 34744 25298
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 34808 22094 34836 28086
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 25498 35388 35866
rect 35452 29510 35480 39200
rect 36096 37126 36124 39200
rect 36726 38856 36782 38865
rect 36726 38791 36782 38800
rect 36266 37496 36322 37505
rect 36266 37431 36322 37440
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 36084 37120 36136 37126
rect 36084 37062 36136 37068
rect 35900 36576 35952 36582
rect 35900 36518 35952 36524
rect 36084 36576 36136 36582
rect 36084 36518 36136 36524
rect 35912 36378 35940 36518
rect 35900 36372 35952 36378
rect 35900 36314 35952 36320
rect 35532 36032 35584 36038
rect 35532 35974 35584 35980
rect 35544 33590 35572 35974
rect 35624 35760 35676 35766
rect 35624 35702 35676 35708
rect 35636 34649 35664 35702
rect 35716 35624 35768 35630
rect 35716 35566 35768 35572
rect 35728 35290 35756 35566
rect 35716 35284 35768 35290
rect 35716 35226 35768 35232
rect 35854 34672 35906 34678
rect 35622 34640 35678 34649
rect 35622 34575 35678 34584
rect 35728 34620 35854 34626
rect 35728 34614 35906 34620
rect 35728 34598 35894 34614
rect 35728 34202 35756 34598
rect 35716 34196 35768 34202
rect 35716 34138 35768 34144
rect 35900 33924 35952 33930
rect 35900 33866 35952 33872
rect 35532 33584 35584 33590
rect 35532 33526 35584 33532
rect 35912 33538 35940 33866
rect 35912 33510 36032 33538
rect 35900 33448 35952 33454
rect 35900 33390 35952 33396
rect 35912 32026 35940 33390
rect 35900 32020 35952 32026
rect 35900 31962 35952 31968
rect 35532 31884 35584 31890
rect 35532 31826 35584 31832
rect 35544 31754 35572 31826
rect 35544 31726 35664 31754
rect 35532 31136 35584 31142
rect 35532 31078 35584 31084
rect 35440 29504 35492 29510
rect 35440 29446 35492 29452
rect 35544 29322 35572 31078
rect 35452 29294 35572 29322
rect 35452 28966 35480 29294
rect 35440 28960 35492 28966
rect 35440 28902 35492 28908
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 35348 25152 35400 25158
rect 35348 25094 35400 25100
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24290 35388 25094
rect 35268 24274 35388 24290
rect 35256 24268 35388 24274
rect 35308 24262 35388 24268
rect 35452 24290 35480 28902
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35544 25242 35572 27270
rect 35636 26926 35664 31726
rect 35808 31476 35860 31482
rect 35808 31418 35860 31424
rect 35820 31346 35848 31418
rect 35808 31340 35860 31346
rect 35808 31282 35860 31288
rect 35624 26920 35676 26926
rect 35624 26862 35676 26868
rect 35636 25401 35664 26862
rect 35716 25968 35768 25974
rect 35716 25910 35768 25916
rect 35622 25392 35678 25401
rect 35622 25327 35678 25336
rect 35544 25214 35664 25242
rect 35452 24262 35572 24290
rect 35256 24210 35308 24216
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34888 22228 34940 22234
rect 34888 22170 34940 22176
rect 34532 22066 34652 22094
rect 34624 21434 34652 22066
rect 34440 21406 34652 21434
rect 34716 22066 34836 22094
rect 34440 20210 34468 21406
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34532 20534 34560 21286
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34716 20890 34744 22066
rect 34796 21956 34848 21962
rect 34796 21898 34848 21904
rect 34808 21146 34836 21898
rect 34900 21350 34928 22170
rect 34980 21956 35032 21962
rect 34980 21898 35032 21904
rect 35072 21956 35124 21962
rect 35072 21898 35124 21904
rect 34992 21486 35020 21898
rect 35084 21690 35112 21898
rect 35072 21684 35124 21690
rect 35072 21626 35124 21632
rect 34980 21480 35032 21486
rect 34980 21422 35032 21428
rect 34888 21344 34940 21350
rect 34888 21286 34940 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21140 34848 21146
rect 34796 21082 34848 21088
rect 34794 21040 34850 21049
rect 34794 20975 34796 20984
rect 34848 20975 34850 20984
rect 35256 21004 35308 21010
rect 34796 20946 34848 20952
rect 35256 20946 35308 20952
rect 34520 20528 34572 20534
rect 34624 20505 34652 20878
rect 34716 20862 34836 20890
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34520 20470 34572 20476
rect 34610 20496 34666 20505
rect 34610 20431 34666 20440
rect 34610 20360 34666 20369
rect 34610 20295 34666 20304
rect 34440 20182 34560 20210
rect 34428 19984 34480 19990
rect 34428 19926 34480 19932
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 34244 19440 34296 19446
rect 34244 19382 34296 19388
rect 34440 19378 34468 19926
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34060 18964 34112 18970
rect 34060 18906 34112 18912
rect 34164 18766 34192 19314
rect 34152 18760 34204 18766
rect 34152 18702 34204 18708
rect 34164 18290 34192 18702
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 34152 17876 34204 17882
rect 34152 17818 34204 17824
rect 34164 17678 34192 17818
rect 34152 17672 34204 17678
rect 34152 17614 34204 17620
rect 34242 16552 34298 16561
rect 34426 16552 34482 16561
rect 34348 16522 34426 16538
rect 34242 16487 34298 16496
rect 34336 16516 34426 16522
rect 34152 15564 34204 15570
rect 34152 15506 34204 15512
rect 33968 14952 34020 14958
rect 33968 14894 34020 14900
rect 33692 14816 33744 14822
rect 33692 14758 33744 14764
rect 33704 14618 33732 14758
rect 33692 14612 33744 14618
rect 33692 14554 33744 14560
rect 34164 14414 34192 15506
rect 34256 14414 34284 16487
rect 34388 16510 34426 16516
rect 34426 16487 34482 16496
rect 34336 16458 34388 16464
rect 34532 16182 34560 20182
rect 34624 18902 34652 20295
rect 34716 18970 34744 20742
rect 34808 20369 34836 20862
rect 34794 20360 34850 20369
rect 34794 20295 34850 20304
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 35268 20210 35296 20946
rect 35360 20398 35388 24262
rect 35544 22094 35572 24262
rect 35636 23186 35664 25214
rect 35624 23180 35676 23186
rect 35624 23122 35676 23128
rect 35544 22066 35664 22094
rect 35440 21956 35492 21962
rect 35440 21898 35492 21904
rect 35452 21010 35480 21898
rect 35532 21344 35584 21350
rect 35532 21286 35584 21292
rect 35440 21004 35492 21010
rect 35440 20946 35492 20952
rect 35348 20392 35400 20398
rect 35348 20334 35400 20340
rect 35440 20324 35492 20330
rect 35440 20266 35492 20272
rect 34808 19802 34836 20198
rect 35268 20182 35388 20210
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35360 20040 35388 20182
rect 35452 20058 35480 20266
rect 35268 20012 35388 20040
rect 35440 20052 35492 20058
rect 34808 19786 35112 19802
rect 34808 19780 35124 19786
rect 34808 19774 35072 19780
rect 35072 19722 35124 19728
rect 34888 19712 34940 19718
rect 34888 19654 34940 19660
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34612 18896 34664 18902
rect 34808 18850 34836 19450
rect 34900 19417 34928 19654
rect 35268 19514 35296 20012
rect 35440 19994 35492 20000
rect 35544 19938 35572 21286
rect 35360 19910 35572 19938
rect 35256 19508 35308 19514
rect 35256 19450 35308 19456
rect 34886 19408 34942 19417
rect 34886 19343 34942 19352
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35256 18964 35308 18970
rect 35256 18906 35308 18912
rect 35268 18873 35296 18906
rect 34612 18838 34664 18844
rect 34716 18822 34836 18850
rect 35254 18864 35310 18873
rect 34612 18420 34664 18426
rect 34612 18362 34664 18368
rect 34624 18290 34652 18362
rect 34612 18284 34664 18290
rect 34612 18226 34664 18232
rect 34624 17134 34652 18226
rect 34612 17128 34664 17134
rect 34612 17070 34664 17076
rect 34428 16176 34480 16182
rect 34428 16118 34480 16124
rect 34520 16176 34572 16182
rect 34520 16118 34572 16124
rect 34152 14408 34204 14414
rect 34152 14350 34204 14356
rect 34244 14408 34296 14414
rect 34244 14350 34296 14356
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33048 12640 33100 12646
rect 33048 12582 33100 12588
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 32220 12096 32272 12102
rect 32220 12038 32272 12044
rect 32140 11082 32168 12038
rect 32232 11694 32260 12038
rect 32968 11898 32996 12174
rect 32956 11892 33008 11898
rect 32956 11834 33008 11840
rect 32220 11688 32272 11694
rect 32220 11630 32272 11636
rect 33060 11626 33088 12582
rect 33232 12096 33284 12102
rect 33232 12038 33284 12044
rect 33244 11762 33272 12038
rect 34440 11830 34468 16118
rect 34520 15972 34572 15978
rect 34520 15914 34572 15920
rect 34532 15706 34560 15914
rect 34520 15700 34572 15706
rect 34520 15642 34572 15648
rect 34624 15094 34652 17070
rect 34612 15088 34664 15094
rect 34612 15030 34664 15036
rect 34520 14952 34572 14958
rect 34520 14894 34572 14900
rect 34532 14074 34560 14894
rect 34716 14770 34744 18822
rect 35254 18799 35310 18808
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17746 35388 19910
rect 35440 19780 35492 19786
rect 35440 19722 35492 19728
rect 35452 18426 35480 19722
rect 35532 19440 35584 19446
rect 35532 19382 35584 19388
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 35348 17740 35400 17746
rect 35348 17682 35400 17688
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 34808 16794 34836 17614
rect 35348 17536 35400 17542
rect 35348 17478 35400 17484
rect 35360 17270 35388 17478
rect 35348 17264 35400 17270
rect 35348 17206 35400 17212
rect 35348 17128 35400 17134
rect 35348 17070 35400 17076
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 34888 16720 34940 16726
rect 34624 14742 34744 14770
rect 34808 16668 34888 16674
rect 34808 16662 34940 16668
rect 34808 16646 34928 16662
rect 35360 16658 35388 17070
rect 35348 16652 35400 16658
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 34520 13320 34572 13326
rect 34520 13262 34572 13268
rect 34532 12442 34560 13262
rect 34520 12436 34572 12442
rect 34520 12378 34572 12384
rect 34624 12186 34652 14742
rect 34808 13410 34836 16646
rect 35348 16594 35400 16600
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34888 15088 34940 15094
rect 34888 15030 34940 15036
rect 34900 14822 34928 15030
rect 34888 14816 34940 14822
rect 34888 14758 34940 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14482 35388 16594
rect 35544 16454 35572 19382
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35636 16114 35664 22066
rect 35728 21690 35756 25910
rect 35820 24410 35848 31282
rect 35912 30802 35940 31962
rect 35900 30796 35952 30802
rect 35900 30738 35952 30744
rect 35808 24404 35860 24410
rect 35808 24346 35860 24352
rect 35900 24132 35952 24138
rect 35900 24074 35952 24080
rect 35912 23882 35940 24074
rect 35820 23854 35940 23882
rect 35820 23610 35848 23854
rect 35820 23582 35940 23610
rect 35808 23180 35860 23186
rect 35808 23122 35860 23128
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 35716 20052 35768 20058
rect 35716 19994 35768 20000
rect 35728 16726 35756 19994
rect 35716 16720 35768 16726
rect 35716 16662 35768 16668
rect 35624 16108 35676 16114
rect 35624 16050 35676 16056
rect 35820 15892 35848 23122
rect 35912 20602 35940 23582
rect 35900 20596 35952 20602
rect 35900 20538 35952 20544
rect 36004 19514 36032 33510
rect 36096 31822 36124 36518
rect 36188 36378 36216 37198
rect 36176 36372 36228 36378
rect 36176 36314 36228 36320
rect 36280 36310 36308 37431
rect 36740 36854 36768 38791
rect 37384 36922 37412 39200
rect 38672 37330 38700 39200
rect 38660 37324 38712 37330
rect 38660 37266 38712 37272
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 36544 36848 36596 36854
rect 36544 36790 36596 36796
rect 36728 36848 36780 36854
rect 36728 36790 36780 36796
rect 36268 36304 36320 36310
rect 36268 36246 36320 36252
rect 36176 36168 36228 36174
rect 36176 36110 36228 36116
rect 36188 34542 36216 36110
rect 36176 34536 36228 34542
rect 36176 34478 36228 34484
rect 36188 33454 36216 34478
rect 36176 33448 36228 33454
rect 36176 33390 36228 33396
rect 36084 31816 36136 31822
rect 36082 31784 36084 31793
rect 36136 31784 36138 31793
rect 36082 31719 36138 31728
rect 36452 31136 36504 31142
rect 36452 31078 36504 31084
rect 36464 30802 36492 31078
rect 36452 30796 36504 30802
rect 36452 30738 36504 30744
rect 36268 30320 36320 30326
rect 36268 30262 36320 30268
rect 36176 25220 36228 25226
rect 36176 25162 36228 25168
rect 36084 22772 36136 22778
rect 36084 22714 36136 22720
rect 36096 20602 36124 22714
rect 36084 20596 36136 20602
rect 36084 20538 36136 20544
rect 36084 20256 36136 20262
rect 36084 20198 36136 20204
rect 36096 19854 36124 20198
rect 36188 20058 36216 25162
rect 36280 22094 36308 30262
rect 36556 29102 36584 36790
rect 37464 36780 37516 36786
rect 37464 36722 37516 36728
rect 36820 35012 36872 35018
rect 36820 34954 36872 34960
rect 36636 31272 36688 31278
rect 36636 31214 36688 31220
rect 36648 30054 36676 31214
rect 36636 30048 36688 30054
rect 36636 29990 36688 29996
rect 36544 29096 36596 29102
rect 36544 29038 36596 29044
rect 36452 24880 36504 24886
rect 36452 24822 36504 24828
rect 36360 23520 36412 23526
rect 36358 23488 36360 23497
rect 36412 23488 36414 23497
rect 36358 23423 36414 23432
rect 36464 22234 36492 24822
rect 36544 22772 36596 22778
rect 36544 22714 36596 22720
rect 36452 22228 36504 22234
rect 36452 22170 36504 22176
rect 36280 22066 36400 22094
rect 36372 21622 36400 22066
rect 36452 22024 36504 22030
rect 36452 21966 36504 21972
rect 36360 21616 36412 21622
rect 36360 21558 36412 21564
rect 36464 20942 36492 21966
rect 36556 21894 36584 22714
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 36544 21548 36596 21554
rect 36544 21490 36596 21496
rect 36556 20942 36584 21490
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36544 20936 36596 20942
rect 36544 20878 36596 20884
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 36176 20052 36228 20058
rect 36176 19994 36228 20000
rect 36280 19922 36308 20402
rect 36464 19990 36492 20878
rect 36452 19984 36504 19990
rect 36452 19926 36504 19932
rect 36268 19916 36320 19922
rect 36268 19858 36320 19864
rect 36556 19854 36584 20878
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36544 19848 36596 19854
rect 36544 19790 36596 19796
rect 35992 19508 36044 19514
rect 35992 19450 36044 19456
rect 35992 19372 36044 19378
rect 36096 19360 36124 19790
rect 36044 19332 36124 19360
rect 36176 19372 36228 19378
rect 35992 19314 36044 19320
rect 36176 19314 36228 19320
rect 36188 18766 36216 19314
rect 36360 19304 36412 19310
rect 36360 19246 36412 19252
rect 35900 18760 35952 18766
rect 35898 18728 35900 18737
rect 36176 18760 36228 18766
rect 35952 18728 35954 18737
rect 36176 18702 36228 18708
rect 35898 18663 35954 18672
rect 36372 18290 36400 19246
rect 36556 18358 36584 19790
rect 36544 18352 36596 18358
rect 36544 18294 36596 18300
rect 36360 18284 36412 18290
rect 36360 18226 36412 18232
rect 36452 18216 36504 18222
rect 36082 18184 36138 18193
rect 36452 18158 36504 18164
rect 36082 18119 36138 18128
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 35912 17241 35940 17682
rect 35898 17232 35954 17241
rect 35898 17167 35954 17176
rect 36096 17134 36124 18119
rect 36084 17128 36136 17134
rect 36084 17070 36136 17076
rect 36360 17128 36412 17134
rect 36360 17070 36412 17076
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 36004 16250 36032 16526
rect 35992 16244 36044 16250
rect 35992 16186 36044 16192
rect 35452 15864 35848 15892
rect 35348 14476 35400 14482
rect 35348 14418 35400 14424
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34808 13382 35020 13410
rect 34796 13252 34848 13258
rect 34796 13194 34848 13200
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34716 12306 34744 12378
rect 34808 12322 34836 13194
rect 34888 13184 34940 13190
rect 34888 13126 34940 13132
rect 34900 12918 34928 13126
rect 34992 12918 35020 13382
rect 35348 13388 35400 13394
rect 35348 13330 35400 13336
rect 34888 12912 34940 12918
rect 34888 12854 34940 12860
rect 34980 12912 35032 12918
rect 34980 12854 35032 12860
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12442 35388 13330
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 34704 12300 34756 12306
rect 34808 12294 35112 12322
rect 34704 12242 34756 12248
rect 34532 12158 34652 12186
rect 35084 12170 35112 12294
rect 35072 12164 35124 12170
rect 34532 11898 34560 12158
rect 35072 12106 35124 12112
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 34428 11824 34480 11830
rect 34428 11766 34480 11772
rect 33232 11756 33284 11762
rect 33232 11698 33284 11704
rect 34624 11694 34652 12038
rect 35452 11762 35480 15864
rect 35624 15700 35676 15706
rect 35624 15642 35676 15648
rect 35636 14890 35664 15642
rect 35900 15496 35952 15502
rect 35900 15438 35952 15444
rect 35912 15162 35940 15438
rect 36372 15434 36400 17070
rect 36360 15428 36412 15434
rect 36360 15370 36412 15376
rect 36372 15314 36400 15370
rect 36004 15286 36400 15314
rect 35900 15156 35952 15162
rect 35900 15098 35952 15104
rect 35624 14884 35676 14890
rect 35624 14826 35676 14832
rect 35808 14816 35860 14822
rect 35808 14758 35860 14764
rect 35900 14816 35952 14822
rect 35900 14758 35952 14764
rect 35624 14340 35676 14346
rect 35624 14282 35676 14288
rect 35636 13258 35664 14282
rect 35820 14090 35848 14758
rect 35912 14414 35940 14758
rect 35900 14408 35952 14414
rect 35900 14350 35952 14356
rect 35820 14062 35940 14090
rect 35808 14000 35860 14006
rect 35808 13942 35860 13948
rect 35716 13864 35768 13870
rect 35716 13806 35768 13812
rect 35624 13252 35676 13258
rect 35624 13194 35676 13200
rect 35532 13184 35584 13190
rect 35532 13126 35584 13132
rect 35544 12782 35572 13126
rect 35624 12912 35676 12918
rect 35624 12854 35676 12860
rect 35532 12776 35584 12782
rect 35532 12718 35584 12724
rect 35636 12306 35664 12854
rect 35624 12300 35676 12306
rect 35624 12242 35676 12248
rect 35728 11898 35756 13806
rect 35820 13530 35848 13942
rect 35912 13870 35940 14062
rect 35900 13864 35952 13870
rect 35900 13806 35952 13812
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35912 13410 35940 13806
rect 35820 13382 35940 13410
rect 35820 12782 35848 13382
rect 35808 12776 35860 12782
rect 35808 12718 35860 12724
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35440 11756 35492 11762
rect 35440 11698 35492 11704
rect 34612 11688 34664 11694
rect 34612 11630 34664 11636
rect 33048 11620 33100 11626
rect 33048 11562 33100 11568
rect 34796 11620 34848 11626
rect 34796 11562 34848 11568
rect 32404 11552 32456 11558
rect 32404 11494 32456 11500
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 32416 8974 32444 11494
rect 34808 11150 34836 11562
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 35452 10742 35480 11698
rect 36004 11354 36032 15286
rect 36464 14414 36492 18158
rect 36648 15570 36676 29990
rect 36728 23656 36780 23662
rect 36728 23598 36780 23604
rect 36740 22778 36768 23598
rect 36728 22772 36780 22778
rect 36728 22714 36780 22720
rect 36726 20088 36782 20097
rect 36726 20023 36728 20032
rect 36780 20023 36782 20032
rect 36728 19994 36780 20000
rect 36832 19514 36860 34954
rect 37476 32994 37504 36722
rect 37832 36168 37884 36174
rect 37832 36110 37884 36116
rect 38198 36136 38254 36145
rect 37740 36100 37792 36106
rect 37740 36042 37792 36048
rect 37556 35488 37608 35494
rect 37556 35430 37608 35436
rect 37568 35086 37596 35430
rect 37556 35080 37608 35086
rect 37556 35022 37608 35028
rect 37476 32966 37596 32994
rect 37464 32904 37516 32910
rect 37464 32846 37516 32852
rect 37280 32836 37332 32842
rect 37280 32778 37332 32784
rect 37292 30802 37320 32778
rect 37476 32745 37504 32846
rect 37462 32736 37518 32745
rect 37462 32671 37518 32680
rect 37372 31408 37424 31414
rect 37372 31350 37424 31356
rect 37280 30796 37332 30802
rect 37280 30738 37332 30744
rect 36912 29572 36964 29578
rect 36912 29514 36964 29520
rect 36924 27674 36952 29514
rect 37004 29504 37056 29510
rect 37004 29446 37056 29452
rect 36912 27668 36964 27674
rect 36912 27610 36964 27616
rect 36912 21888 36964 21894
rect 36912 21830 36964 21836
rect 36820 19508 36872 19514
rect 36820 19450 36872 19456
rect 36728 16108 36780 16114
rect 36728 16050 36780 16056
rect 36636 15564 36688 15570
rect 36636 15506 36688 15512
rect 36740 14482 36768 16050
rect 36924 14822 36952 21830
rect 37016 18426 37044 29446
rect 37280 27532 37332 27538
rect 37280 27474 37332 27480
rect 37096 25288 37148 25294
rect 37096 25230 37148 25236
rect 37108 21554 37136 25230
rect 37188 22024 37240 22030
rect 37188 21966 37240 21972
rect 37200 21554 37228 21966
rect 37096 21548 37148 21554
rect 37096 21490 37148 21496
rect 37188 21548 37240 21554
rect 37188 21490 37240 21496
rect 37292 20602 37320 27474
rect 37384 21146 37412 31350
rect 37568 30122 37596 32966
rect 37556 30116 37608 30122
rect 37556 30058 37608 30064
rect 37648 26376 37700 26382
rect 37648 26318 37700 26324
rect 37660 25922 37688 26318
rect 37752 26042 37780 36042
rect 37740 26036 37792 26042
rect 37740 25978 37792 25984
rect 37660 25894 37780 25922
rect 37464 23792 37516 23798
rect 37464 23734 37516 23740
rect 37476 22098 37504 23734
rect 37556 22704 37608 22710
rect 37556 22646 37608 22652
rect 37464 22092 37516 22098
rect 37464 22034 37516 22040
rect 37568 21690 37596 22646
rect 37648 22636 37700 22642
rect 37648 22578 37700 22584
rect 37556 21684 37608 21690
rect 37556 21626 37608 21632
rect 37372 21140 37424 21146
rect 37372 21082 37424 21088
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37200 19854 37228 20402
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37200 19378 37228 19790
rect 37278 19680 37334 19689
rect 37278 19615 37334 19624
rect 37188 19372 37240 19378
rect 37188 19314 37240 19320
rect 37292 18698 37320 19615
rect 37280 18692 37332 18698
rect 37280 18634 37332 18640
rect 37372 18692 37424 18698
rect 37372 18634 37424 18640
rect 37004 18420 37056 18426
rect 37004 18362 37056 18368
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 37200 17678 37228 18226
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37004 16584 37056 16590
rect 37004 16526 37056 16532
rect 37016 15026 37044 16526
rect 37384 16182 37412 18634
rect 37476 17270 37504 19790
rect 37556 18896 37608 18902
rect 37556 18838 37608 18844
rect 37568 18193 37596 18838
rect 37554 18184 37610 18193
rect 37554 18119 37610 18128
rect 37464 17264 37516 17270
rect 37464 17206 37516 17212
rect 37660 16454 37688 22578
rect 37752 20602 37780 25894
rect 37844 23322 37872 36110
rect 38198 36071 38254 36080
rect 38212 36038 38240 36071
rect 38200 36032 38252 36038
rect 38200 35974 38252 35980
rect 38384 35692 38436 35698
rect 38384 35634 38436 35640
rect 38200 35488 38252 35494
rect 38198 35456 38200 35465
rect 38252 35456 38254 35465
rect 38198 35391 38254 35400
rect 37924 34604 37976 34610
rect 37924 34546 37976 34552
rect 37832 23316 37884 23322
rect 37832 23258 37884 23264
rect 37832 23044 37884 23050
rect 37832 22986 37884 22992
rect 37740 20596 37792 20602
rect 37740 20538 37792 20544
rect 37740 18828 37792 18834
rect 37740 18770 37792 18776
rect 37752 18306 37780 18770
rect 37844 18426 37872 22986
rect 37936 20058 37964 34546
rect 38200 34400 38252 34406
rect 38200 34342 38252 34348
rect 38212 34105 38240 34342
rect 38198 34096 38254 34105
rect 38198 34031 38254 34040
rect 38108 33380 38160 33386
rect 38108 33322 38160 33328
rect 38120 32570 38148 33322
rect 38108 32564 38160 32570
rect 38108 32506 38160 32512
rect 38292 32428 38344 32434
rect 38292 32370 38344 32376
rect 38304 32065 38332 32370
rect 38290 32056 38346 32065
rect 38290 31991 38346 32000
rect 38290 30696 38346 30705
rect 38290 30631 38346 30640
rect 38304 30258 38332 30631
rect 38292 30252 38344 30258
rect 38292 30194 38344 30200
rect 38108 29572 38160 29578
rect 38108 29514 38160 29520
rect 38120 29345 38148 29514
rect 38200 29504 38252 29510
rect 38200 29446 38252 29452
rect 38106 29336 38162 29345
rect 38106 29271 38162 29280
rect 38108 29028 38160 29034
rect 38108 28970 38160 28976
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 38028 24954 38056 25230
rect 38016 24948 38068 24954
rect 38016 24890 38068 24896
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 37924 20052 37976 20058
rect 37924 19994 37976 20000
rect 37924 18624 37976 18630
rect 37924 18566 37976 18572
rect 37832 18420 37884 18426
rect 37832 18362 37884 18368
rect 37752 18290 37872 18306
rect 37752 18284 37884 18290
rect 37752 18278 37832 18284
rect 37832 18226 37884 18232
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 37648 16448 37700 16454
rect 37648 16390 37700 16396
rect 37372 16176 37424 16182
rect 37372 16118 37424 16124
rect 37648 15972 37700 15978
rect 37648 15914 37700 15920
rect 37096 15904 37148 15910
rect 37096 15846 37148 15852
rect 37004 15020 37056 15026
rect 37004 14962 37056 14968
rect 36912 14816 36964 14822
rect 36912 14758 36964 14764
rect 36912 14612 36964 14618
rect 36912 14554 36964 14560
rect 36728 14476 36780 14482
rect 36728 14418 36780 14424
rect 36452 14408 36504 14414
rect 36452 14350 36504 14356
rect 36360 13932 36412 13938
rect 36360 13874 36412 13880
rect 36176 13184 36228 13190
rect 36176 13126 36228 13132
rect 36188 12918 36216 13126
rect 36176 12912 36228 12918
rect 36176 12854 36228 12860
rect 36176 12640 36228 12646
rect 36176 12582 36228 12588
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 35440 10736 35492 10742
rect 35440 10678 35492 10684
rect 36188 10674 36216 12582
rect 36372 10810 36400 13874
rect 36818 12336 36874 12345
rect 36818 12271 36874 12280
rect 36452 11756 36504 11762
rect 36452 11698 36504 11704
rect 36360 10804 36412 10810
rect 36360 10746 36412 10752
rect 36176 10668 36228 10674
rect 36176 10610 36228 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 33600 8832 33652 8838
rect 33600 8774 33652 8780
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32416 7886 32444 8026
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32036 2508 32088 2514
rect 32036 2450 32088 2456
rect 33612 2446 33640 8774
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34336 7744 34388 7750
rect 34336 7686 34388 7692
rect 34348 2514 34376 7686
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34336 2508 34388 2514
rect 34336 2450 34388 2456
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 31668 2372 31720 2378
rect 31668 2314 31720 2320
rect 32232 800 32260 2382
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 33520 800 33548 2246
rect 34164 800 34192 2246
rect 35452 800 35480 2994
rect 35912 2446 35940 3878
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36004 3058 36032 3402
rect 36464 3194 36492 11698
rect 36832 11150 36860 12271
rect 36820 11144 36872 11150
rect 36820 11086 36872 11092
rect 36728 11076 36780 11082
rect 36728 11018 36780 11024
rect 36740 4622 36768 11018
rect 36924 10062 36952 14554
rect 37108 13258 37136 15846
rect 37556 15564 37608 15570
rect 37556 15506 37608 15512
rect 37280 14340 37332 14346
rect 37280 14282 37332 14288
rect 37004 13252 37056 13258
rect 37004 13194 37056 13200
rect 37096 13252 37148 13258
rect 37096 13194 37148 13200
rect 37016 12442 37044 13194
rect 37004 12436 37056 12442
rect 37004 12378 37056 12384
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 37292 9450 37320 14282
rect 37568 13462 37596 15506
rect 37660 15434 37688 15914
rect 37648 15428 37700 15434
rect 37648 15370 37700 15376
rect 37752 15366 37780 17682
rect 37844 17678 37872 18226
rect 37832 17672 37884 17678
rect 37832 17614 37884 17620
rect 37936 16590 37964 18566
rect 38028 18154 38056 21966
rect 38016 18148 38068 18154
rect 38016 18090 38068 18096
rect 38120 16726 38148 28970
rect 38212 26897 38240 29446
rect 38292 29164 38344 29170
rect 38292 29106 38344 29112
rect 38304 28665 38332 29106
rect 38290 28656 38346 28665
rect 38290 28591 38346 28600
rect 38292 27464 38344 27470
rect 38292 27406 38344 27412
rect 38304 27305 38332 27406
rect 38290 27296 38346 27305
rect 38290 27231 38346 27240
rect 38198 26888 38254 26897
rect 38198 26823 38254 26832
rect 38292 26376 38344 26382
rect 38292 26318 38344 26324
rect 38304 25945 38332 26318
rect 38290 25936 38346 25945
rect 38290 25871 38346 25880
rect 38198 25256 38254 25265
rect 38198 25191 38254 25200
rect 38212 25158 38240 25191
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38292 24200 38344 24206
rect 38292 24142 38344 24148
rect 38200 24064 38252 24070
rect 38200 24006 38252 24012
rect 38212 23118 38240 24006
rect 38304 23905 38332 24142
rect 38290 23896 38346 23905
rect 38290 23831 38346 23840
rect 38200 23112 38252 23118
rect 38200 23054 38252 23060
rect 38198 22536 38254 22545
rect 38198 22471 38200 22480
rect 38252 22471 38254 22480
rect 38200 22442 38252 22448
rect 38200 21888 38252 21894
rect 38198 21856 38200 21865
rect 38252 21856 38254 21865
rect 38198 21791 38254 21800
rect 38200 19168 38252 19174
rect 38198 19136 38200 19145
rect 38252 19136 38254 19145
rect 38198 19071 38254 19080
rect 38198 17096 38254 17105
rect 38198 17031 38200 17040
rect 38252 17031 38254 17040
rect 38200 17002 38252 17008
rect 38108 16720 38160 16726
rect 38108 16662 38160 16668
rect 37924 16584 37976 16590
rect 37924 16526 37976 16532
rect 38016 16108 38068 16114
rect 38016 16050 38068 16056
rect 37740 15360 37792 15366
rect 37740 15302 37792 15308
rect 37648 14544 37700 14550
rect 37648 14486 37700 14492
rect 37556 13456 37608 13462
rect 37556 13398 37608 13404
rect 37372 12844 37424 12850
rect 37372 12786 37424 12792
rect 37384 10266 37412 12786
rect 37568 11762 37596 13398
rect 37556 11756 37608 11762
rect 37556 11698 37608 11704
rect 37568 11218 37596 11698
rect 37556 11212 37608 11218
rect 37556 11154 37608 11160
rect 37660 11082 37688 14486
rect 38028 14278 38056 16050
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 15745 38240 15846
rect 38198 15736 38254 15745
rect 38198 15671 38254 15680
rect 38106 15056 38162 15065
rect 38106 14991 38108 15000
rect 38160 14991 38162 15000
rect 38108 14962 38160 14968
rect 38016 14272 38068 14278
rect 38016 14214 38068 14220
rect 38200 13728 38252 13734
rect 38198 13696 38200 13705
rect 38252 13696 38254 13705
rect 38198 13631 38254 13640
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 38212 12345 38240 12582
rect 38198 12336 38254 12345
rect 38198 12271 38254 12280
rect 37740 12164 37792 12170
rect 37740 12106 37792 12112
rect 37556 11076 37608 11082
rect 37556 11018 37608 11024
rect 37648 11076 37700 11082
rect 37648 11018 37700 11024
rect 37372 10260 37424 10266
rect 37372 10202 37424 10208
rect 37280 9444 37332 9450
rect 37280 9386 37332 9392
rect 37568 9042 37596 11018
rect 37556 9036 37608 9042
rect 37556 8978 37608 8984
rect 37464 7880 37516 7886
rect 37464 7822 37516 7828
rect 37476 7585 37504 7822
rect 37462 7576 37518 7585
rect 37752 7546 37780 12106
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 10062 37872 11494
rect 38016 11280 38068 11286
rect 38016 11222 38068 11228
rect 38028 10674 38056 11222
rect 38198 10976 38254 10985
rect 38198 10911 38254 10920
rect 38212 10810 38240 10911
rect 38200 10804 38252 10810
rect 38200 10746 38252 10752
rect 38016 10668 38068 10674
rect 38016 10610 38068 10616
rect 38108 10600 38160 10606
rect 38108 10542 38160 10548
rect 37924 10464 37976 10470
rect 37924 10406 37976 10412
rect 37832 10056 37884 10062
rect 37832 9998 37884 10004
rect 37936 9586 37964 10406
rect 37924 9580 37976 9586
rect 37924 9522 37976 9528
rect 38120 8634 38148 10542
rect 38198 10296 38254 10305
rect 38198 10231 38200 10240
rect 38252 10231 38254 10240
rect 38200 10202 38252 10208
rect 38290 8936 38346 8945
rect 38290 8871 38346 8880
rect 38108 8628 38160 8634
rect 38108 8570 38160 8576
rect 38304 8498 38332 8871
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38396 8022 38424 35634
rect 39316 35290 39344 39200
rect 39304 35284 39356 35290
rect 39304 35226 39356 35232
rect 38844 34740 38896 34746
rect 38844 34682 38896 34688
rect 38752 32904 38804 32910
rect 38752 32846 38804 32852
rect 38476 30048 38528 30054
rect 38476 29990 38528 29996
rect 38488 18222 38516 29990
rect 38568 27056 38620 27062
rect 38568 26998 38620 27004
rect 38476 18216 38528 18222
rect 38476 18158 38528 18164
rect 38580 17882 38608 26998
rect 38660 25900 38712 25906
rect 38660 25842 38712 25848
rect 38568 17876 38620 17882
rect 38568 17818 38620 17824
rect 38672 13530 38700 25842
rect 38764 16522 38792 32846
rect 38856 18970 38884 34682
rect 39212 29096 39264 29102
rect 39212 29038 39264 29044
rect 39028 23112 39080 23118
rect 39028 23054 39080 23060
rect 38844 18964 38896 18970
rect 38844 18906 38896 18912
rect 38752 16516 38804 16522
rect 38752 16458 38804 16464
rect 38660 13524 38712 13530
rect 38660 13466 38712 13472
rect 39040 12238 39068 23054
rect 39224 19990 39252 29038
rect 39580 27396 39632 27402
rect 39580 27338 39632 27344
rect 39304 27328 39356 27334
rect 39304 27270 39356 27276
rect 39212 19984 39264 19990
rect 39212 19926 39264 19932
rect 39316 16658 39344 27270
rect 39396 26512 39448 26518
rect 39396 26454 39448 26460
rect 39408 16794 39436 26454
rect 39592 17814 39620 27338
rect 39580 17808 39632 17814
rect 39580 17750 39632 17756
rect 39396 16788 39448 16794
rect 39396 16730 39448 16736
rect 39304 16652 39356 16658
rect 39304 16594 39356 16600
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 38384 8016 38436 8022
rect 38384 7958 38436 7964
rect 37462 7511 37518 7520
rect 37740 7540 37792 7546
rect 37740 7482 37792 7488
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38304 6905 38332 7346
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38200 5568 38252 5574
rect 38198 5536 38200 5545
rect 38252 5536 38254 5545
rect 38198 5471 38254 5480
rect 37740 5160 37792 5166
rect 37740 5102 37792 5108
rect 37752 4690 37780 5102
rect 37740 4684 37792 4690
rect 37740 4626 37792 4632
rect 36728 4616 36780 4622
rect 36728 4558 36780 4564
rect 37464 4616 37516 4622
rect 37464 4558 37516 4564
rect 37476 4185 37504 4558
rect 37462 4176 37518 4185
rect 36728 4140 36780 4146
rect 37462 4111 37518 4120
rect 36728 4082 36780 4088
rect 36740 3738 36768 4082
rect 36728 3732 36780 3738
rect 36728 3674 36780 3680
rect 37740 3596 37792 3602
rect 37740 3538 37792 3544
rect 36452 3188 36504 3194
rect 36452 3130 36504 3136
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 37188 2372 37240 2378
rect 37188 2314 37240 2320
rect 36820 2304 36872 2310
rect 36820 2246 36872 2252
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 36832 2145 36860 2246
rect 36818 2136 36874 2145
rect 36818 2071 36874 2080
rect 36740 870 36860 898
rect 36740 800 36768 870
rect 2870 776 2926 785
rect 2870 711 2926 720
rect 3238 200 3294 800
rect 3882 200 3938 800
rect 5170 200 5226 800
rect 6458 200 6514 800
rect 7102 200 7158 800
rect 8390 200 8446 800
rect 9678 200 9734 800
rect 10322 200 10378 800
rect 11610 200 11666 800
rect 12898 200 12954 800
rect 13542 200 13598 800
rect 14830 200 14886 800
rect 16118 200 16174 800
rect 16762 200 16818 800
rect 18050 200 18106 800
rect 19338 200 19394 800
rect 19982 200 20038 800
rect 21270 200 21326 800
rect 22558 200 22614 800
rect 23202 200 23258 800
rect 24490 200 24546 800
rect 25778 200 25834 800
rect 27066 200 27122 800
rect 27710 200 27766 800
rect 28998 200 29054 800
rect 30286 200 30342 800
rect 30930 200 30986 800
rect 32218 200 32274 800
rect 33506 200 33562 800
rect 34150 200 34206 800
rect 35438 200 35494 800
rect 36726 200 36782 800
rect 36832 762 36860 870
rect 37108 762 37136 2246
rect 36832 734 37136 762
rect 37200 105 37228 2314
rect 37384 800 37412 2994
rect 37370 200 37426 800
rect 37752 785 37780 3538
rect 38198 3496 38254 3505
rect 38198 3431 38254 3440
rect 38212 3398 38240 3431
rect 38200 3392 38252 3398
rect 38200 3334 38252 3340
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 38672 800 38700 2790
rect 37738 776 37794 785
rect 37738 711 37794 720
rect 38658 200 38714 800
rect 37186 96 37242 105
rect 37186 31 37242 40
<< via2 >>
rect 3422 39480 3478 39536
rect 1582 36236 1638 36272
rect 1582 36216 1584 36236
rect 1584 36216 1636 36236
rect 1636 36216 1638 36236
rect 1398 36080 1454 36136
rect 1766 34040 1822 34096
rect 2870 38800 2926 38856
rect 2870 37440 2926 37496
rect 2318 35536 2374 35592
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 3054 35708 3056 35728
rect 3056 35708 3108 35728
rect 3108 35708 3110 35728
rect 3054 35672 3110 35708
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 1766 32716 1768 32736
rect 1768 32716 1820 32736
rect 1820 32716 1822 32736
rect 1766 32680 1822 32716
rect 1766 32000 1822 32056
rect 1766 30640 1822 30696
rect 1766 29280 1822 29336
rect 1582 28600 1638 28656
rect 1674 27240 1730 27296
rect 1766 25880 1822 25936
rect 1766 24556 1768 24576
rect 1768 24556 1820 24576
rect 1820 24556 1822 24576
rect 1766 24520 1822 24556
rect 1582 23840 1638 23896
rect 1766 22480 1822 22536
rect 1674 21120 1730 21176
rect 1674 20440 1730 20496
rect 1766 19080 1822 19136
rect 1582 17720 1638 17776
rect 1766 17040 1822 17096
rect 1766 15680 1822 15736
rect 1766 14356 1768 14376
rect 1768 14356 1820 14376
rect 1820 14356 1822 14376
rect 1766 14320 1822 14356
rect 1766 13676 1768 13696
rect 1768 13676 1820 13696
rect 1820 13676 1822 13696
rect 1766 13640 1822 13676
rect 1766 12280 1822 12336
rect 1674 10920 1730 10976
rect 1766 10240 1822 10296
rect 1766 8880 1822 8936
rect 1766 7520 1822 7576
rect 1766 6840 1822 6896
rect 1766 5480 1822 5536
rect 1766 4120 1822 4176
rect 1766 3440 1822 3496
rect 2318 33904 2374 33960
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 2778 2080 2834 2136
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 6458 35128 6514 35184
rect 8022 36644 8078 36680
rect 8022 36624 8024 36644
rect 8024 36624 8076 36644
rect 8076 36624 8078 36644
rect 6734 36116 6736 36136
rect 6736 36116 6788 36136
rect 6788 36116 6790 36136
rect 6734 36080 6790 36116
rect 8206 33768 8262 33824
rect 9402 33904 9458 33960
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 9678 36780 9734 36816
rect 9678 36760 9680 36780
rect 9680 36760 9732 36780
rect 9732 36760 9734 36780
rect 10598 36780 10654 36816
rect 10598 36760 10600 36780
rect 10600 36760 10652 36780
rect 10652 36760 10654 36780
rect 10046 36352 10102 36408
rect 9770 32680 9826 32736
rect 10138 35436 10140 35456
rect 10140 35436 10192 35456
rect 10192 35436 10194 35456
rect 10138 35400 10194 35436
rect 10506 35264 10562 35320
rect 10230 32952 10286 33008
rect 10782 35828 10838 35864
rect 10782 35808 10784 35828
rect 10784 35808 10836 35828
rect 10836 35808 10838 35828
rect 9770 20848 9826 20904
rect 10966 34740 11022 34776
rect 10966 34720 10968 34740
rect 10968 34720 11020 34740
rect 11020 34720 11022 34740
rect 11518 35944 11574 36000
rect 10966 33496 11022 33552
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11426 30368 11482 30424
rect 10966 23740 10968 23760
rect 10968 23740 11020 23760
rect 11020 23740 11022 23760
rect 10966 23704 11022 23740
rect 10966 20984 11022 21040
rect 11242 21256 11298 21312
rect 11794 35808 11850 35864
rect 11978 35808 12034 35864
rect 12070 33632 12126 33688
rect 11702 32272 11758 32328
rect 12346 32408 12402 32464
rect 11794 21256 11850 21312
rect 12254 21836 12256 21856
rect 12256 21836 12308 21856
rect 12308 21836 12310 21856
rect 12254 21800 12310 21836
rect 12254 21528 12310 21584
rect 13818 35944 13874 36000
rect 14278 35944 14334 36000
rect 13542 35400 13598 35456
rect 12898 33224 12954 33280
rect 12806 32408 12862 32464
rect 12990 32544 13046 32600
rect 13082 27956 13084 27976
rect 13084 27956 13136 27976
rect 13136 27956 13138 27976
rect 13082 27920 13138 27956
rect 12530 21836 12532 21856
rect 12532 21836 12584 21856
rect 12584 21836 12586 21856
rect 12530 21800 12586 21836
rect 12530 21392 12586 21448
rect 13726 21528 13782 21584
rect 13266 17720 13322 17776
rect 14186 34604 14242 34640
rect 14186 34584 14188 34604
rect 14188 34584 14240 34604
rect 14240 34584 14242 34604
rect 14370 30252 14426 30288
rect 14370 30232 14372 30252
rect 14372 30232 14424 30252
rect 14424 30232 14426 30252
rect 14278 20848 14334 20904
rect 15934 37188 15990 37224
rect 15934 37168 15936 37188
rect 15936 37168 15988 37188
rect 15988 37168 15990 37188
rect 18878 37188 18934 37224
rect 18878 37168 18880 37188
rect 18880 37168 18932 37188
rect 18932 37168 18934 37188
rect 15290 34720 15346 34776
rect 15198 32272 15254 32328
rect 15474 33088 15530 33144
rect 14646 20984 14702 21040
rect 16854 36760 16910 36816
rect 16210 36352 16266 36408
rect 17682 36352 17738 36408
rect 16946 35944 17002 36000
rect 15750 34584 15806 34640
rect 15934 33924 15990 33960
rect 15934 33904 15936 33924
rect 15936 33904 15988 33924
rect 15988 33904 15990 33924
rect 17130 35572 17132 35592
rect 17132 35572 17184 35592
rect 17184 35572 17186 35592
rect 16302 33088 16358 33144
rect 16946 32852 16948 32872
rect 16948 32852 17000 32872
rect 17000 32852 17002 32872
rect 16946 32816 17002 32852
rect 15474 30232 15530 30288
rect 15290 23568 15346 23624
rect 15382 21004 15438 21040
rect 15382 20984 15384 21004
rect 15384 20984 15436 21004
rect 15436 20984 15438 21004
rect 15842 21428 15844 21448
rect 15844 21428 15896 21448
rect 15896 21428 15898 21448
rect 15842 21392 15898 21428
rect 17130 35536 17186 35572
rect 17130 33804 17132 33824
rect 17132 33804 17184 33824
rect 17184 33804 17186 33824
rect 17130 33768 17186 33804
rect 17406 35264 17462 35320
rect 17498 32816 17554 32872
rect 17222 21256 17278 21312
rect 17774 35536 17830 35592
rect 17774 33396 17776 33416
rect 17776 33396 17828 33416
rect 17828 33396 17830 33416
rect 17774 33360 17830 33396
rect 18418 35808 18474 35864
rect 17958 35128 18014 35184
rect 18418 33088 18474 33144
rect 18050 32544 18106 32600
rect 18602 23568 18658 23624
rect 18602 23432 18658 23488
rect 18694 21528 18750 21584
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19430 33632 19486 33688
rect 19430 33088 19486 33144
rect 19246 32680 19302 32736
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 20350 35028 20352 35048
rect 20352 35028 20404 35048
rect 20404 35028 20406 35048
rect 20350 34992 20406 35028
rect 20902 35672 20958 35728
rect 20902 33360 20958 33416
rect 22098 35944 22154 36000
rect 21178 33924 21234 33960
rect 21178 33904 21180 33924
rect 21180 33904 21232 33924
rect 21232 33904 21234 33924
rect 21546 33088 21602 33144
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 21454 26288 21510 26344
rect 21546 24792 21602 24848
rect 21178 21140 21234 21176
rect 21178 21120 21180 21140
rect 21180 21120 21232 21140
rect 21232 21120 21234 21140
rect 21270 20984 21326 21040
rect 21362 20884 21364 20904
rect 21364 20884 21416 20904
rect 21416 20884 21418 20904
rect 21362 20848 21418 20884
rect 21270 19080 21326 19136
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 23478 36624 23534 36680
rect 22926 35028 22928 35048
rect 22928 35028 22980 35048
rect 22980 35028 22982 35048
rect 22926 34992 22982 35028
rect 22006 13504 22062 13560
rect 23846 23432 23902 23488
rect 23018 17856 23074 17912
rect 23294 15428 23350 15464
rect 23294 15408 23296 15428
rect 23296 15408 23348 15428
rect 23348 15408 23350 15428
rect 23662 15136 23718 15192
rect 22282 9832 22338 9888
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 24214 18400 24270 18456
rect 24490 24792 24546 24848
rect 28078 37204 28080 37224
rect 28080 37204 28132 37224
rect 28132 37204 28134 37224
rect 28078 37168 28134 37204
rect 26146 36488 26202 36544
rect 26054 36080 26110 36136
rect 26422 36216 26478 36272
rect 26238 35944 26294 36000
rect 27710 36116 27712 36136
rect 27712 36116 27764 36136
rect 27764 36116 27766 36136
rect 27710 36080 27766 36116
rect 26238 34448 26294 34504
rect 26238 33496 26294 33552
rect 25962 27668 26018 27704
rect 25962 27648 25964 27668
rect 25964 27648 26016 27668
rect 26016 27648 26018 27668
rect 25318 20576 25374 20632
rect 25778 20868 25834 20904
rect 25778 20848 25780 20868
rect 25780 20848 25832 20868
rect 25832 20848 25834 20868
rect 25686 20304 25742 20360
rect 26054 18420 26110 18456
rect 26054 18400 26056 18420
rect 26056 18400 26108 18420
rect 26108 18400 26110 18420
rect 26330 19116 26332 19136
rect 26332 19116 26384 19136
rect 26384 19116 26386 19136
rect 26330 19080 26386 19116
rect 26330 18964 26386 19000
rect 26330 18944 26332 18964
rect 26332 18944 26384 18964
rect 26384 18944 26386 18964
rect 27434 26288 27490 26344
rect 27342 23296 27398 23352
rect 27986 36236 28042 36272
rect 27986 36216 27988 36236
rect 27988 36216 28040 36236
rect 28040 36216 28042 36236
rect 28814 36488 28870 36544
rect 28446 36236 28502 36272
rect 28446 36216 28448 36236
rect 28448 36216 28500 36236
rect 28500 36216 28502 36236
rect 31298 37204 31300 37224
rect 31300 37204 31352 37224
rect 31352 37204 31354 37224
rect 31298 37168 31354 37204
rect 28630 36080 28686 36136
rect 28354 35980 28356 36000
rect 28356 35980 28408 36000
rect 28408 35980 28410 36000
rect 28354 35944 28410 35980
rect 29182 35980 29184 36000
rect 29184 35980 29236 36000
rect 29236 35980 29238 36000
rect 29182 35944 29238 35980
rect 28722 34720 28778 34776
rect 28538 34604 28594 34640
rect 28538 34584 28540 34604
rect 28540 34584 28592 34604
rect 28592 34584 28594 34604
rect 28446 33224 28502 33280
rect 28446 32836 28502 32872
rect 28446 32816 28448 32836
rect 28448 32816 28500 32836
rect 28500 32816 28502 32836
rect 27986 19216 28042 19272
rect 28538 20576 28594 20632
rect 30562 35944 30618 36000
rect 29826 33224 29882 33280
rect 28262 16788 28318 16824
rect 28262 16768 28264 16788
rect 28264 16768 28316 16788
rect 28316 16768 28318 16788
rect 27710 14320 27766 14376
rect 28906 20340 28908 20360
rect 28908 20340 28960 20360
rect 28960 20340 28962 20360
rect 28906 20304 28962 20340
rect 28906 20052 28962 20088
rect 28906 20032 28908 20052
rect 28908 20032 28960 20052
rect 28960 20032 28962 20052
rect 28998 19252 29000 19272
rect 29000 19252 29052 19272
rect 29052 19252 29054 19272
rect 28998 19216 29054 19252
rect 28630 17876 28686 17912
rect 28630 17856 28632 17876
rect 28632 17856 28684 17876
rect 28684 17856 28686 17876
rect 29182 17332 29238 17368
rect 29182 17312 29184 17332
rect 29184 17312 29236 17332
rect 29236 17312 29238 17332
rect 28998 16360 29054 16416
rect 28446 15428 28502 15464
rect 28446 15408 28448 15428
rect 28448 15408 28500 15428
rect 28500 15408 28502 15428
rect 28538 14340 28594 14376
rect 28538 14320 28540 14340
rect 28540 14320 28592 14340
rect 28592 14320 28594 14340
rect 28446 13524 28502 13560
rect 28446 13504 28448 13524
rect 28448 13504 28500 13524
rect 28500 13504 28502 13524
rect 31022 34604 31078 34640
rect 31022 34584 31024 34604
rect 31024 34584 31076 34604
rect 31076 34584 31078 34604
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 31206 34584 31262 34640
rect 29734 19932 29736 19952
rect 29736 19932 29788 19952
rect 29788 19932 29790 19952
rect 29734 19896 29790 19932
rect 29826 19624 29882 19680
rect 29734 19216 29790 19272
rect 30378 23468 30380 23488
rect 30380 23468 30432 23488
rect 30432 23468 30434 23488
rect 30378 23432 30434 23468
rect 30378 20576 30434 20632
rect 30286 18672 30342 18728
rect 30378 17740 30434 17776
rect 30378 17720 30380 17740
rect 30380 17720 30432 17740
rect 30432 17720 30434 17740
rect 29734 9832 29790 9888
rect 31206 16224 31262 16280
rect 30838 14900 30840 14920
rect 30840 14900 30892 14920
rect 30892 14900 30894 14920
rect 30838 14864 30894 14900
rect 31206 14864 31262 14920
rect 31942 20476 31944 20496
rect 31944 20476 31996 20496
rect 31996 20476 31998 20496
rect 31942 20440 31998 20476
rect 32310 32952 32366 33008
rect 32678 34348 32680 34368
rect 32680 34348 32732 34368
rect 32732 34348 32734 34368
rect 32678 34312 32734 34348
rect 32770 30504 32826 30560
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 31666 15544 31722 15600
rect 32678 19896 32734 19952
rect 33046 26152 33102 26208
rect 33322 26152 33378 26208
rect 33138 22208 33194 22264
rect 32310 17856 32366 17912
rect 32954 19352 33010 19408
rect 32770 16516 32826 16552
rect 32770 16496 32772 16516
rect 32772 16496 32824 16516
rect 32824 16496 32826 16516
rect 32954 13640 33010 13696
rect 33966 27648 34022 27704
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34794 31184 34850 31240
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34610 30096 34666 30152
rect 35254 30132 35256 30152
rect 35256 30132 35308 30152
rect 35308 30132 35310 30152
rect 35254 30096 35310 30132
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34242 23432 34298 23488
rect 34058 19488 34114 19544
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 36726 38800 36782 38856
rect 36266 37440 36322 37496
rect 35622 34584 35678 34640
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35622 25336 35678 25392
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34794 21004 34850 21040
rect 34794 20984 34796 21004
rect 34796 20984 34848 21004
rect 34848 20984 34850 21004
rect 34610 20440 34666 20496
rect 34610 20304 34666 20360
rect 34242 16496 34298 16552
rect 34426 16496 34482 16552
rect 34794 20304 34850 20360
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34886 19352 34942 19408
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35254 18808 35310 18864
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 36082 31764 36084 31784
rect 36084 31764 36136 31784
rect 36136 31764 36138 31784
rect 36082 31728 36138 31764
rect 36358 23468 36360 23488
rect 36360 23468 36412 23488
rect 36412 23468 36414 23488
rect 36358 23432 36414 23468
rect 35898 18708 35900 18728
rect 35900 18708 35952 18728
rect 35952 18708 35954 18728
rect 35898 18672 35954 18708
rect 36082 18128 36138 18184
rect 35898 17176 35954 17232
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 36726 20052 36782 20088
rect 36726 20032 36728 20052
rect 36728 20032 36780 20052
rect 36780 20032 36782 20052
rect 37462 32680 37518 32736
rect 37278 19624 37334 19680
rect 37554 18128 37610 18184
rect 38198 36080 38254 36136
rect 38198 35436 38200 35456
rect 38200 35436 38252 35456
rect 38252 35436 38254 35456
rect 38198 35400 38254 35436
rect 38198 34040 38254 34096
rect 38290 32000 38346 32056
rect 38290 30640 38346 30696
rect 38106 29280 38162 29336
rect 36818 12280 36874 12336
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38290 28600 38346 28656
rect 38290 27240 38346 27296
rect 38198 26832 38254 26888
rect 38290 25880 38346 25936
rect 38198 25200 38254 25256
rect 38290 23840 38346 23896
rect 38198 22500 38254 22536
rect 38198 22480 38200 22500
rect 38200 22480 38252 22500
rect 38252 22480 38254 22500
rect 38198 21836 38200 21856
rect 38200 21836 38252 21856
rect 38252 21836 38254 21856
rect 38198 21800 38254 21836
rect 38198 19116 38200 19136
rect 38200 19116 38252 19136
rect 38252 19116 38254 19136
rect 38198 19080 38254 19116
rect 38198 17060 38254 17096
rect 38198 17040 38200 17060
rect 38200 17040 38252 17060
rect 38252 17040 38254 17060
rect 38198 15680 38254 15736
rect 38106 15020 38162 15056
rect 38106 15000 38108 15020
rect 38108 15000 38160 15020
rect 38160 15000 38162 15020
rect 38198 13676 38200 13696
rect 38200 13676 38252 13696
rect 38252 13676 38254 13696
rect 38198 13640 38254 13676
rect 38198 12280 38254 12336
rect 37462 7520 37518 7576
rect 38198 10920 38254 10976
rect 38198 10260 38254 10296
rect 38198 10240 38200 10260
rect 38200 10240 38252 10260
rect 38252 10240 38254 10260
rect 38290 8880 38346 8936
rect 38290 6840 38346 6896
rect 38198 5516 38200 5536
rect 38200 5516 38252 5536
rect 38252 5516 38254 5536
rect 38198 5480 38254 5516
rect 37462 4120 37518 4176
rect 36818 2080 36874 2136
rect 2870 720 2926 776
rect 38198 3440 38254 3496
rect 37738 720 37794 776
rect 37186 40 37242 96
<< metal3 >>
rect 200 39538 800 39568
rect 3417 39538 3483 39541
rect 200 39536 3483 39538
rect 200 39480 3422 39536
rect 3478 39480 3483 39536
rect 200 39478 3483 39480
rect 200 39448 800 39478
rect 3417 39475 3483 39478
rect 200 38858 800 38888
rect 2865 38858 2931 38861
rect 200 38856 2931 38858
rect 200 38800 2870 38856
rect 2926 38800 2931 38856
rect 200 38798 2931 38800
rect 200 38768 800 38798
rect 2865 38795 2931 38798
rect 36721 38858 36787 38861
rect 39200 38858 39800 38888
rect 36721 38856 39800 38858
rect 36721 38800 36726 38856
rect 36782 38800 39800 38856
rect 36721 38798 39800 38800
rect 36721 38795 36787 38798
rect 39200 38768 39800 38798
rect 4210 37568 4526 37569
rect 200 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 2865 37498 2931 37501
rect 200 37496 2931 37498
rect 200 37440 2870 37496
rect 2926 37440 2931 37496
rect 200 37438 2931 37440
rect 200 37408 800 37438
rect 2865 37435 2931 37438
rect 36261 37498 36327 37501
rect 39200 37498 39800 37528
rect 36261 37496 39800 37498
rect 36261 37440 36266 37496
rect 36322 37440 39800 37496
rect 36261 37438 39800 37440
rect 36261 37435 36327 37438
rect 39200 37408 39800 37438
rect 15929 37226 15995 37229
rect 18873 37226 18939 37229
rect 15929 37224 18939 37226
rect 15929 37168 15934 37224
rect 15990 37168 18878 37224
rect 18934 37168 18939 37224
rect 15929 37166 18939 37168
rect 15929 37163 15995 37166
rect 18873 37163 18939 37166
rect 28073 37226 28139 37229
rect 31293 37226 31359 37229
rect 28073 37224 31359 37226
rect 28073 37168 28078 37224
rect 28134 37168 31298 37224
rect 31354 37168 31359 37224
rect 28073 37166 31359 37168
rect 28073 37163 28139 37166
rect 31293 37163 31359 37166
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 9673 36818 9739 36821
rect 10593 36818 10659 36821
rect 9673 36816 10659 36818
rect 9673 36760 9678 36816
rect 9734 36760 10598 36816
rect 10654 36760 10659 36816
rect 9673 36758 10659 36760
rect 9673 36755 9739 36758
rect 10593 36755 10659 36758
rect 16849 36818 16915 36821
rect 16982 36818 16988 36820
rect 16849 36816 16988 36818
rect 16849 36760 16854 36816
rect 16910 36760 16988 36816
rect 16849 36758 16988 36760
rect 16849 36755 16915 36758
rect 16982 36756 16988 36758
rect 17052 36756 17058 36820
rect 8017 36682 8083 36685
rect 23473 36682 23539 36685
rect 8017 36680 23539 36682
rect 8017 36624 8022 36680
rect 8078 36624 23478 36680
rect 23534 36624 23539 36680
rect 8017 36622 23539 36624
rect 8017 36619 8083 36622
rect 23473 36619 23539 36622
rect 26141 36546 26207 36549
rect 28809 36546 28875 36549
rect 26141 36544 28875 36546
rect 26141 36488 26146 36544
rect 26202 36488 28814 36544
rect 28870 36488 28875 36544
rect 26141 36486 28875 36488
rect 26141 36483 26207 36486
rect 28809 36483 28875 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 10041 36410 10107 36413
rect 16205 36410 16271 36413
rect 17677 36410 17743 36413
rect 10041 36408 17743 36410
rect 10041 36352 10046 36408
rect 10102 36352 16210 36408
rect 16266 36352 17682 36408
rect 17738 36352 17743 36408
rect 10041 36350 17743 36352
rect 10041 36347 10107 36350
rect 16205 36347 16271 36350
rect 17677 36347 17743 36350
rect 1577 36274 1643 36277
rect 26417 36274 26483 36277
rect 1577 36272 26483 36274
rect 1577 36216 1582 36272
rect 1638 36216 26422 36272
rect 26478 36216 26483 36272
rect 1577 36214 26483 36216
rect 1577 36211 1643 36214
rect 26417 36211 26483 36214
rect 27981 36274 28047 36277
rect 28441 36274 28507 36277
rect 27981 36272 28507 36274
rect 27981 36216 27986 36272
rect 28042 36216 28446 36272
rect 28502 36216 28507 36272
rect 27981 36214 28507 36216
rect 27981 36211 28047 36214
rect 28441 36211 28507 36214
rect 200 36138 800 36168
rect 1393 36138 1459 36141
rect 200 36136 1459 36138
rect 200 36080 1398 36136
rect 1454 36080 1459 36136
rect 200 36078 1459 36080
rect 200 36048 800 36078
rect 1393 36075 1459 36078
rect 6729 36138 6795 36141
rect 26049 36138 26115 36141
rect 6729 36136 26115 36138
rect 6729 36080 6734 36136
rect 6790 36080 26054 36136
rect 26110 36080 26115 36136
rect 6729 36078 26115 36080
rect 6729 36075 6795 36078
rect 26049 36075 26115 36078
rect 27705 36138 27771 36141
rect 28625 36138 28691 36141
rect 27705 36136 28691 36138
rect 27705 36080 27710 36136
rect 27766 36080 28630 36136
rect 28686 36080 28691 36136
rect 27705 36078 28691 36080
rect 27705 36075 27771 36078
rect 28625 36075 28691 36078
rect 38193 36138 38259 36141
rect 39200 36138 39800 36168
rect 38193 36136 39800 36138
rect 38193 36080 38198 36136
rect 38254 36080 39800 36136
rect 38193 36078 39800 36080
rect 38193 36075 38259 36078
rect 39200 36048 39800 36078
rect 11513 36002 11579 36005
rect 13813 36002 13879 36005
rect 11513 36000 13879 36002
rect 11513 35944 11518 36000
rect 11574 35944 13818 36000
rect 13874 35944 13879 36000
rect 11513 35942 13879 35944
rect 11513 35939 11579 35942
rect 13813 35939 13879 35942
rect 14273 36002 14339 36005
rect 16941 36002 17007 36005
rect 14273 36000 17007 36002
rect 14273 35944 14278 36000
rect 14334 35944 16946 36000
rect 17002 35944 17007 36000
rect 14273 35942 17007 35944
rect 14273 35939 14339 35942
rect 16941 35939 17007 35942
rect 22093 36004 22159 36005
rect 26233 36004 26299 36005
rect 22093 36000 22140 36004
rect 22204 36002 22210 36004
rect 26182 36002 26188 36004
rect 22093 35944 22098 36000
rect 22093 35940 22140 35944
rect 22204 35942 22250 36002
rect 26142 35942 26188 36002
rect 26252 36000 26299 36004
rect 26294 35944 26299 36000
rect 22204 35940 22210 35942
rect 26182 35940 26188 35942
rect 26252 35940 26299 35944
rect 22093 35939 22159 35940
rect 26233 35939 26299 35940
rect 28349 36002 28415 36005
rect 29177 36002 29243 36005
rect 28349 36000 29243 36002
rect 28349 35944 28354 36000
rect 28410 35944 29182 36000
rect 29238 35944 29243 36000
rect 28349 35942 29243 35944
rect 28349 35939 28415 35942
rect 29177 35939 29243 35942
rect 29310 35940 29316 36004
rect 29380 36002 29386 36004
rect 30557 36002 30623 36005
rect 29380 36000 30623 36002
rect 29380 35944 30562 36000
rect 30618 35944 30623 36000
rect 29380 35942 30623 35944
rect 29380 35940 29386 35942
rect 30557 35939 30623 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 10777 35866 10843 35869
rect 11789 35866 11855 35869
rect 10777 35864 11855 35866
rect 10777 35808 10782 35864
rect 10838 35808 11794 35864
rect 11850 35808 11855 35864
rect 10777 35806 11855 35808
rect 10777 35803 10843 35806
rect 11789 35803 11855 35806
rect 11973 35866 12039 35869
rect 18413 35866 18479 35869
rect 11973 35864 18479 35866
rect 11973 35808 11978 35864
rect 12034 35808 18418 35864
rect 18474 35808 18479 35864
rect 11973 35806 18479 35808
rect 11973 35803 12039 35806
rect 18413 35803 18479 35806
rect 3049 35730 3115 35733
rect 20897 35730 20963 35733
rect 3049 35728 20963 35730
rect 3049 35672 3054 35728
rect 3110 35672 20902 35728
rect 20958 35672 20963 35728
rect 3049 35670 20963 35672
rect 3049 35667 3115 35670
rect 20897 35667 20963 35670
rect 2313 35594 2379 35597
rect 17125 35594 17191 35597
rect 17769 35594 17835 35597
rect 2313 35592 17835 35594
rect 2313 35536 2318 35592
rect 2374 35536 17130 35592
rect 17186 35536 17774 35592
rect 17830 35536 17835 35592
rect 2313 35534 17835 35536
rect 2313 35531 2379 35534
rect 17125 35531 17191 35534
rect 17769 35531 17835 35534
rect 200 35368 800 35488
rect 10133 35458 10199 35461
rect 13537 35458 13603 35461
rect 10133 35456 13603 35458
rect 10133 35400 10138 35456
rect 10194 35400 13542 35456
rect 13598 35400 13603 35456
rect 10133 35398 13603 35400
rect 10133 35395 10199 35398
rect 13537 35395 13603 35398
rect 38193 35458 38259 35461
rect 39200 35458 39800 35488
rect 38193 35456 39800 35458
rect 38193 35400 38198 35456
rect 38254 35400 39800 35456
rect 38193 35398 39800 35400
rect 38193 35395 38259 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 39800 35398
rect 34930 35327 35246 35328
rect 10501 35322 10567 35325
rect 17401 35322 17467 35325
rect 10501 35320 17467 35322
rect 10501 35264 10506 35320
rect 10562 35264 17406 35320
rect 17462 35264 17467 35320
rect 10501 35262 17467 35264
rect 10501 35259 10567 35262
rect 17401 35259 17467 35262
rect 6453 35186 6519 35189
rect 17953 35186 18019 35189
rect 6453 35184 18019 35186
rect 6453 35128 6458 35184
rect 6514 35128 17958 35184
rect 18014 35128 18019 35184
rect 6453 35126 18019 35128
rect 6453 35123 6519 35126
rect 17953 35123 18019 35126
rect 20345 35050 20411 35053
rect 22921 35050 22987 35053
rect 20345 35048 22987 35050
rect 20345 34992 20350 35048
rect 20406 34992 22926 35048
rect 22982 34992 22987 35048
rect 20345 34990 22987 34992
rect 20345 34987 20411 34990
rect 22921 34987 22987 34990
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 10961 34778 11027 34781
rect 15285 34778 15351 34781
rect 10961 34776 15351 34778
rect 10961 34720 10966 34776
rect 11022 34720 15290 34776
rect 15346 34720 15351 34776
rect 10961 34718 15351 34720
rect 10961 34715 11027 34718
rect 15285 34715 15351 34718
rect 28717 34780 28783 34781
rect 28717 34776 28764 34780
rect 28828 34778 28834 34780
rect 28717 34720 28722 34776
rect 28717 34716 28764 34720
rect 28828 34718 28874 34778
rect 28828 34716 28834 34718
rect 28717 34715 28783 34716
rect 14181 34642 14247 34645
rect 15745 34642 15811 34645
rect 14181 34640 15811 34642
rect 14181 34584 14186 34640
rect 14242 34584 15750 34640
rect 15806 34584 15811 34640
rect 14181 34582 15811 34584
rect 14181 34579 14247 34582
rect 15745 34579 15811 34582
rect 28533 34644 28599 34645
rect 28533 34640 28580 34644
rect 28644 34642 28650 34644
rect 31017 34642 31083 34645
rect 28533 34584 28538 34640
rect 28533 34580 28580 34584
rect 28644 34582 28690 34642
rect 30974 34640 31083 34642
rect 30974 34584 31022 34640
rect 31078 34584 31083 34640
rect 28644 34580 28650 34582
rect 28533 34579 28599 34580
rect 30974 34579 31083 34584
rect 31201 34642 31267 34645
rect 31334 34642 31340 34644
rect 31201 34640 31340 34642
rect 31201 34584 31206 34640
rect 31262 34584 31340 34640
rect 31201 34582 31340 34584
rect 31201 34579 31267 34582
rect 31334 34580 31340 34582
rect 31404 34580 31410 34644
rect 35617 34642 35683 34645
rect 35750 34642 35756 34644
rect 35617 34640 35756 34642
rect 35617 34584 35622 34640
rect 35678 34584 35756 34640
rect 35617 34582 35756 34584
rect 35617 34579 35683 34582
rect 35750 34580 35756 34582
rect 35820 34580 35826 34644
rect 26233 34506 26299 34509
rect 30974 34508 31034 34579
rect 30966 34506 30972 34508
rect 26233 34504 30972 34506
rect 26233 34448 26238 34504
rect 26294 34448 30972 34504
rect 26233 34446 30972 34448
rect 26233 34443 26299 34446
rect 30966 34444 30972 34446
rect 31036 34444 31042 34508
rect 32673 34370 32739 34373
rect 32990 34370 32996 34372
rect 32673 34368 32996 34370
rect 32673 34312 32678 34368
rect 32734 34312 32996 34368
rect 32673 34310 32996 34312
rect 32673 34307 32739 34310
rect 32990 34308 32996 34310
rect 33060 34308 33066 34372
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 200 34098 800 34128
rect 1761 34098 1827 34101
rect 200 34096 1827 34098
rect 200 34040 1766 34096
rect 1822 34040 1827 34096
rect 200 34038 1827 34040
rect 200 34008 800 34038
rect 1761 34035 1827 34038
rect 38193 34098 38259 34101
rect 39200 34098 39800 34128
rect 38193 34096 39800 34098
rect 38193 34040 38198 34096
rect 38254 34040 39800 34096
rect 38193 34038 39800 34040
rect 38193 34035 38259 34038
rect 39200 34008 39800 34038
rect 2313 33962 2379 33965
rect 9397 33962 9463 33965
rect 2313 33960 9463 33962
rect 2313 33904 2318 33960
rect 2374 33904 9402 33960
rect 9458 33904 9463 33960
rect 2313 33902 9463 33904
rect 2313 33899 2379 33902
rect 9397 33899 9463 33902
rect 15929 33962 15995 33965
rect 21173 33962 21239 33965
rect 15929 33960 21239 33962
rect 15929 33904 15934 33960
rect 15990 33904 21178 33960
rect 21234 33904 21239 33960
rect 15929 33902 21239 33904
rect 15929 33899 15995 33902
rect 21173 33899 21239 33902
rect 8201 33826 8267 33829
rect 17125 33826 17191 33829
rect 8201 33824 17191 33826
rect 8201 33768 8206 33824
rect 8262 33768 17130 33824
rect 17186 33768 17191 33824
rect 8201 33766 17191 33768
rect 8201 33763 8267 33766
rect 17125 33763 17191 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 12065 33690 12131 33693
rect 19425 33690 19491 33693
rect 12065 33688 19491 33690
rect 12065 33632 12070 33688
rect 12126 33632 19430 33688
rect 19486 33632 19491 33688
rect 12065 33630 19491 33632
rect 12065 33627 12131 33630
rect 19425 33627 19491 33630
rect 10961 33554 11027 33557
rect 26233 33554 26299 33557
rect 10961 33552 26299 33554
rect 10961 33496 10966 33552
rect 11022 33496 26238 33552
rect 26294 33496 26299 33552
rect 10961 33494 26299 33496
rect 10961 33491 11027 33494
rect 26233 33491 26299 33494
rect 17769 33418 17835 33421
rect 20897 33418 20963 33421
rect 17769 33416 20963 33418
rect 17769 33360 17774 33416
rect 17830 33360 20902 33416
rect 20958 33360 20963 33416
rect 17769 33358 20963 33360
rect 17769 33355 17835 33358
rect 20897 33355 20963 33358
rect 12893 33282 12959 33285
rect 28022 33282 28028 33284
rect 12893 33280 28028 33282
rect 12893 33224 12898 33280
rect 12954 33224 28028 33280
rect 12893 33222 28028 33224
rect 12893 33219 12959 33222
rect 28022 33220 28028 33222
rect 28092 33282 28098 33284
rect 28441 33282 28507 33285
rect 28092 33280 28507 33282
rect 28092 33224 28446 33280
rect 28502 33224 28507 33280
rect 28092 33222 28507 33224
rect 28092 33220 28098 33222
rect 28441 33219 28507 33222
rect 29821 33284 29887 33285
rect 29821 33280 29868 33284
rect 29932 33282 29938 33284
rect 29821 33224 29826 33280
rect 29821 33220 29868 33224
rect 29932 33222 29978 33282
rect 29932 33220 29938 33222
rect 29821 33219 29887 33220
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 15469 33146 15535 33149
rect 16297 33146 16363 33149
rect 18413 33146 18479 33149
rect 15469 33144 18479 33146
rect 15469 33088 15474 33144
rect 15530 33088 16302 33144
rect 16358 33088 18418 33144
rect 18474 33088 18479 33144
rect 15469 33086 18479 33088
rect 15469 33083 15535 33086
rect 16297 33083 16363 33086
rect 18413 33083 18479 33086
rect 19425 33146 19491 33149
rect 21541 33146 21607 33149
rect 19425 33144 21607 33146
rect 19425 33088 19430 33144
rect 19486 33088 21546 33144
rect 21602 33088 21607 33144
rect 19425 33086 21607 33088
rect 19425 33083 19491 33086
rect 21541 33083 21607 33086
rect 10225 33010 10291 33013
rect 32305 33010 32371 33013
rect 10225 33008 32371 33010
rect 10225 32952 10230 33008
rect 10286 32952 32310 33008
rect 32366 32952 32371 33008
rect 10225 32950 32371 32952
rect 10225 32947 10291 32950
rect 32305 32947 32371 32950
rect 16941 32874 17007 32877
rect 17493 32874 17559 32877
rect 28441 32876 28507 32877
rect 16941 32872 17559 32874
rect 16941 32816 16946 32872
rect 17002 32816 17498 32872
rect 17554 32816 17559 32872
rect 16941 32814 17559 32816
rect 16941 32811 17007 32814
rect 17493 32811 17559 32814
rect 28390 32812 28396 32876
rect 28460 32874 28507 32876
rect 28460 32872 28552 32874
rect 28502 32816 28552 32872
rect 28460 32814 28552 32816
rect 28460 32812 28507 32814
rect 28441 32811 28507 32812
rect 200 32738 800 32768
rect 1761 32738 1827 32741
rect 200 32736 1827 32738
rect 200 32680 1766 32736
rect 1822 32680 1827 32736
rect 200 32678 1827 32680
rect 200 32648 800 32678
rect 1761 32675 1827 32678
rect 9765 32738 9831 32741
rect 19241 32738 19307 32741
rect 9765 32736 19307 32738
rect 9765 32680 9770 32736
rect 9826 32680 19246 32736
rect 19302 32680 19307 32736
rect 9765 32678 19307 32680
rect 9765 32675 9831 32678
rect 19241 32675 19307 32678
rect 37457 32738 37523 32741
rect 39200 32738 39800 32768
rect 37457 32736 39800 32738
rect 37457 32680 37462 32736
rect 37518 32680 39800 32736
rect 37457 32678 39800 32680
rect 37457 32675 37523 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 39800 32678
rect 19570 32607 19886 32608
rect 12985 32602 13051 32605
rect 18045 32602 18111 32605
rect 12985 32600 18111 32602
rect 12985 32544 12990 32600
rect 13046 32544 18050 32600
rect 18106 32544 18111 32600
rect 12985 32542 18111 32544
rect 12985 32539 13051 32542
rect 18045 32539 18111 32542
rect 12341 32466 12407 32469
rect 12801 32466 12867 32469
rect 12341 32464 12867 32466
rect 12341 32408 12346 32464
rect 12402 32408 12806 32464
rect 12862 32408 12867 32464
rect 12341 32406 12867 32408
rect 12341 32403 12407 32406
rect 12801 32403 12867 32406
rect 11697 32330 11763 32333
rect 15193 32330 15259 32333
rect 11697 32328 15259 32330
rect 11697 32272 11702 32328
rect 11758 32272 15198 32328
rect 15254 32272 15259 32328
rect 11697 32270 15259 32272
rect 11697 32267 11763 32270
rect 15193 32267 15259 32270
rect 4210 32128 4526 32129
rect 200 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1761 32058 1827 32061
rect 200 32056 1827 32058
rect 200 32000 1766 32056
rect 1822 32000 1827 32056
rect 200 31998 1827 32000
rect 200 31968 800 31998
rect 1761 31995 1827 31998
rect 38285 32058 38351 32061
rect 39200 32058 39800 32088
rect 38285 32056 39800 32058
rect 38285 32000 38290 32056
rect 38346 32000 39800 32056
rect 38285 31998 39800 32000
rect 38285 31995 38351 31998
rect 39200 31968 39800 31998
rect 36077 31786 36143 31789
rect 36854 31786 36860 31788
rect 36077 31784 36860 31786
rect 36077 31728 36082 31784
rect 36138 31728 36860 31784
rect 36077 31726 36860 31728
rect 36077 31723 36143 31726
rect 36854 31724 36860 31726
rect 36924 31724 36930 31788
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 25814 31180 25820 31244
rect 25884 31242 25890 31244
rect 34789 31242 34855 31245
rect 25884 31240 34855 31242
rect 25884 31184 34794 31240
rect 34850 31184 34855 31240
rect 25884 31182 34855 31184
rect 25884 31180 25890 31182
rect 34789 31179 34855 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 38285 30698 38351 30701
rect 39200 30698 39800 30728
rect 38285 30696 39800 30698
rect 38285 30640 38290 30696
rect 38346 30640 39800 30696
rect 38285 30638 39800 30640
rect 38285 30635 38351 30638
rect 39200 30608 39800 30638
rect 25998 30500 26004 30564
rect 26068 30562 26074 30564
rect 32765 30562 32831 30565
rect 26068 30560 32831 30562
rect 26068 30504 32770 30560
rect 32826 30504 32831 30560
rect 26068 30502 32831 30504
rect 26068 30500 26074 30502
rect 32765 30499 32831 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 11421 30426 11487 30429
rect 12934 30426 12940 30428
rect 11421 30424 12940 30426
rect 11421 30368 11426 30424
rect 11482 30368 12940 30424
rect 11421 30366 12940 30368
rect 11421 30363 11487 30366
rect 12934 30364 12940 30366
rect 13004 30364 13010 30428
rect 14365 30290 14431 30293
rect 15469 30290 15535 30293
rect 14365 30288 15535 30290
rect 14365 30232 14370 30288
rect 14426 30232 15474 30288
rect 15530 30232 15535 30288
rect 14365 30230 15535 30232
rect 14365 30227 14431 30230
rect 15469 30227 15535 30230
rect 34462 30092 34468 30156
rect 34532 30154 34538 30156
rect 34605 30154 34671 30157
rect 35249 30154 35315 30157
rect 34532 30152 35315 30154
rect 34532 30096 34610 30152
rect 34666 30096 35254 30152
rect 35310 30096 35315 30152
rect 34532 30094 35315 30096
rect 34532 30092 34538 30094
rect 34605 30091 34671 30094
rect 35249 30091 35315 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1761 29338 1827 29341
rect 200 29336 1827 29338
rect 200 29280 1766 29336
rect 1822 29280 1827 29336
rect 200 29278 1827 29280
rect 200 29248 800 29278
rect 1761 29275 1827 29278
rect 38101 29338 38167 29341
rect 39200 29338 39800 29368
rect 38101 29336 39800 29338
rect 38101 29280 38106 29336
rect 38162 29280 39800 29336
rect 38101 29278 39800 29280
rect 38101 29275 38167 29278
rect 39200 29248 39800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 200 28658 800 28688
rect 1577 28658 1643 28661
rect 200 28656 1643 28658
rect 200 28600 1582 28656
rect 1638 28600 1643 28656
rect 200 28598 1643 28600
rect 200 28568 800 28598
rect 1577 28595 1643 28598
rect 38285 28658 38351 28661
rect 39200 28658 39800 28688
rect 38285 28656 39800 28658
rect 38285 28600 38290 28656
rect 38346 28600 39800 28656
rect 38285 28598 39800 28600
rect 38285 28595 38351 28598
rect 39200 28568 39800 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 12934 27916 12940 27980
rect 13004 27978 13010 27980
rect 13077 27978 13143 27981
rect 13004 27976 13143 27978
rect 13004 27920 13082 27976
rect 13138 27920 13143 27976
rect 13004 27918 13143 27920
rect 13004 27916 13010 27918
rect 13077 27915 13143 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 25957 27708 26023 27709
rect 25446 27644 25452 27708
rect 25516 27706 25522 27708
rect 25957 27706 26004 27708
rect 25516 27704 26004 27706
rect 25516 27648 25962 27704
rect 25516 27646 26004 27648
rect 25516 27644 25522 27646
rect 25957 27644 26004 27646
rect 26068 27644 26074 27708
rect 33174 27644 33180 27708
rect 33244 27706 33250 27708
rect 33961 27706 34027 27709
rect 33244 27704 34027 27706
rect 33244 27648 33966 27704
rect 34022 27648 34027 27704
rect 33244 27646 34027 27648
rect 33244 27644 33250 27646
rect 25957 27643 26023 27644
rect 33961 27643 34027 27646
rect 200 27298 800 27328
rect 1669 27298 1735 27301
rect 200 27296 1735 27298
rect 200 27240 1674 27296
rect 1730 27240 1735 27296
rect 200 27238 1735 27240
rect 200 27208 800 27238
rect 1669 27235 1735 27238
rect 38285 27298 38351 27301
rect 39200 27298 39800 27328
rect 38285 27296 39800 27298
rect 38285 27240 38290 27296
rect 38346 27240 39800 27296
rect 38285 27238 39800 27240
rect 38285 27235 38351 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 39800 27238
rect 19570 27167 19886 27168
rect 23974 26828 23980 26892
rect 24044 26890 24050 26892
rect 38193 26890 38259 26893
rect 24044 26888 38259 26890
rect 24044 26832 38198 26888
rect 38254 26832 38259 26888
rect 24044 26830 38259 26832
rect 24044 26828 24050 26830
rect 38193 26827 38259 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 21449 26346 21515 26349
rect 26734 26346 26740 26348
rect 21449 26344 26740 26346
rect 21449 26288 21454 26344
rect 21510 26288 26740 26344
rect 21449 26286 26740 26288
rect 21449 26283 21515 26286
rect 26734 26284 26740 26286
rect 26804 26346 26810 26348
rect 27429 26346 27495 26349
rect 26804 26344 27495 26346
rect 26804 26288 27434 26344
rect 27490 26288 27495 26344
rect 26804 26286 27495 26288
rect 26804 26284 26810 26286
rect 27429 26283 27495 26286
rect 32438 26148 32444 26212
rect 32508 26210 32514 26212
rect 33041 26210 33107 26213
rect 32508 26208 33107 26210
rect 32508 26152 33046 26208
rect 33102 26152 33107 26208
rect 32508 26150 33107 26152
rect 32508 26148 32514 26150
rect 33041 26147 33107 26150
rect 33317 26210 33383 26213
rect 36670 26210 36676 26212
rect 33317 26208 36676 26210
rect 33317 26152 33322 26208
rect 33378 26152 36676 26208
rect 33317 26150 36676 26152
rect 33317 26147 33383 26150
rect 36670 26148 36676 26150
rect 36740 26148 36746 26212
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 200 25938 800 25968
rect 1761 25938 1827 25941
rect 200 25936 1827 25938
rect 200 25880 1766 25936
rect 1822 25880 1827 25936
rect 200 25878 1827 25880
rect 200 25848 800 25878
rect 1761 25875 1827 25878
rect 38285 25938 38351 25941
rect 39200 25938 39800 25968
rect 38285 25936 39800 25938
rect 38285 25880 38290 25936
rect 38346 25880 39800 25936
rect 38285 25878 39800 25880
rect 38285 25875 38351 25878
rect 39200 25848 39800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 35617 25394 35683 25397
rect 35574 25392 35683 25394
rect 35574 25336 35622 25392
rect 35678 25336 35683 25392
rect 35574 25331 35683 25336
rect 30230 25196 30236 25260
rect 30300 25258 30306 25260
rect 35574 25258 35634 25331
rect 30300 25198 35634 25258
rect 38193 25258 38259 25261
rect 39200 25258 39800 25288
rect 38193 25256 39800 25258
rect 38193 25200 38198 25256
rect 38254 25200 39800 25256
rect 38193 25198 39800 25200
rect 30300 25196 30306 25198
rect 38193 25195 38259 25198
rect 39200 25168 39800 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 21398 24788 21404 24852
rect 21468 24850 21474 24852
rect 21541 24850 21607 24853
rect 21468 24848 21607 24850
rect 21468 24792 21546 24848
rect 21602 24792 21607 24848
rect 21468 24790 21607 24792
rect 21468 24788 21474 24790
rect 21541 24787 21607 24790
rect 24485 24850 24551 24853
rect 27470 24850 27476 24852
rect 24485 24848 27476 24850
rect 24485 24792 24490 24848
rect 24546 24792 27476 24848
rect 24485 24790 27476 24792
rect 24485 24787 24551 24790
rect 27470 24788 27476 24790
rect 27540 24788 27546 24852
rect 200 24578 800 24608
rect 1761 24578 1827 24581
rect 200 24576 1827 24578
rect 200 24520 1766 24576
rect 1822 24520 1827 24576
rect 200 24518 1827 24520
rect 200 24488 800 24518
rect 1761 24515 1827 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 200 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1577 23898 1643 23901
rect 200 23896 1643 23898
rect 200 23840 1582 23896
rect 1638 23840 1643 23896
rect 200 23838 1643 23840
rect 200 23808 800 23838
rect 1577 23835 1643 23838
rect 38285 23898 38351 23901
rect 39200 23898 39800 23928
rect 38285 23896 39800 23898
rect 38285 23840 38290 23896
rect 38346 23840 39800 23896
rect 38285 23838 39800 23840
rect 38285 23835 38351 23838
rect 39200 23808 39800 23838
rect 10961 23762 11027 23765
rect 12934 23762 12940 23764
rect 10961 23760 12940 23762
rect 10961 23704 10966 23760
rect 11022 23704 12940 23760
rect 10961 23702 12940 23704
rect 10961 23699 11027 23702
rect 12934 23700 12940 23702
rect 13004 23700 13010 23764
rect 15285 23626 15351 23629
rect 18597 23626 18663 23629
rect 15285 23624 18663 23626
rect 15285 23568 15290 23624
rect 15346 23568 18602 23624
rect 18658 23568 18663 23624
rect 15285 23566 18663 23568
rect 15285 23563 15351 23566
rect 18597 23563 18663 23566
rect 16982 23428 16988 23492
rect 17052 23490 17058 23492
rect 18597 23490 18663 23493
rect 17052 23488 18663 23490
rect 17052 23432 18602 23488
rect 18658 23432 18663 23488
rect 17052 23430 18663 23432
rect 17052 23428 17058 23430
rect 18597 23427 18663 23430
rect 21214 23428 21220 23492
rect 21284 23490 21290 23492
rect 23841 23490 23907 23493
rect 21284 23488 23907 23490
rect 21284 23432 23846 23488
rect 23902 23432 23907 23488
rect 21284 23430 23907 23432
rect 21284 23428 21290 23430
rect 23841 23427 23907 23430
rect 30373 23492 30439 23493
rect 30373 23488 30420 23492
rect 30484 23490 30490 23492
rect 30373 23432 30378 23488
rect 30373 23428 30420 23432
rect 30484 23430 30530 23490
rect 30484 23428 30490 23430
rect 33726 23428 33732 23492
rect 33796 23490 33802 23492
rect 34237 23490 34303 23493
rect 36353 23492 36419 23493
rect 36302 23490 36308 23492
rect 33796 23488 34303 23490
rect 33796 23432 34242 23488
rect 34298 23432 34303 23488
rect 33796 23430 34303 23432
rect 36262 23430 36308 23490
rect 36372 23488 36419 23492
rect 36414 23432 36419 23488
rect 33796 23428 33802 23430
rect 30373 23427 30439 23428
rect 34237 23427 34303 23430
rect 36302 23428 36308 23430
rect 36372 23428 36419 23432
rect 36353 23427 36419 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 27337 23354 27403 23357
rect 30598 23354 30604 23356
rect 27337 23352 30604 23354
rect 27337 23296 27342 23352
rect 27398 23296 30604 23352
rect 27337 23294 30604 23296
rect 27337 23291 27403 23294
rect 30598 23292 30604 23294
rect 30668 23292 30674 23356
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 200 22538 800 22568
rect 1761 22538 1827 22541
rect 200 22536 1827 22538
rect 200 22480 1766 22536
rect 1822 22480 1827 22536
rect 200 22478 1827 22480
rect 200 22448 800 22478
rect 1761 22475 1827 22478
rect 38193 22538 38259 22541
rect 39200 22538 39800 22568
rect 38193 22536 39800 22538
rect 38193 22480 38198 22536
rect 38254 22480 39800 22536
rect 38193 22478 39800 22480
rect 38193 22475 38259 22478
rect 39200 22448 39800 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 30598 22204 30604 22268
rect 30668 22266 30674 22268
rect 33133 22266 33199 22269
rect 30668 22264 33199 22266
rect 30668 22208 33138 22264
rect 33194 22208 33199 22264
rect 30668 22206 33199 22208
rect 30668 22204 30674 22206
rect 33133 22203 33199 22206
rect 12249 21858 12315 21861
rect 12525 21858 12591 21861
rect 12249 21856 12591 21858
rect 12249 21800 12254 21856
rect 12310 21800 12530 21856
rect 12586 21800 12591 21856
rect 12249 21798 12591 21800
rect 12249 21795 12315 21798
rect 12525 21795 12591 21798
rect 38193 21858 38259 21861
rect 39200 21858 39800 21888
rect 38193 21856 39800 21858
rect 38193 21800 38198 21856
rect 38254 21800 39800 21856
rect 38193 21798 39800 21800
rect 38193 21795 38259 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 39800 21798
rect 19570 21727 19886 21728
rect 12249 21586 12315 21589
rect 13721 21586 13787 21589
rect 18689 21586 18755 21589
rect 12249 21584 18755 21586
rect 12249 21528 12254 21584
rect 12310 21528 13726 21584
rect 13782 21528 18694 21584
rect 18750 21528 18755 21584
rect 12249 21526 18755 21528
rect 12249 21523 12315 21526
rect 13721 21523 13787 21526
rect 18689 21523 18755 21526
rect 12525 21450 12591 21453
rect 15837 21450 15903 21453
rect 12525 21448 15903 21450
rect 12525 21392 12530 21448
rect 12586 21392 15842 21448
rect 15898 21392 15903 21448
rect 12525 21390 15903 21392
rect 12525 21387 12591 21390
rect 15837 21387 15903 21390
rect 11237 21314 11303 21317
rect 10964 21312 11303 21314
rect 10964 21256 11242 21312
rect 11298 21256 11303 21312
rect 10964 21254 11303 21256
rect 4210 21248 4526 21249
rect 200 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 1669 21178 1735 21181
rect 200 21176 1735 21178
rect 200 21120 1674 21176
rect 1730 21120 1735 21176
rect 200 21118 1735 21120
rect 200 21088 800 21118
rect 1669 21115 1735 21118
rect 10964 21045 11024 21254
rect 11237 21251 11303 21254
rect 11789 21314 11855 21317
rect 17217 21314 17283 21317
rect 11789 21312 17283 21314
rect 11789 21256 11794 21312
rect 11850 21256 17222 21312
rect 17278 21256 17283 21312
rect 11789 21254 17283 21256
rect 11789 21251 11855 21254
rect 17217 21251 17283 21254
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 21173 21180 21239 21181
rect 21173 21178 21220 21180
rect 21128 21176 21220 21178
rect 21128 21120 21178 21176
rect 21128 21118 21220 21120
rect 21173 21116 21220 21118
rect 21284 21116 21290 21180
rect 21173 21115 21239 21116
rect 10961 21040 11027 21045
rect 10961 20984 10966 21040
rect 11022 20984 11027 21040
rect 10961 20979 11027 20984
rect 14641 21042 14707 21045
rect 15377 21042 15443 21045
rect 14641 21040 15443 21042
rect 14641 20984 14646 21040
rect 14702 20984 15382 21040
rect 15438 20984 15443 21040
rect 14641 20982 15443 20984
rect 14641 20979 14707 20982
rect 15377 20979 15443 20982
rect 21265 21042 21331 21045
rect 21398 21042 21404 21044
rect 21265 21040 21404 21042
rect 21265 20984 21270 21040
rect 21326 20984 21404 21040
rect 21265 20982 21404 20984
rect 21265 20979 21331 20982
rect 21398 20980 21404 20982
rect 21468 20980 21474 21044
rect 34646 20980 34652 21044
rect 34716 21042 34722 21044
rect 34789 21042 34855 21045
rect 34716 21040 34855 21042
rect 34716 20984 34794 21040
rect 34850 20984 34855 21040
rect 34716 20982 34855 20984
rect 34716 20980 34722 20982
rect 34789 20979 34855 20982
rect 9765 20906 9831 20909
rect 14273 20906 14339 20909
rect 9765 20904 14339 20906
rect 9765 20848 9770 20904
rect 9826 20848 14278 20904
rect 14334 20848 14339 20904
rect 9765 20846 14339 20848
rect 9765 20843 9831 20846
rect 14273 20843 14339 20846
rect 21357 20906 21423 20909
rect 25773 20908 25839 20909
rect 23422 20906 23428 20908
rect 21357 20904 23428 20906
rect 21357 20848 21362 20904
rect 21418 20848 23428 20904
rect 21357 20846 23428 20848
rect 21357 20843 21423 20846
rect 23422 20844 23428 20846
rect 23492 20844 23498 20908
rect 25773 20906 25820 20908
rect 25728 20904 25820 20906
rect 25728 20848 25778 20904
rect 25728 20846 25820 20848
rect 25773 20844 25820 20846
rect 25884 20844 25890 20908
rect 25773 20843 25839 20844
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 25313 20634 25379 20637
rect 28533 20634 28599 20637
rect 25313 20632 28599 20634
rect 25313 20576 25318 20632
rect 25374 20576 28538 20632
rect 28594 20576 28599 20632
rect 25313 20574 28599 20576
rect 25313 20571 25379 20574
rect 28533 20571 28599 20574
rect 30373 20634 30439 20637
rect 30598 20634 30604 20636
rect 30373 20632 30604 20634
rect 30373 20576 30378 20632
rect 30434 20576 30604 20632
rect 30373 20574 30604 20576
rect 30373 20571 30439 20574
rect 30598 20572 30604 20574
rect 30668 20572 30674 20636
rect 200 20498 800 20528
rect 1669 20498 1735 20501
rect 200 20496 1735 20498
rect 200 20440 1674 20496
rect 1730 20440 1735 20496
rect 200 20438 1735 20440
rect 200 20408 800 20438
rect 1669 20435 1735 20438
rect 28574 20436 28580 20500
rect 28644 20498 28650 20500
rect 31937 20498 32003 20501
rect 28644 20496 32003 20498
rect 28644 20440 31942 20496
rect 31998 20440 32003 20496
rect 28644 20438 32003 20440
rect 28644 20436 28650 20438
rect 31937 20435 32003 20438
rect 34605 20498 34671 20501
rect 39200 20498 39800 20528
rect 34605 20496 39800 20498
rect 34605 20440 34610 20496
rect 34666 20440 39800 20496
rect 34605 20438 39800 20440
rect 34605 20435 34671 20438
rect 39200 20408 39800 20438
rect 25681 20362 25747 20365
rect 28901 20362 28967 20365
rect 25681 20360 28967 20362
rect 25681 20304 25686 20360
rect 25742 20304 28906 20360
rect 28962 20304 28967 20360
rect 25681 20302 28967 20304
rect 25681 20299 25747 20302
rect 28901 20299 28967 20302
rect 34605 20362 34671 20365
rect 34789 20362 34855 20365
rect 34605 20360 34855 20362
rect 34605 20304 34610 20360
rect 34666 20304 34794 20360
rect 34850 20304 34855 20360
rect 34605 20302 34855 20304
rect 34605 20299 34671 20302
rect 34789 20299 34855 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 27470 20028 27476 20092
rect 27540 20090 27546 20092
rect 28901 20090 28967 20093
rect 36721 20092 36787 20093
rect 27540 20088 28967 20090
rect 27540 20032 28906 20088
rect 28962 20032 28967 20088
rect 27540 20030 28967 20032
rect 27540 20028 27546 20030
rect 28901 20027 28967 20030
rect 36670 20028 36676 20092
rect 36740 20090 36787 20092
rect 36740 20088 36832 20090
rect 36782 20032 36832 20088
rect 36740 20030 36832 20032
rect 36740 20028 36787 20030
rect 36721 20027 36787 20028
rect 29729 19954 29795 19957
rect 32673 19954 32739 19957
rect 29729 19952 32739 19954
rect 29729 19896 29734 19952
rect 29790 19896 32678 19952
rect 32734 19896 32739 19952
rect 29729 19894 32739 19896
rect 29729 19891 29795 19894
rect 32673 19891 32739 19894
rect 29821 19682 29887 19685
rect 37273 19682 37339 19685
rect 29821 19680 37339 19682
rect 29821 19624 29826 19680
rect 29882 19624 37278 19680
rect 37334 19624 37339 19680
rect 29821 19622 37339 19624
rect 29821 19619 29887 19622
rect 37273 19619 37339 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 34053 19546 34119 19549
rect 34462 19546 34468 19548
rect 34053 19544 34468 19546
rect 34053 19488 34058 19544
rect 34114 19488 34468 19544
rect 34053 19486 34468 19488
rect 34053 19483 34119 19486
rect 34462 19484 34468 19486
rect 34532 19484 34538 19548
rect 32949 19410 33015 19413
rect 33174 19410 33180 19412
rect 32949 19408 33180 19410
rect 32949 19352 32954 19408
rect 33010 19352 33180 19408
rect 32949 19350 33180 19352
rect 32949 19347 33015 19350
rect 33174 19348 33180 19350
rect 33244 19348 33250 19412
rect 34462 19348 34468 19412
rect 34532 19410 34538 19412
rect 34881 19410 34947 19413
rect 34532 19408 34947 19410
rect 34532 19352 34886 19408
rect 34942 19352 34947 19408
rect 34532 19350 34947 19352
rect 34532 19348 34538 19350
rect 34881 19347 34947 19350
rect 27981 19276 28047 19277
rect 27981 19272 28028 19276
rect 28092 19274 28098 19276
rect 27981 19216 27986 19272
rect 27981 19212 28028 19216
rect 28092 19214 28138 19274
rect 28092 19212 28098 19214
rect 28758 19212 28764 19276
rect 28828 19274 28834 19276
rect 28993 19274 29059 19277
rect 28828 19272 29059 19274
rect 28828 19216 28998 19272
rect 29054 19216 29059 19272
rect 28828 19214 29059 19216
rect 28828 19212 28834 19214
rect 27981 19211 28047 19212
rect 28993 19211 29059 19214
rect 29729 19274 29795 19277
rect 30230 19274 30236 19276
rect 29729 19272 30236 19274
rect 29729 19216 29734 19272
rect 29790 19216 30236 19272
rect 29729 19214 30236 19216
rect 29729 19211 29795 19214
rect 30230 19212 30236 19214
rect 30300 19212 30306 19276
rect 200 19138 800 19168
rect 1761 19138 1827 19141
rect 200 19136 1827 19138
rect 200 19080 1766 19136
rect 1822 19080 1827 19136
rect 200 19078 1827 19080
rect 200 19048 800 19078
rect 1761 19075 1827 19078
rect 21265 19138 21331 19141
rect 26325 19138 26391 19141
rect 21265 19136 26391 19138
rect 21265 19080 21270 19136
rect 21326 19080 26330 19136
rect 26386 19080 26391 19136
rect 21265 19078 26391 19080
rect 21265 19075 21331 19078
rect 26325 19075 26391 19078
rect 38193 19138 38259 19141
rect 39200 19138 39800 19168
rect 38193 19136 39800 19138
rect 38193 19080 38198 19136
rect 38254 19080 39800 19136
rect 38193 19078 39800 19080
rect 38193 19075 38259 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 22134 18940 22140 19004
rect 22204 19002 22210 19004
rect 26325 19002 26391 19005
rect 22204 19000 26391 19002
rect 22204 18944 26330 19000
rect 26386 18944 26391 19000
rect 22204 18942 26391 18944
rect 22204 18940 22210 18942
rect 26325 18939 26391 18942
rect 35249 18866 35315 18869
rect 35750 18866 35756 18868
rect 35249 18864 35756 18866
rect 35249 18808 35254 18864
rect 35310 18808 35756 18864
rect 35249 18806 35756 18808
rect 35249 18803 35315 18806
rect 35750 18804 35756 18806
rect 35820 18804 35826 18868
rect 30281 18730 30347 18733
rect 35893 18730 35959 18733
rect 30281 18728 35959 18730
rect 30281 18672 30286 18728
rect 30342 18672 35898 18728
rect 35954 18672 35959 18728
rect 30281 18670 35959 18672
rect 30281 18667 30347 18670
rect 35893 18667 35959 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 24209 18458 24275 18461
rect 25446 18458 25452 18460
rect 24209 18456 25452 18458
rect 24209 18400 24214 18456
rect 24270 18400 25452 18456
rect 24209 18398 25452 18400
rect 24209 18395 24275 18398
rect 25446 18396 25452 18398
rect 25516 18396 25522 18460
rect 26049 18458 26115 18461
rect 26182 18458 26188 18460
rect 26049 18456 26188 18458
rect 26049 18400 26054 18456
rect 26110 18400 26188 18456
rect 26049 18398 26188 18400
rect 26049 18395 26115 18398
rect 26182 18396 26188 18398
rect 26252 18396 26258 18460
rect 39200 18368 39800 18488
rect 31334 18124 31340 18188
rect 31404 18186 31410 18188
rect 36077 18186 36143 18189
rect 37549 18186 37615 18189
rect 31404 18184 37615 18186
rect 31404 18128 36082 18184
rect 36138 18128 37554 18184
rect 37610 18128 37615 18184
rect 31404 18126 37615 18128
rect 31404 18124 31410 18126
rect 36077 18123 36143 18126
rect 37549 18123 37615 18126
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 23013 17914 23079 17917
rect 23974 17914 23980 17916
rect 23013 17912 23980 17914
rect 23013 17856 23018 17912
rect 23074 17856 23980 17912
rect 23013 17854 23980 17856
rect 23013 17851 23079 17854
rect 23974 17852 23980 17854
rect 24044 17852 24050 17916
rect 28625 17914 28691 17917
rect 29862 17914 29868 17916
rect 28625 17912 29868 17914
rect 28625 17856 28630 17912
rect 28686 17856 29868 17912
rect 28625 17854 29868 17856
rect 28625 17851 28691 17854
rect 29862 17852 29868 17854
rect 29932 17852 29938 17916
rect 32305 17914 32371 17917
rect 32438 17914 32444 17916
rect 32305 17912 32444 17914
rect 32305 17856 32310 17912
rect 32366 17856 32444 17912
rect 32305 17854 32444 17856
rect 32305 17851 32371 17854
rect 32438 17852 32444 17854
rect 32508 17852 32514 17916
rect 200 17778 800 17808
rect 1577 17778 1643 17781
rect 200 17776 1643 17778
rect 200 17720 1582 17776
rect 1638 17720 1643 17776
rect 200 17718 1643 17720
rect 200 17688 800 17718
rect 1577 17715 1643 17718
rect 13261 17778 13327 17781
rect 30373 17778 30439 17781
rect 34462 17778 34468 17780
rect 13261 17776 34468 17778
rect 13261 17720 13266 17776
rect 13322 17720 30378 17776
rect 30434 17720 34468 17776
rect 13261 17718 34468 17720
rect 13261 17715 13327 17718
rect 30373 17715 30439 17718
rect 34462 17716 34468 17718
rect 34532 17716 34538 17780
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 29177 17370 29243 17373
rect 29310 17370 29316 17372
rect 29177 17368 29316 17370
rect 29177 17312 29182 17368
rect 29238 17312 29316 17368
rect 29177 17310 29316 17312
rect 29177 17307 29243 17310
rect 29310 17308 29316 17310
rect 29380 17308 29386 17372
rect 12934 17172 12940 17236
rect 13004 17234 13010 17236
rect 35893 17234 35959 17237
rect 13004 17232 35959 17234
rect 13004 17176 35898 17232
rect 35954 17176 35959 17232
rect 13004 17174 35959 17176
rect 13004 17172 13010 17174
rect 35893 17171 35959 17174
rect 200 17098 800 17128
rect 1761 17098 1827 17101
rect 200 17096 1827 17098
rect 200 17040 1766 17096
rect 1822 17040 1827 17096
rect 200 17038 1827 17040
rect 200 17008 800 17038
rect 1761 17035 1827 17038
rect 38193 17098 38259 17101
rect 39200 17098 39800 17128
rect 38193 17096 39800 17098
rect 38193 17040 38198 17096
rect 38254 17040 39800 17096
rect 38193 17038 39800 17040
rect 38193 17035 38259 17038
rect 39200 17008 39800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 28257 16826 28323 16829
rect 28390 16826 28396 16828
rect 28257 16824 28396 16826
rect 28257 16768 28262 16824
rect 28318 16768 28396 16824
rect 28257 16766 28396 16768
rect 28257 16763 28323 16766
rect 28390 16764 28396 16766
rect 28460 16764 28466 16828
rect 30966 16492 30972 16556
rect 31036 16554 31042 16556
rect 32765 16554 32831 16557
rect 31036 16552 32831 16554
rect 31036 16496 32770 16552
rect 32826 16496 32831 16552
rect 31036 16494 32831 16496
rect 31036 16492 31042 16494
rect 32765 16491 32831 16494
rect 33726 16492 33732 16556
rect 33796 16554 33802 16556
rect 34237 16554 34303 16557
rect 33796 16552 34303 16554
rect 33796 16496 34242 16552
rect 34298 16496 34303 16552
rect 33796 16494 34303 16496
rect 33796 16492 33802 16494
rect 34237 16491 34303 16494
rect 34421 16554 34487 16557
rect 34646 16554 34652 16556
rect 34421 16552 34652 16554
rect 34421 16496 34426 16552
rect 34482 16496 34652 16552
rect 34421 16494 34652 16496
rect 34421 16491 34487 16494
rect 34646 16492 34652 16494
rect 34716 16492 34722 16556
rect 28993 16418 29059 16421
rect 34424 16418 34484 16491
rect 28993 16416 34484 16418
rect 28993 16360 28998 16416
rect 29054 16360 34484 16416
rect 28993 16358 34484 16360
rect 28993 16355 29059 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 26734 16220 26740 16284
rect 26804 16282 26810 16284
rect 31201 16282 31267 16285
rect 26804 16280 31267 16282
rect 26804 16224 31206 16280
rect 31262 16224 31267 16280
rect 26804 16222 31267 16224
rect 26804 16220 26810 16222
rect 31201 16219 31267 16222
rect 4210 15808 4526 15809
rect 200 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1761 15738 1827 15741
rect 200 15736 1827 15738
rect 200 15680 1766 15736
rect 1822 15680 1827 15736
rect 200 15678 1827 15680
rect 200 15648 800 15678
rect 1761 15675 1827 15678
rect 38193 15738 38259 15741
rect 39200 15738 39800 15768
rect 38193 15736 39800 15738
rect 38193 15680 38198 15736
rect 38254 15680 39800 15736
rect 38193 15678 39800 15680
rect 38193 15675 38259 15678
rect 39200 15648 39800 15678
rect 31661 15602 31727 15605
rect 36302 15602 36308 15604
rect 31661 15600 36308 15602
rect 31661 15544 31666 15600
rect 31722 15544 36308 15600
rect 31661 15542 36308 15544
rect 31661 15539 31727 15542
rect 36302 15540 36308 15542
rect 36372 15540 36378 15604
rect 23289 15466 23355 15469
rect 28441 15466 28507 15469
rect 23289 15464 28507 15466
rect 23289 15408 23294 15464
rect 23350 15408 28446 15464
rect 28502 15408 28507 15464
rect 23289 15406 28507 15408
rect 23289 15403 23355 15406
rect 28441 15403 28507 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 23422 15132 23428 15196
rect 23492 15194 23498 15196
rect 23657 15194 23723 15197
rect 23492 15192 23723 15194
rect 23492 15136 23662 15192
rect 23718 15136 23723 15192
rect 23492 15134 23723 15136
rect 23492 15132 23498 15134
rect 23657 15131 23723 15134
rect 38101 15058 38167 15061
rect 39200 15058 39800 15088
rect 38101 15056 39800 15058
rect 38101 15000 38106 15056
rect 38162 15000 39800 15056
rect 38101 14998 39800 15000
rect 38101 14995 38167 14998
rect 39200 14968 39800 14998
rect 30833 14922 30899 14925
rect 31201 14922 31267 14925
rect 30833 14920 31267 14922
rect 30833 14864 30838 14920
rect 30894 14864 31206 14920
rect 31262 14864 31267 14920
rect 30833 14862 31267 14864
rect 30833 14859 30899 14862
rect 31201 14859 31267 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 200 14378 800 14408
rect 1761 14378 1827 14381
rect 200 14376 1827 14378
rect 200 14320 1766 14376
rect 1822 14320 1827 14376
rect 200 14318 1827 14320
rect 200 14288 800 14318
rect 1761 14315 1827 14318
rect 25814 14316 25820 14380
rect 25884 14378 25890 14380
rect 27705 14378 27771 14381
rect 28533 14378 28599 14381
rect 25884 14376 28599 14378
rect 25884 14320 27710 14376
rect 27766 14320 28538 14376
rect 28594 14320 28599 14376
rect 25884 14318 28599 14320
rect 25884 14316 25890 14318
rect 27705 14315 27771 14318
rect 28533 14315 28599 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 200 13698 800 13728
rect 1761 13698 1827 13701
rect 200 13696 1827 13698
rect 200 13640 1766 13696
rect 1822 13640 1827 13696
rect 200 13638 1827 13640
rect 200 13608 800 13638
rect 1761 13635 1827 13638
rect 32949 13700 33015 13701
rect 32949 13696 32996 13700
rect 33060 13698 33066 13700
rect 38193 13698 38259 13701
rect 39200 13698 39800 13728
rect 32949 13640 32954 13696
rect 32949 13636 32996 13640
rect 33060 13638 33106 13698
rect 38193 13696 39800 13698
rect 38193 13640 38198 13696
rect 38254 13640 39800 13696
rect 38193 13638 39800 13640
rect 33060 13636 33066 13638
rect 32949 13635 33015 13636
rect 38193 13635 38259 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 39800 13638
rect 34930 13567 35246 13568
rect 22001 13562 22067 13565
rect 28441 13562 28507 13565
rect 22001 13560 28507 13562
rect 22001 13504 22006 13560
rect 22062 13504 28446 13560
rect 28502 13504 28507 13560
rect 22001 13502 28507 13504
rect 22001 13499 22067 13502
rect 28441 13499 28507 13502
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 200 12338 800 12368
rect 1761 12338 1827 12341
rect 200 12336 1827 12338
rect 200 12280 1766 12336
rect 1822 12280 1827 12336
rect 200 12278 1827 12280
rect 200 12248 800 12278
rect 1761 12275 1827 12278
rect 36813 12340 36879 12341
rect 36813 12336 36860 12340
rect 36924 12338 36930 12340
rect 38193 12338 38259 12341
rect 39200 12338 39800 12368
rect 36813 12280 36818 12336
rect 36813 12276 36860 12280
rect 36924 12278 36970 12338
rect 38193 12336 39800 12338
rect 38193 12280 38198 12336
rect 38254 12280 39800 12336
rect 38193 12278 39800 12280
rect 36924 12276 36930 12278
rect 36813 12275 36879 12276
rect 38193 12275 38259 12278
rect 39200 12248 39800 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 200 10978 800 11008
rect 1669 10978 1735 10981
rect 200 10976 1735 10978
rect 200 10920 1674 10976
rect 1730 10920 1735 10976
rect 200 10918 1735 10920
rect 200 10888 800 10918
rect 1669 10915 1735 10918
rect 38193 10978 38259 10981
rect 39200 10978 39800 11008
rect 38193 10976 39800 10978
rect 38193 10920 38198 10976
rect 38254 10920 39800 10976
rect 38193 10918 39800 10920
rect 38193 10915 38259 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 39800 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1761 10298 1827 10301
rect 200 10296 1827 10298
rect 200 10240 1766 10296
rect 1822 10240 1827 10296
rect 200 10238 1827 10240
rect 200 10208 800 10238
rect 1761 10235 1827 10238
rect 38193 10298 38259 10301
rect 39200 10298 39800 10328
rect 38193 10296 39800 10298
rect 38193 10240 38198 10296
rect 38254 10240 39800 10296
rect 38193 10238 39800 10240
rect 38193 10235 38259 10238
rect 39200 10208 39800 10238
rect 22277 9890 22343 9893
rect 29729 9890 29795 9893
rect 30414 9890 30420 9892
rect 22277 9888 30420 9890
rect 22277 9832 22282 9888
rect 22338 9832 29734 9888
rect 29790 9832 30420 9888
rect 22277 9830 30420 9832
rect 22277 9827 22343 9830
rect 29729 9827 29795 9830
rect 30414 9828 30420 9830
rect 30484 9828 30490 9892
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 200 8938 800 8968
rect 1761 8938 1827 8941
rect 200 8936 1827 8938
rect 200 8880 1766 8936
rect 1822 8880 1827 8936
rect 200 8878 1827 8880
rect 200 8848 800 8878
rect 1761 8875 1827 8878
rect 38285 8938 38351 8941
rect 39200 8938 39800 8968
rect 38285 8936 39800 8938
rect 38285 8880 38290 8936
rect 38346 8880 39800 8936
rect 38285 8878 39800 8880
rect 38285 8875 38351 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 200 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 1761 7578 1827 7581
rect 200 7576 1827 7578
rect 200 7520 1766 7576
rect 1822 7520 1827 7576
rect 200 7518 1827 7520
rect 200 7488 800 7518
rect 1761 7515 1827 7518
rect 37457 7578 37523 7581
rect 39200 7578 39800 7608
rect 37457 7576 39800 7578
rect 37457 7520 37462 7576
rect 37518 7520 39800 7576
rect 37457 7518 39800 7520
rect 37457 7515 37523 7518
rect 39200 7488 39800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 200 6898 800 6928
rect 1761 6898 1827 6901
rect 200 6896 1827 6898
rect 200 6840 1766 6896
rect 1822 6840 1827 6896
rect 200 6838 1827 6840
rect 200 6808 800 6838
rect 1761 6835 1827 6838
rect 38285 6898 38351 6901
rect 39200 6898 39800 6928
rect 38285 6896 39800 6898
rect 38285 6840 38290 6896
rect 38346 6840 39800 6896
rect 38285 6838 39800 6840
rect 38285 6835 38351 6838
rect 39200 6808 39800 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 200 5538 800 5568
rect 1761 5538 1827 5541
rect 200 5536 1827 5538
rect 200 5480 1766 5536
rect 1822 5480 1827 5536
rect 200 5478 1827 5480
rect 200 5448 800 5478
rect 1761 5475 1827 5478
rect 38193 5538 38259 5541
rect 39200 5538 39800 5568
rect 38193 5536 39800 5538
rect 38193 5480 38198 5536
rect 38254 5480 39800 5536
rect 38193 5478 39800 5480
rect 38193 5475 38259 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 39800 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 200 4178 800 4208
rect 1761 4178 1827 4181
rect 200 4176 1827 4178
rect 200 4120 1766 4176
rect 1822 4120 1827 4176
rect 200 4118 1827 4120
rect 200 4088 800 4118
rect 1761 4115 1827 4118
rect 37457 4178 37523 4181
rect 39200 4178 39800 4208
rect 37457 4176 39800 4178
rect 37457 4120 37462 4176
rect 37518 4120 39800 4176
rect 37457 4118 39800 4120
rect 37457 4115 37523 4118
rect 39200 4088 39800 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 200 3498 800 3528
rect 1761 3498 1827 3501
rect 200 3496 1827 3498
rect 200 3440 1766 3496
rect 1822 3440 1827 3496
rect 200 3438 1827 3440
rect 200 3408 800 3438
rect 1761 3435 1827 3438
rect 38193 3498 38259 3501
rect 39200 3498 39800 3528
rect 38193 3496 39800 3498
rect 38193 3440 38198 3496
rect 38254 3440 39800 3496
rect 38193 3438 39800 3440
rect 38193 3435 38259 3438
rect 39200 3408 39800 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 200 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 2773 2138 2839 2141
rect 200 2136 2839 2138
rect 200 2080 2778 2136
rect 2834 2080 2839 2136
rect 200 2078 2839 2080
rect 200 2048 800 2078
rect 2773 2075 2839 2078
rect 36813 2138 36879 2141
rect 39200 2138 39800 2168
rect 36813 2136 39800 2138
rect 36813 2080 36818 2136
rect 36874 2080 39800 2136
rect 36813 2078 39800 2080
rect 36813 2075 36879 2078
rect 39200 2048 39800 2078
rect 200 778 800 808
rect 2865 778 2931 781
rect 200 776 2931 778
rect 200 720 2870 776
rect 2926 720 2931 776
rect 200 718 2931 720
rect 200 688 800 718
rect 2865 715 2931 718
rect 37733 778 37799 781
rect 39200 778 39800 808
rect 37733 776 39800 778
rect 37733 720 37738 776
rect 37794 720 39800 776
rect 37733 718 39800 720
rect 37733 715 37799 718
rect 39200 688 39800 718
rect 37181 98 37247 101
rect 39200 98 39800 128
rect 37181 96 39800 98
rect 37181 40 37186 96
rect 37242 40 39800 96
rect 37181 38 39800 40
rect 37181 35 37247 38
rect 39200 8 39800 38
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 16988 36756 17052 36820
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 22140 36000 22204 36004
rect 22140 35944 22154 36000
rect 22154 35944 22204 36000
rect 22140 35940 22204 35944
rect 26188 36000 26252 36004
rect 26188 35944 26238 36000
rect 26238 35944 26252 36000
rect 26188 35940 26252 35944
rect 29316 35940 29380 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 28764 34776 28828 34780
rect 28764 34720 28778 34776
rect 28778 34720 28828 34776
rect 28764 34716 28828 34720
rect 28580 34640 28644 34644
rect 28580 34584 28594 34640
rect 28594 34584 28644 34640
rect 28580 34580 28644 34584
rect 31340 34580 31404 34644
rect 35756 34580 35820 34644
rect 30972 34444 31036 34508
rect 32996 34308 33060 34372
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 28028 33220 28092 33284
rect 29868 33280 29932 33284
rect 29868 33224 29882 33280
rect 29882 33224 29932 33280
rect 29868 33220 29932 33224
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 28396 32872 28460 32876
rect 28396 32816 28446 32872
rect 28446 32816 28460 32872
rect 28396 32812 28460 32816
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 36860 31724 36924 31788
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 25820 31180 25884 31244
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 26004 30500 26068 30564
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 12940 30364 13004 30428
rect 34468 30092 34532 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 12940 27916 13004 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 25452 27644 25516 27708
rect 26004 27704 26068 27708
rect 26004 27648 26018 27704
rect 26018 27648 26068 27704
rect 26004 27644 26068 27648
rect 33180 27644 33244 27708
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 23980 26828 24044 26892
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 26740 26284 26804 26348
rect 32444 26148 32508 26212
rect 36676 26148 36740 26212
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 30236 25196 30300 25260
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 21404 24788 21468 24852
rect 27476 24788 27540 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 12940 23700 13004 23764
rect 16988 23428 17052 23492
rect 21220 23428 21284 23492
rect 30420 23488 30484 23492
rect 30420 23432 30434 23488
rect 30434 23432 30484 23488
rect 30420 23428 30484 23432
rect 33732 23428 33796 23492
rect 36308 23488 36372 23492
rect 36308 23432 36358 23488
rect 36358 23432 36372 23488
rect 36308 23428 36372 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 30604 23292 30668 23356
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 30604 22204 30668 22268
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 21220 21176 21284 21180
rect 21220 21120 21234 21176
rect 21234 21120 21284 21176
rect 21220 21116 21284 21120
rect 21404 20980 21468 21044
rect 34652 20980 34716 21044
rect 23428 20844 23492 20908
rect 25820 20904 25884 20908
rect 25820 20848 25834 20904
rect 25834 20848 25884 20904
rect 25820 20844 25884 20848
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 30604 20572 30668 20636
rect 28580 20436 28644 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 27476 20028 27540 20092
rect 36676 20088 36740 20092
rect 36676 20032 36726 20088
rect 36726 20032 36740 20088
rect 36676 20028 36740 20032
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 34468 19484 34532 19548
rect 33180 19348 33244 19412
rect 34468 19348 34532 19412
rect 28028 19272 28092 19276
rect 28028 19216 28042 19272
rect 28042 19216 28092 19272
rect 28028 19212 28092 19216
rect 28764 19212 28828 19276
rect 30236 19212 30300 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 22140 18940 22204 19004
rect 35756 18804 35820 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 25452 18396 25516 18460
rect 26188 18396 26252 18460
rect 31340 18124 31404 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 23980 17852 24044 17916
rect 29868 17852 29932 17916
rect 32444 17852 32508 17916
rect 34468 17716 34532 17780
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 29316 17308 29380 17372
rect 12940 17172 13004 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 28396 16764 28460 16828
rect 30972 16492 31036 16556
rect 33732 16492 33796 16556
rect 34652 16492 34716 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 26740 16220 26804 16284
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 36308 15540 36372 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 23428 15132 23492 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 25820 14316 25884 14380
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 32996 13696 33060 13700
rect 32996 13640 33010 13696
rect 33010 13640 33060 13696
rect 32996 13636 33060 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 36860 12336 36924 12340
rect 36860 12280 36874 12336
rect 36874 12280 36924 12336
rect 36860 12276 36924 12280
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 30420 9828 30484 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 16987 36820 17053 36821
rect 16987 36756 16988 36820
rect 17052 36756 17053 36820
rect 16987 36755 17053 36756
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 12939 30428 13005 30429
rect 12939 30364 12940 30428
rect 13004 30364 13005 30428
rect 12939 30363 13005 30364
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 12942 27981 13002 30363
rect 12939 27980 13005 27981
rect 12939 27916 12940 27980
rect 13004 27916 13005 27980
rect 12939 27915 13005 27916
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 12942 23765 13002 27915
rect 12939 23764 13005 23765
rect 12939 23700 12940 23764
rect 13004 23700 13005 23764
rect 12939 23699 13005 23700
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 12942 17237 13002 23699
rect 16990 23493 17050 36755
rect 19568 35936 19888 36960
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 22139 36004 22205 36005
rect 22139 35940 22140 36004
rect 22204 35940 22205 36004
rect 22139 35939 22205 35940
rect 26187 36004 26253 36005
rect 26187 35940 26188 36004
rect 26252 35940 26253 36004
rect 26187 35939 26253 35940
rect 29315 36004 29381 36005
rect 29315 35940 29316 36004
rect 29380 35940 29381 36004
rect 29315 35939 29381 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 21403 24852 21469 24853
rect 21403 24788 21404 24852
rect 21468 24788 21469 24852
rect 21403 24787 21469 24788
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 16987 23492 17053 23493
rect 16987 23428 16988 23492
rect 17052 23428 17053 23492
rect 16987 23427 17053 23428
rect 19568 22880 19888 23904
rect 21219 23492 21285 23493
rect 21219 23428 21220 23492
rect 21284 23428 21285 23492
rect 21219 23427 21285 23428
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 21222 21181 21282 23427
rect 21219 21180 21285 21181
rect 21219 21116 21220 21180
rect 21284 21116 21285 21180
rect 21219 21115 21285 21116
rect 21406 21045 21466 24787
rect 21403 21044 21469 21045
rect 21403 20980 21404 21044
rect 21468 20980 21469 21044
rect 21403 20979 21469 20980
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 22142 19005 22202 35939
rect 25819 31244 25885 31245
rect 25819 31180 25820 31244
rect 25884 31180 25885 31244
rect 25819 31179 25885 31180
rect 25451 27708 25517 27709
rect 25451 27644 25452 27708
rect 25516 27644 25517 27708
rect 25451 27643 25517 27644
rect 23979 26892 24045 26893
rect 23979 26828 23980 26892
rect 24044 26828 24045 26892
rect 23979 26827 24045 26828
rect 23427 20908 23493 20909
rect 23427 20844 23428 20908
rect 23492 20844 23493 20908
rect 23427 20843 23493 20844
rect 22139 19004 22205 19005
rect 22139 18940 22140 19004
rect 22204 18940 22205 19004
rect 22139 18939 22205 18940
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 12939 17236 13005 17237
rect 12939 17172 12940 17236
rect 13004 17172 13005 17236
rect 12939 17171 13005 17172
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 23430 15197 23490 20843
rect 23982 17917 24042 26827
rect 25454 18461 25514 27643
rect 25822 20909 25882 31179
rect 26003 30564 26069 30565
rect 26003 30500 26004 30564
rect 26068 30500 26069 30564
rect 26003 30499 26069 30500
rect 26006 27709 26066 30499
rect 26003 27708 26069 27709
rect 26003 27644 26004 27708
rect 26068 27644 26069 27708
rect 26003 27643 26069 27644
rect 25819 20908 25885 20909
rect 25819 20844 25820 20908
rect 25884 20844 25885 20908
rect 25819 20843 25885 20844
rect 25451 18460 25517 18461
rect 25451 18396 25452 18460
rect 25516 18396 25517 18460
rect 25451 18395 25517 18396
rect 23979 17916 24045 17917
rect 23979 17852 23980 17916
rect 24044 17852 24045 17916
rect 23979 17851 24045 17852
rect 23427 15196 23493 15197
rect 23427 15132 23428 15196
rect 23492 15132 23493 15196
rect 23427 15131 23493 15132
rect 25822 14381 25882 20843
rect 26190 18461 26250 35939
rect 28763 34780 28829 34781
rect 28763 34716 28764 34780
rect 28828 34716 28829 34780
rect 28763 34715 28829 34716
rect 28579 34644 28645 34645
rect 28579 34580 28580 34644
rect 28644 34580 28645 34644
rect 28579 34579 28645 34580
rect 28027 33284 28093 33285
rect 28027 33220 28028 33284
rect 28092 33220 28093 33284
rect 28027 33219 28093 33220
rect 26739 26348 26805 26349
rect 26739 26284 26740 26348
rect 26804 26284 26805 26348
rect 26739 26283 26805 26284
rect 26187 18460 26253 18461
rect 26187 18396 26188 18460
rect 26252 18396 26253 18460
rect 26187 18395 26253 18396
rect 26742 16285 26802 26283
rect 27475 24852 27541 24853
rect 27475 24788 27476 24852
rect 27540 24788 27541 24852
rect 27475 24787 27541 24788
rect 27478 20093 27538 24787
rect 27475 20092 27541 20093
rect 27475 20028 27476 20092
rect 27540 20028 27541 20092
rect 27475 20027 27541 20028
rect 28030 19277 28090 33219
rect 28395 32876 28461 32877
rect 28395 32812 28396 32876
rect 28460 32812 28461 32876
rect 28395 32811 28461 32812
rect 28027 19276 28093 19277
rect 28027 19212 28028 19276
rect 28092 19212 28093 19276
rect 28027 19211 28093 19212
rect 28398 16829 28458 32811
rect 28582 20501 28642 34579
rect 28579 20500 28645 20501
rect 28579 20436 28580 20500
rect 28644 20436 28645 20500
rect 28579 20435 28645 20436
rect 28766 19277 28826 34715
rect 28763 19276 28829 19277
rect 28763 19212 28764 19276
rect 28828 19212 28829 19276
rect 28763 19211 28829 19212
rect 29318 17373 29378 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 31339 34644 31405 34645
rect 31339 34580 31340 34644
rect 31404 34580 31405 34644
rect 31339 34579 31405 34580
rect 30971 34508 31037 34509
rect 30971 34444 30972 34508
rect 31036 34444 31037 34508
rect 30971 34443 31037 34444
rect 29867 33284 29933 33285
rect 29867 33220 29868 33284
rect 29932 33220 29933 33284
rect 29867 33219 29933 33220
rect 29870 17917 29930 33219
rect 30235 25260 30301 25261
rect 30235 25196 30236 25260
rect 30300 25196 30301 25260
rect 30235 25195 30301 25196
rect 30238 19277 30298 25195
rect 30419 23492 30485 23493
rect 30419 23428 30420 23492
rect 30484 23428 30485 23492
rect 30419 23427 30485 23428
rect 30235 19276 30301 19277
rect 30235 19212 30236 19276
rect 30300 19212 30301 19276
rect 30235 19211 30301 19212
rect 29867 17916 29933 17917
rect 29867 17852 29868 17916
rect 29932 17852 29933 17916
rect 29867 17851 29933 17852
rect 29315 17372 29381 17373
rect 29315 17308 29316 17372
rect 29380 17308 29381 17372
rect 29315 17307 29381 17308
rect 28395 16828 28461 16829
rect 28395 16764 28396 16828
rect 28460 16764 28461 16828
rect 28395 16763 28461 16764
rect 26739 16284 26805 16285
rect 26739 16220 26740 16284
rect 26804 16220 26805 16284
rect 26739 16219 26805 16220
rect 25819 14380 25885 14381
rect 25819 14316 25820 14380
rect 25884 14316 25885 14380
rect 25819 14315 25885 14316
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 30422 9893 30482 23427
rect 30603 23356 30669 23357
rect 30603 23292 30604 23356
rect 30668 23292 30669 23356
rect 30603 23291 30669 23292
rect 30606 22269 30666 23291
rect 30603 22268 30669 22269
rect 30603 22204 30604 22268
rect 30668 22204 30669 22268
rect 30603 22203 30669 22204
rect 30606 20637 30666 22203
rect 30603 20636 30669 20637
rect 30603 20572 30604 20636
rect 30668 20572 30669 20636
rect 30603 20571 30669 20572
rect 30974 16557 31034 34443
rect 31342 18189 31402 34579
rect 32995 34372 33061 34373
rect 32995 34308 32996 34372
rect 33060 34308 33061 34372
rect 32995 34307 33061 34308
rect 32443 26212 32509 26213
rect 32443 26148 32444 26212
rect 32508 26148 32509 26212
rect 32443 26147 32509 26148
rect 31339 18188 31405 18189
rect 31339 18124 31340 18188
rect 31404 18124 31405 18188
rect 31339 18123 31405 18124
rect 32446 17917 32506 26147
rect 32443 17916 32509 17917
rect 32443 17852 32444 17916
rect 32508 17852 32509 17916
rect 32443 17851 32509 17852
rect 30971 16556 31037 16557
rect 30971 16492 30972 16556
rect 31036 16492 31037 16556
rect 30971 16491 31037 16492
rect 32998 13701 33058 34307
rect 34928 34304 35248 35328
rect 35755 34644 35821 34645
rect 35755 34580 35756 34644
rect 35820 34580 35821 34644
rect 35755 34579 35821 34580
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34467 30156 34533 30157
rect 34467 30092 34468 30156
rect 34532 30092 34533 30156
rect 34467 30091 34533 30092
rect 33179 27708 33245 27709
rect 33179 27644 33180 27708
rect 33244 27644 33245 27708
rect 33179 27643 33245 27644
rect 33182 19413 33242 27643
rect 33731 23492 33797 23493
rect 33731 23428 33732 23492
rect 33796 23428 33797 23492
rect 33731 23427 33797 23428
rect 33179 19412 33245 19413
rect 33179 19348 33180 19412
rect 33244 19348 33245 19412
rect 33179 19347 33245 19348
rect 33734 16557 33794 23427
rect 34470 19549 34530 30091
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34651 21044 34717 21045
rect 34651 20980 34652 21044
rect 34716 20980 34717 21044
rect 34651 20979 34717 20980
rect 34467 19548 34533 19549
rect 34467 19484 34468 19548
rect 34532 19484 34533 19548
rect 34467 19483 34533 19484
rect 34467 19412 34533 19413
rect 34467 19348 34468 19412
rect 34532 19348 34533 19412
rect 34467 19347 34533 19348
rect 34470 17781 34530 19347
rect 34467 17780 34533 17781
rect 34467 17716 34468 17780
rect 34532 17716 34533 17780
rect 34467 17715 34533 17716
rect 34654 16557 34714 20979
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 35758 18869 35818 34579
rect 36859 31788 36925 31789
rect 36859 31724 36860 31788
rect 36924 31724 36925 31788
rect 36859 31723 36925 31724
rect 36675 26212 36741 26213
rect 36675 26148 36676 26212
rect 36740 26148 36741 26212
rect 36675 26147 36741 26148
rect 36307 23492 36373 23493
rect 36307 23428 36308 23492
rect 36372 23428 36373 23492
rect 36307 23427 36373 23428
rect 35755 18868 35821 18869
rect 35755 18804 35756 18868
rect 35820 18804 35821 18868
rect 35755 18803 35821 18804
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 33731 16556 33797 16557
rect 33731 16492 33732 16556
rect 33796 16492 33797 16556
rect 33731 16491 33797 16492
rect 34651 16556 34717 16557
rect 34651 16492 34652 16556
rect 34716 16492 34717 16556
rect 34651 16491 34717 16492
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 36310 15605 36370 23427
rect 36678 20093 36738 26147
rect 36675 20092 36741 20093
rect 36675 20028 36676 20092
rect 36740 20028 36741 20092
rect 36675 20027 36741 20028
rect 36307 15604 36373 15605
rect 36307 15540 36308 15604
rect 36372 15540 36373 15604
rect 36307 15539 36373 15540
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 32995 13700 33061 13701
rect 32995 13636 32996 13700
rect 33060 13636 33061 13700
rect 32995 13635 33061 13636
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 36862 12341 36922 31723
rect 36859 12340 36925 12341
rect 36859 12276 36860 12340
rect 36924 12276 36925 12340
rect 36859 12275 36925 12276
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 30419 9892 30485 9893
rect 30419 9828 30420 9892
rect 30484 9828 30485 9892
rect 30419 9827 30485 9828
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31832 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 37628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1667941163
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1667941163
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1667941163
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1667941163
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1667941163
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1667941163
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 7544 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1667941163
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1667941163
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1667941163
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1667941163
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1667941163
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1667941163
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1667941163
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1667941163
transform 1 0 15824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1667941163
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1667941163
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1667941163
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_230
timestamp 1667941163
transform 1 0 22264 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_238
timestamp 1667941163
transform 1 0 23000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1667941163
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_258
timestamp 1667941163
transform 1 0 24840 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_266
timestamp 1667941163
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1667941163
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1667941163
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_294
timestamp 1667941163
transform 1 0 28152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1667941163
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_315
timestamp 1667941163
transform 1 0 30084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_323
timestamp 1667941163
transform 1 0 30820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1667941163
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1667941163
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_371
timestamp 1667941163
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1667941163
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1667941163
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_399
timestamp 1667941163
transform 1 0 37812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1667941163
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1667941163
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1667941163
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23
timestamp 1667941163
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1667941163
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1667941163
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp 1667941163
transform 1 0 12972 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_133
timestamp 1667941163
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1667941163
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1667941163
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1667941163
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_174
timestamp 1667941163
transform 1 0 17112 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_186
timestamp 1667941163
transform 1 0 18216 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_198
timestamp 1667941163
transform 1 0 19320 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_210
timestamp 1667941163
transform 1 0 20424 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1667941163
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1667941163
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_322
timestamp 1667941163
transform 1 0 30728 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1667941163
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_369
timestamp 1667941163
transform 1 0 35052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1667941163
transform 1 0 35512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_381
timestamp 1667941163
transform 1 0 36156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1667941163
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_9
timestamp 1667941163
transform 1 0 1932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1667941163
transform 1 0 3036 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_385
timestamp 1667941163
transform 1 0 36524 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_390
timestamp 1667941163
transform 1 0 36984 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_397
timestamp 1667941163
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_405
timestamp 1667941163
transform 1 0 38364 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_402
timestamp 1667941163
transform 1 0 38088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_406
timestamp 1667941163
transform 1 0 38456 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1667941163
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_13
timestamp 1667941163
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1667941163
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_405
timestamp 1667941163
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_231
timestamp 1667941163
transform 1 0 22356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_236
timestamp 1667941163
transform 1 0 22816 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_244
timestamp 1667941163
transform 1 0 23552 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1667941163
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1667941163
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1667941163
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_310
timestamp 1667941163
transform 1 0 29624 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_322
timestamp 1667941163
transform 1 0 30728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1667941163
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_8
timestamp 1667941163
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1667941163
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_271
timestamp 1667941163
transform 1 0 26036 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_275
timestamp 1667941163
transform 1 0 26404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_287
timestamp 1667941163
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_299
timestamp 1667941163
transform 1 0 28612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_399
timestamp 1667941163
transform 1 0 37812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_405
timestamp 1667941163
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_153
timestamp 1667941163
transform 1 0 15180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1667941163
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_253
timestamp 1667941163
transform 1 0 24380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_257
timestamp 1667941163
transform 1 0 24748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1667941163
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1667941163
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_320
timestamp 1667941163
transform 1 0 30544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1667941163
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_90
timestamp 1667941163
transform 1 0 9384 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_102
timestamp 1667941163
transform 1 0 10488 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_114
timestamp 1667941163
transform 1 0 11592 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_126
timestamp 1667941163
transform 1 0 12696 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1667941163
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_241
timestamp 1667941163
transform 1 0 23276 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1667941163
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_258
timestamp 1667941163
transform 1 0 24840 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_270
timestamp 1667941163
transform 1 0 25944 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_282
timestamp 1667941163
transform 1 0 27048 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1667941163
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1667941163
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_314
timestamp 1667941163
transform 1 0 29992 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_331
timestamp 1667941163
transform 1 0 31556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_343
timestamp 1667941163
transform 1 0 32660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_355
timestamp 1667941163
transform 1 0 33764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_8
timestamp 1667941163
transform 1 0 1840 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1667941163
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_32
timestamp 1667941163
transform 1 0 4048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1667941163
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_211
timestamp 1667941163
transform 1 0 20516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1667941163
transform 1 0 23460 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_247
timestamp 1667941163
transform 1 0 23828 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_259
timestamp 1667941163
transform 1 0 24932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_267
timestamp 1667941163
transform 1 0 25668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1667941163
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_401
timestamp 1667941163
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_8
timestamp 1667941163
transform 1 0 1840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1667941163
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1667941163
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_227
timestamp 1667941163
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_239
timestamp 1667941163
transform 1 0 23092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1667941163
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_293
timestamp 1667941163
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1667941163
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_327
timestamp 1667941163
transform 1 0 31188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_332
timestamp 1667941163
transform 1 0 31648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_336
timestamp 1667941163
transform 1 0 32016 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_341
timestamp 1667941163
transform 1 0 32476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_353
timestamp 1667941163
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_361
timestamp 1667941163
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1667941163
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1667941163
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1667941163
transform 1 0 10580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1667941163
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_236
timestamp 1667941163
transform 1 0 22816 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_248
timestamp 1667941163
transform 1 0 23920 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_260
timestamp 1667941163
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_272
timestamp 1667941163
transform 1 0 26128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1667941163
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_296
timestamp 1667941163
transform 1 0 28336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_313
timestamp 1667941163
transform 1 0 29900 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_318
timestamp 1667941163
transform 1 0 30360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_330
timestamp 1667941163
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_401
timestamp 1667941163
transform 1 0 37996 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_9
timestamp 1667941163
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1667941163
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_151
timestamp 1667941163
transform 1 0 14996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1667941163
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1667941163
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1667941163
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_205
timestamp 1667941163
transform 1 0 19964 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_210
timestamp 1667941163
transform 1 0 20424 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_222
timestamp 1667941163
transform 1 0 21528 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_241
timestamp 1667941163
transform 1 0 23276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_249
timestamp 1667941163
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1667941163
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_276
timestamp 1667941163
transform 1 0 26496 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_282
timestamp 1667941163
transform 1 0 27048 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_286
timestamp 1667941163
transform 1 0 27416 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_298
timestamp 1667941163
transform 1 0 28520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1667941163
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_313
timestamp 1667941163
transform 1 0 29900 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_323
timestamp 1667941163
transform 1 0 30820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_335
timestamp 1667941163
transform 1 0 31924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_343
timestamp 1667941163
transform 1 0 32660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_347
timestamp 1667941163
transform 1 0 33028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1667941163
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_395
timestamp 1667941163
transform 1 0 37444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_399
timestamp 1667941163
transform 1 0 37812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1667941163
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1667941163
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1667941163
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1667941163
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1667941163
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp 1667941163
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 1667941163
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1667941163
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1667941163
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1667941163
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1667941163
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_180
timestamp 1667941163
transform 1 0 17664 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1667941163
transform 1 0 18768 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1667941163
transform 1 0 19504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_233
timestamp 1667941163
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_250
timestamp 1667941163
transform 1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_308
timestamp 1667941163
transform 1 0 29440 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_320
timestamp 1667941163
transform 1 0 30544 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1667941163
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_397
timestamp 1667941163
transform 1 0 37628 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_401
timestamp 1667941163
transform 1 0 37996 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1667941163
transform 1 0 1932 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_14
timestamp 1667941163
transform 1 0 2392 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1667941163
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1667941163
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_167
timestamp 1667941163
transform 1 0 16468 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_179
timestamp 1667941163
transform 1 0 17572 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_184
timestamp 1667941163
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_224
timestamp 1667941163
transform 1 0 21712 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_263
timestamp 1667941163
transform 1 0 25300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_275
timestamp 1667941163
transform 1 0 26404 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_283
timestamp 1667941163
transform 1 0 27140 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_287
timestamp 1667941163
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_299
timestamp 1667941163
transform 1 0 28612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_317
timestamp 1667941163
transform 1 0 30268 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_385
timestamp 1667941163
transform 1 0 36524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_390
timestamp 1667941163
transform 1 0 36984 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_397
timestamp 1667941163
transform 1 0 37628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_405
timestamp 1667941163
transform 1 0 38364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1667941163
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1667941163
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_85
timestamp 1667941163
transform 1 0 8924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_89
timestamp 1667941163
transform 1 0 9292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1667941163
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1667941163
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_145
timestamp 1667941163
transform 1 0 14444 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_208
timestamp 1667941163
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1667941163
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_232
timestamp 1667941163
transform 1 0 22448 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_244
timestamp 1667941163
transform 1 0 23552 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_253
timestamp 1667941163
transform 1 0 24380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_265
timestamp 1667941163
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1667941163
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_292
timestamp 1667941163
transform 1 0 27968 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_300
timestamp 1667941163
transform 1 0 28704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_310
timestamp 1667941163
transform 1 0 29624 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_382
timestamp 1667941163
transform 1 0 36248 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_386
timestamp 1667941163
transform 1 0 36616 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1667941163
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_9
timestamp 1667941163
transform 1 0 1932 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1667941163
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_57
timestamp 1667941163
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_61
timestamp 1667941163
transform 1 0 6716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1667941163
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_71
timestamp 1667941163
transform 1 0 7636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_95
timestamp 1667941163
transform 1 0 9844 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_103
timestamp 1667941163
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_107
timestamp 1667941163
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_119
timestamp 1667941163
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1667941163
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_159
timestamp 1667941163
transform 1 0 15732 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_163
timestamp 1667941163
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1667941163
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1667941163
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_207
timestamp 1667941163
transform 1 0 20148 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1667941163
transform 1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_225
timestamp 1667941163
transform 1 0 21804 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_232
timestamp 1667941163
transform 1 0 22448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1667941163
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1667941163
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_316
timestamp 1667941163
transform 1 0 30176 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_320
timestamp 1667941163
transform 1 0 30544 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_324
timestamp 1667941163
transform 1 0 30912 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_331
timestamp 1667941163
transform 1 0 31556 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_343
timestamp 1667941163
transform 1 0 32660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_355
timestamp 1667941163
transform 1 0 33764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_370
timestamp 1667941163
transform 1 0 35144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_385
timestamp 1667941163
transform 1 0 36524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_391
timestamp 1667941163
transform 1 0 37076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_404
timestamp 1667941163
transform 1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_64
timestamp 1667941163
transform 1 0 6992 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_76
timestamp 1667941163
transform 1 0 8096 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_88
timestamp 1667941163
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_100
timestamp 1667941163
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_121
timestamp 1667941163
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_127
timestamp 1667941163
transform 1 0 12788 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_139
timestamp 1667941163
transform 1 0 13892 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_151
timestamp 1667941163
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1667941163
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_174
timestamp 1667941163
transform 1 0 17112 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_191
timestamp 1667941163
transform 1 0 18676 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_203
timestamp 1667941163
transform 1 0 19780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1667941163
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1667941163
transform 1 0 22264 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1667941163
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_261
timestamp 1667941163
transform 1 0 25116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_271
timestamp 1667941163
transform 1 0 26036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1667941163
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_312
timestamp 1667941163
transform 1 0 29808 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_320
timestamp 1667941163
transform 1 0 30544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1667941163
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_342
timestamp 1667941163
transform 1 0 32568 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_372
timestamp 1667941163
transform 1 0 35328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_376
timestamp 1667941163
transform 1 0 35696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_380
timestamp 1667941163
transform 1 0 36064 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1667941163
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_397
timestamp 1667941163
transform 1 0 37628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_401
timestamp 1667941163
transform 1 0 37996 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_37
timestamp 1667941163
transform 1 0 4508 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_43
timestamp 1667941163
transform 1 0 5060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_55
timestamp 1667941163
transform 1 0 6164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_67
timestamp 1667941163
transform 1 0 7268 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1667941163
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_146
timestamp 1667941163
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_158
timestamp 1667941163
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_170
timestamp 1667941163
transform 1 0 16744 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_182
timestamp 1667941163
transform 1 0 17848 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1667941163
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_212
timestamp 1667941163
transform 1 0 20608 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_224
timestamp 1667941163
transform 1 0 21712 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1667941163
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1667941163
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1667941163
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1667941163
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1667941163
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1667941163
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_340
timestamp 1667941163
transform 1 0 32384 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_348
timestamp 1667941163
transform 1 0 33120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_352
timestamp 1667941163
transform 1 0 33488 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1667941163
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_376
timestamp 1667941163
transform 1 0 35696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_383
timestamp 1667941163
transform 1 0 36340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_392
timestamp 1667941163
transform 1 0 37168 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_396
timestamp 1667941163
transform 1 0 37536 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_400
timestamp 1667941163
transform 1 0 37904 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1667941163
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_9
timestamp 1667941163
transform 1 0 1932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_21
timestamp 1667941163
transform 1 0 3036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_29
timestamp 1667941163
transform 1 0 3772 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1667941163
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1667941163
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1667941163
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1667941163
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_123
timestamp 1667941163
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_135
timestamp 1667941163
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_147
timestamp 1667941163
transform 1 0 14628 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_152
timestamp 1667941163
transform 1 0 15088 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1667941163
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_194
timestamp 1667941163
transform 1 0 18952 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1667941163
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1667941163
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_235
timestamp 1667941163
transform 1 0 22724 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_252
timestamp 1667941163
transform 1 0 24288 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_267
timestamp 1667941163
transform 1 0 25668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1667941163
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_296
timestamp 1667941163
transform 1 0 28336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_312
timestamp 1667941163
transform 1 0 29808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_324
timestamp 1667941163
transform 1 0 30912 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1667941163
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1667941163
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_345
timestamp 1667941163
transform 1 0 32844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_352
timestamp 1667941163
transform 1 0 33488 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_374
timestamp 1667941163
transform 1 0 35512 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1667941163
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_103
timestamp 1667941163
transform 1 0 10580 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_117
timestamp 1667941163
transform 1 0 11868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1667941163
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1667941163
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1667941163
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_151
timestamp 1667941163
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1667941163
transform 1 0 16100 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_184
timestamp 1667941163
transform 1 0 18032 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_208
timestamp 1667941163
transform 1 0 20240 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_220
timestamp 1667941163
transform 1 0 21344 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_225
timestamp 1667941163
transform 1 0 21804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_233
timestamp 1667941163
transform 1 0 22540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1667941163
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1667941163
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_258
timestamp 1667941163
transform 1 0 24840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1667941163
transform 1 0 25944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_282
timestamp 1667941163
transform 1 0 27048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_290
timestamp 1667941163
transform 1 0 27784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1667941163
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_319
timestamp 1667941163
transform 1 0 30452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_335
timestamp 1667941163
transform 1 0 31924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_342
timestamp 1667941163
transform 1 0 32568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_349
timestamp 1667941163
transform 1 0 33212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_357
timestamp 1667941163
transform 1 0 33948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1667941163
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_370
timestamp 1667941163
transform 1 0 35144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_384
timestamp 1667941163
transform 1 0 36432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_388
timestamp 1667941163
transform 1 0 36800 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_398
timestamp 1667941163
transform 1 0 37720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_405
timestamp 1667941163
transform 1 0 38364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_9
timestamp 1667941163
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1667941163
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1667941163
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1667941163
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1667941163
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_90
timestamp 1667941163
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1667941163
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1667941163
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_128
timestamp 1667941163
transform 1 0 12880 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_140
timestamp 1667941163
transform 1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_151
timestamp 1667941163
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1667941163
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_177
timestamp 1667941163
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_189
timestamp 1667941163
transform 1 0 18492 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_196
timestamp 1667941163
transform 1 0 19136 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1667941163
transform 1 0 19872 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_213
timestamp 1667941163
transform 1 0 20700 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1667941163
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1667941163
transform 1 0 23184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_247
timestamp 1667941163
transform 1 0 23828 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1667941163
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_302
timestamp 1667941163
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_309
timestamp 1667941163
transform 1 0 29532 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_318
timestamp 1667941163
transform 1 0 30360 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_324
timestamp 1667941163
transform 1 0 30912 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1667941163
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_343
timestamp 1667941163
transform 1 0 32660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_358
timestamp 1667941163
transform 1 0 34040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_362
timestamp 1667941163
transform 1 0 34408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_366
timestamp 1667941163
transform 1 0 34776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_374
timestamp 1667941163
transform 1 0 35512 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1667941163
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_8
timestamp 1667941163
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_20
timestamp 1667941163
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_90
timestamp 1667941163
transform 1 0 9384 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_102
timestamp 1667941163
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_114
timestamp 1667941163
transform 1 0 11592 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_120
timestamp 1667941163
transform 1 0 12144 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 1667941163
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1667941163
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1667941163
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1667941163
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_182
timestamp 1667941163
transform 1 0 17848 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1667941163
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1667941163
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_217
timestamp 1667941163
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1667941163
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_241
timestamp 1667941163
transform 1 0 23276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1667941163
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_258
timestamp 1667941163
transform 1 0 24840 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_270
timestamp 1667941163
transform 1 0 25944 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_282
timestamp 1667941163
transform 1 0 27048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1667941163
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1667941163
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_314
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_327
timestamp 1667941163
transform 1 0 31188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_334
timestamp 1667941163
transform 1 0 31832 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_342
timestamp 1667941163
transform 1 0 32568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_351
timestamp 1667941163
transform 1 0 33396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1667941163
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_370
timestamp 1667941163
transform 1 0 35144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_376
timestamp 1667941163
transform 1 0 35696 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_380
timestamp 1667941163
transform 1 0 36064 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1667941163
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_400
timestamp 1667941163
transform 1 0 37904 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1667941163
transform 1 0 38456 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1667941163
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_90
timestamp 1667941163
transform 1 0 9384 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1667941163
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1667941163
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1667941163
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_138
timestamp 1667941163
transform 1 0 13800 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_151
timestamp 1667941163
transform 1 0 14996 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1667941163
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_175
timestamp 1667941163
transform 1 0 17204 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_187
timestamp 1667941163
transform 1 0 18308 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_199
timestamp 1667941163
transform 1 0 19412 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_209
timestamp 1667941163
transform 1 0 20332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1667941163
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_232
timestamp 1667941163
transform 1 0 22448 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1667941163
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_250
timestamp 1667941163
transform 1 0 24104 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1667941163
transform 1 0 24840 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_263
timestamp 1667941163
transform 1 0 25300 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_286
timestamp 1667941163
transform 1 0 27416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_294
timestamp 1667941163
transform 1 0 28152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_304
timestamp 1667941163
transform 1 0 29072 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_311
timestamp 1667941163
transform 1 0 29716 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_319
timestamp 1667941163
transform 1 0 30452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1667941163
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_342
timestamp 1667941163
transform 1 0 32568 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_357
timestamp 1667941163
transform 1 0 33948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1667941163
transform 1 0 34868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1667941163
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_381
timestamp 1667941163
transform 1 0 36156 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1667941163
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_59
timestamp 1667941163
transform 1 0 6532 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_63
timestamp 1667941163
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1667941163
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_112
timestamp 1667941163
transform 1 0 11408 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_124
timestamp 1667941163
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1667941163
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_162
timestamp 1667941163
transform 1 0 16008 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_174
timestamp 1667941163
transform 1 0 17112 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1667941163
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1667941163
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_214
timestamp 1667941163
transform 1 0 20792 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_226
timestamp 1667941163
transform 1 0 21896 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_258
timestamp 1667941163
transform 1 0 24840 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_264
timestamp 1667941163
transform 1 0 25392 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_268
timestamp 1667941163
transform 1 0 25760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_275
timestamp 1667941163
transform 1 0 26404 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_283
timestamp 1667941163
transform 1 0 27140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_292
timestamp 1667941163
transform 1 0 27968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1667941163
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1667941163
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_321
timestamp 1667941163
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_328
timestamp 1667941163
transform 1 0 31280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_335
timestamp 1667941163
transform 1 0 31924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_342
timestamp 1667941163
transform 1 0 32568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_349
timestamp 1667941163
transform 1 0 33212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1667941163
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1667941163
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 1667941163
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_381
timestamp 1667941163
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_391
timestamp 1667941163
transform 1 0 37076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_404
timestamp 1667941163
transform 1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_9
timestamp 1667941163
transform 1 0 1932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1667941163
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1667941163
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1667941163
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1667941163
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_62
timestamp 1667941163
transform 1 0 6808 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_77
timestamp 1667941163
transform 1 0 8188 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_89
timestamp 1667941163
transform 1 0 9292 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_101
timestamp 1667941163
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1667941163
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_180
timestamp 1667941163
transform 1 0 17664 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_186
timestamp 1667941163
transform 1 0 18216 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_196
timestamp 1667941163
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_208
timestamp 1667941163
transform 1 0 20240 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1667941163
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 1667941163
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1667941163
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1667941163
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1667941163
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1667941163
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_297
timestamp 1667941163
transform 1 0 28428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_305
timestamp 1667941163
transform 1 0 29164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_319
timestamp 1667941163
transform 1 0 30452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_326
timestamp 1667941163
transform 1 0 31096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1667941163
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1667941163
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1667941163
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_359
timestamp 1667941163
transform 1 0 34132 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_369
timestamp 1667941163
transform 1 0 35052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_376
timestamp 1667941163
transform 1 0 35696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_383
timestamp 1667941163
transform 1 0 36340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1667941163
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1667941163
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1667941163
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_214
timestamp 1667941163
transform 1 0 20792 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1667941163
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_233
timestamp 1667941163
transform 1 0 22540 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_239
timestamp 1667941163
transform 1 0 23092 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1667941163
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_261
timestamp 1667941163
transform 1 0 25116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_266
timestamp 1667941163
transform 1 0 25576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_291
timestamp 1667941163
transform 1 0 27876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_298
timestamp 1667941163
transform 1 0 28520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1667941163
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_324
timestamp 1667941163
transform 1 0 30912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_345
timestamp 1667941163
transform 1 0 32844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_369
timestamp 1667941163
transform 1 0 35052 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_373
timestamp 1667941163
transform 1 0 35420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_380
timestamp 1667941163
transform 1 0 36064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_387
timestamp 1667941163
transform 1 0 36708 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_394
timestamp 1667941163
transform 1 0 37352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1667941163
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_8
timestamp 1667941163
transform 1 0 1840 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_20
timestamp 1667941163
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_32
timestamp 1667941163
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1667941163
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_91
timestamp 1667941163
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1667941163
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_177
timestamp 1667941163
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_183
timestamp 1667941163
transform 1 0 17940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1667941163
transform 1 0 19044 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1667941163
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1667941163
transform 1 0 20700 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1667941163
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_230
timestamp 1667941163
transform 1 0 22264 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1667941163
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1667941163
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1667941163
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1667941163
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_286
timestamp 1667941163
transform 1 0 27416 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_298
timestamp 1667941163
transform 1 0 28520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_307
timestamp 1667941163
transform 1 0 29348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_311
timestamp 1667941163
transform 1 0 29716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1667941163
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1667941163
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_342
timestamp 1667941163
transform 1 0 32568 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_359
timestamp 1667941163
transform 1 0 34132 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_367
timestamp 1667941163
transform 1 0 34868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_383
timestamp 1667941163
transform 1 0 36340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_390
timestamp 1667941163
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1667941163
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1667941163
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_96
timestamp 1667941163
transform 1 0 9936 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_104
timestamp 1667941163
transform 1 0 10672 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_120
timestamp 1667941163
transform 1 0 12144 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_128
timestamp 1667941163
transform 1 0 12880 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1667941163
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_146
timestamp 1667941163
transform 1 0 14536 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_158
timestamp 1667941163
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_170
timestamp 1667941163
transform 1 0 16744 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp 1667941163
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_190
timestamp 1667941163
transform 1 0 18584 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1667941163
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_202
timestamp 1667941163
transform 1 0 19688 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_214
timestamp 1667941163
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_226
timestamp 1667941163
transform 1 0 21896 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_241
timestamp 1667941163
transform 1 0 23276 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1667941163
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_265
timestamp 1667941163
transform 1 0 25484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_270
timestamp 1667941163
transform 1 0 25944 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_287
timestamp 1667941163
transform 1 0 27508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1667941163
transform 1 0 28152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1667941163
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1667941163
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1667941163
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_331
timestamp 1667941163
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_343
timestamp 1667941163
transform 1 0 32660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_348
timestamp 1667941163
transform 1 0 33120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_355
timestamp 1667941163
transform 1 0 33764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_362
timestamp 1667941163
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_388
timestamp 1667941163
transform 1 0 36800 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1667941163
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_402
timestamp 1667941163
transform 1 0 38088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1667941163
transform 1 0 38456 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_73
timestamp 1667941163
transform 1 0 7820 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1667941163
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_89
timestamp 1667941163
transform 1 0 9292 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_97
timestamp 1667941163
transform 1 0 10028 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_101
timestamp 1667941163
transform 1 0 10396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1667941163
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1667941163
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_133
timestamp 1667941163
transform 1 0 13340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_142
timestamp 1667941163
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_200
timestamp 1667941163
transform 1 0 19504 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_212
timestamp 1667941163
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_234
timestamp 1667941163
transform 1 0 22632 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_241
timestamp 1667941163
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_248
timestamp 1667941163
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_255
timestamp 1667941163
transform 1 0 24564 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_264
timestamp 1667941163
transform 1 0 25392 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1667941163
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1667941163
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_288
timestamp 1667941163
transform 1 0 27600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_295
timestamp 1667941163
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_302
timestamp 1667941163
transform 1 0 28888 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_309
timestamp 1667941163
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_321
timestamp 1667941163
transform 1 0 30636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1667941163
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1667941163
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_355
timestamp 1667941163
transform 1 0 33764 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_359
timestamp 1667941163
transform 1 0 34132 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_364
timestamp 1667941163
transform 1 0 34592 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_371
timestamp 1667941163
transform 1 0 35236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_378
timestamp 1667941163
transform 1 0 35880 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_386
timestamp 1667941163
transform 1 0 36616 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1667941163
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_402
timestamp 1667941163
transform 1 0 38088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1667941163
transform 1 0 38456 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1667941163
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1667941163
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_95
timestamp 1667941163
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_99
timestamp 1667941163
transform 1 0 10212 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1667941163
transform 1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1667941163
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_150
timestamp 1667941163
transform 1 0 14904 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1667941163
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_166
timestamp 1667941163
transform 1 0 16376 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_178
timestamp 1667941163
transform 1 0 17480 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_220
timestamp 1667941163
transform 1 0 21344 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_237
timestamp 1667941163
transform 1 0 22908 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_243
timestamp 1667941163
transform 1 0 23460 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1667941163
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1667941163
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1667941163
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1667941163
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1667941163
transform 1 0 26496 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_293
timestamp 1667941163
transform 1 0 28060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1667941163
transform 1 0 28980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1667941163
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_314
timestamp 1667941163
transform 1 0 29992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_329
timestamp 1667941163
transform 1 0 31372 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1667941163
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_345
timestamp 1667941163
transform 1 0 32844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_351
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_357
timestamp 1667941163
transform 1 0 33948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1667941163
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_371
timestamp 1667941163
transform 1 0 35236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_378
timestamp 1667941163
transform 1 0 35880 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_385
timestamp 1667941163
transform 1 0 36524 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_391
timestamp 1667941163
transform 1 0 37076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_405
timestamp 1667941163
transform 1 0 38364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_8
timestamp 1667941163
transform 1 0 1840 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_20
timestamp 1667941163
transform 1 0 2944 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_32
timestamp 1667941163
transform 1 0 4048 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_44
timestamp 1667941163
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_72
timestamp 1667941163
transform 1 0 7728 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1667941163
transform 1 0 8464 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_90
timestamp 1667941163
transform 1 0 9384 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_96
timestamp 1667941163
transform 1 0 9936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1667941163
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1667941163
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_135
timestamp 1667941163
transform 1 0 13524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_144
timestamp 1667941163
transform 1 0 14352 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_152
timestamp 1667941163
transform 1 0 15088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1667941163
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1667941163
transform 1 0 17112 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1667941163
transform 1 0 17480 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_182
timestamp 1667941163
transform 1 0 17848 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_190
timestamp 1667941163
transform 1 0 18584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_196
timestamp 1667941163
transform 1 0 19136 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_204
timestamp 1667941163
transform 1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1667941163
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1667941163
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_230
timestamp 1667941163
transform 1 0 22264 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_242
timestamp 1667941163
transform 1 0 23368 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_250
timestamp 1667941163
transform 1 0 24104 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_257
timestamp 1667941163
transform 1 0 24748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_263
timestamp 1667941163
transform 1 0 25300 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1667941163
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1667941163
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1667941163
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_297
timestamp 1667941163
transform 1 0 28428 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_319
timestamp 1667941163
transform 1 0 30452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1667941163
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1667941163
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_342
timestamp 1667941163
transform 1 0 32568 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_351
timestamp 1667941163
transform 1 0 33396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_358
timestamp 1667941163
transform 1 0 34040 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_367
timestamp 1667941163
transform 1 0 34868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_374
timestamp 1667941163
transform 1 0 35512 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_383
timestamp 1667941163
transform 1 0 36340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1667941163
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1667941163
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_59
timestamp 1667941163
transform 1 0 6532 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_63
timestamp 1667941163
transform 1 0 6900 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_70
timestamp 1667941163
transform 1 0 7544 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_78
timestamp 1667941163
transform 1 0 8280 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1667941163
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1667941163
transform 1 0 9476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_100
timestamp 1667941163
transform 1 0 10304 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_108
timestamp 1667941163
transform 1 0 11040 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_112
timestamp 1667941163
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_120
timestamp 1667941163
transform 1 0 12144 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1667941163
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1667941163
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1667941163
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_156
timestamp 1667941163
transform 1 0 15456 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1667941163
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_179
timestamp 1667941163
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1667941163
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1667941163
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_222
timestamp 1667941163
transform 1 0 21528 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_237
timestamp 1667941163
transform 1 0 22908 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1667941163
transform 1 0 25668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_275
timestamp 1667941163
transform 1 0 26404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_283
timestamp 1667941163
transform 1 0 27140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_290
timestamp 1667941163
transform 1 0 27784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_297
timestamp 1667941163
transform 1 0 28428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1667941163
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_324
timestamp 1667941163
transform 1 0 30912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1667941163
transform 1 0 31556 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1667941163
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_345
timestamp 1667941163
transform 1 0 32844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_353
timestamp 1667941163
transform 1 0 33580 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1667941163
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_383
timestamp 1667941163
transform 1 0 36340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_390
timestamp 1667941163
transform 1 0 36984 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_397
timestamp 1667941163
transform 1 0 37628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_404
timestamp 1667941163
transform 1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_10
timestamp 1667941163
transform 1 0 2024 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_22
timestamp 1667941163
transform 1 0 3128 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_34
timestamp 1667941163
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1667941163
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1667941163
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_68
timestamp 1667941163
transform 1 0 7360 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_74
timestamp 1667941163
transform 1 0 7912 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_78
timestamp 1667941163
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp 1667941163
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_95
timestamp 1667941163
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1667941163
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_124
timestamp 1667941163
transform 1 0 12512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_145
timestamp 1667941163
transform 1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1667941163
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1667941163
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_184
timestamp 1667941163
transform 1 0 18032 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_188
timestamp 1667941163
transform 1 0 18400 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_195
timestamp 1667941163
transform 1 0 19044 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_207
timestamp 1667941163
transform 1 0 20148 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1667941163
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1667941163
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_233
timestamp 1667941163
transform 1 0 22540 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_263
timestamp 1667941163
transform 1 0 25300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_270
timestamp 1667941163
transform 1 0 25944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1667941163
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_289
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1667941163
transform 1 0 28704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_307
timestamp 1667941163
transform 1 0 29348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_314
timestamp 1667941163
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_321
timestamp 1667941163
transform 1 0 30636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1667941163
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_342
timestamp 1667941163
transform 1 0 32568 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_349
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_356
timestamp 1667941163
transform 1 0 33856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_371
timestamp 1667941163
transform 1 0 35236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_378
timestamp 1667941163
transform 1 0 35880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1667941163
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1667941163
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_398
timestamp 1667941163
transform 1 0 37720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_9
timestamp 1667941163
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1667941163
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1667941163
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1667941163
transform 1 0 10856 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_113
timestamp 1667941163
transform 1 0 11500 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_119
timestamp 1667941163
transform 1 0 12052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_123
timestamp 1667941163
transform 1 0 12420 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1667941163
transform 1 0 12788 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_131
timestamp 1667941163
transform 1 0 13156 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1667941163
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1667941163
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1667941163
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_174
timestamp 1667941163
transform 1 0 17112 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_182
timestamp 1667941163
transform 1 0 17848 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_187
timestamp 1667941163
transform 1 0 18308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1667941163
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_202
timestamp 1667941163
transform 1 0 19688 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1667941163
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_231
timestamp 1667941163
transform 1 0 22356 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_239
timestamp 1667941163
transform 1 0 23092 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1667941163
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_268
timestamp 1667941163
transform 1 0 25760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_272
timestamp 1667941163
transform 1 0 26128 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_279
timestamp 1667941163
transform 1 0 26772 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_286
timestamp 1667941163
transform 1 0 27416 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_298
timestamp 1667941163
transform 1 0 28520 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1667941163
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_314
timestamp 1667941163
transform 1 0 29992 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_320
timestamp 1667941163
transform 1 0 30544 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_324
timestamp 1667941163
transform 1 0 30912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_331
timestamp 1667941163
transform 1 0 31556 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_338
timestamp 1667941163
transform 1 0 32200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_351
timestamp 1667941163
transform 1 0 33396 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1667941163
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_380
timestamp 1667941163
transform 1 0 36064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_387
timestamp 1667941163
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_394
timestamp 1667941163
transform 1 0 37352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1667941163
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_9
timestamp 1667941163
transform 1 0 1932 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_16
timestamp 1667941163
transform 1 0 2576 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_28
timestamp 1667941163
transform 1 0 3680 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_43
timestamp 1667941163
transform 1 0 5060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1667941163
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_74
timestamp 1667941163
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_78
timestamp 1667941163
transform 1 0 8280 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1667941163
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1667941163
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_106
timestamp 1667941163
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 1667941163
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_129
timestamp 1667941163
transform 1 0 12972 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_133
timestamp 1667941163
transform 1 0 13340 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_145
timestamp 1667941163
transform 1 0 14444 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_157
timestamp 1667941163
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1667941163
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_174
timestamp 1667941163
transform 1 0 17112 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_183
timestamp 1667941163
transform 1 0 17940 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_195
timestamp 1667941163
transform 1 0 19044 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_207
timestamp 1667941163
transform 1 0 20148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1667941163
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1667941163
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_238
timestamp 1667941163
transform 1 0 23000 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_250
timestamp 1667941163
transform 1 0 24104 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_258
timestamp 1667941163
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1667941163
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1667941163
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1667941163
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1667941163
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1667941163
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_317
timestamp 1667941163
transform 1 0 30268 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_321
timestamp 1667941163
transform 1 0 30636 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_329
timestamp 1667941163
transform 1 0 31372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1667941163
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_345
timestamp 1667941163
transform 1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_369
timestamp 1667941163
transform 1 0 35052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_378
timestamp 1667941163
transform 1 0 35880 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_384
timestamp 1667941163
transform 1 0 36432 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1667941163
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_398
timestamp 1667941163
transform 1 0 37720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_35
timestamp 1667941163
transform 1 0 4324 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_44
timestamp 1667941163
transform 1 0 5152 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_56
timestamp 1667941163
transform 1 0 6256 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_68
timestamp 1667941163
transform 1 0 7360 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_76
timestamp 1667941163
transform 1 0 8096 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1667941163
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_96
timestamp 1667941163
transform 1 0 9936 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_108
timestamp 1667941163
transform 1 0 11040 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1667941163
transform 1 0 12144 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_130
timestamp 1667941163
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1667941163
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1667941163
transform 1 0 14444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1667941163
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_166
timestamp 1667941163
transform 1 0 16376 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_178
timestamp 1667941163
transform 1 0 17480 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_209
timestamp 1667941163
transform 1 0 20332 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1667941163
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_219
timestamp 1667941163
transform 1 0 21252 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_231
timestamp 1667941163
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_241
timestamp 1667941163
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1667941163
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_285
timestamp 1667941163
transform 1 0 27324 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_297
timestamp 1667941163
transform 1 0 28428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1667941163
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_321
timestamp 1667941163
transform 1 0 30636 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1667941163
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1667941163
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_380
timestamp 1667941163
transform 1 0 36064 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_386
timestamp 1667941163
transform 1 0 36616 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_390
timestamp 1667941163
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_8
timestamp 1667941163
transform 1 0 1840 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_20
timestamp 1667941163
transform 1 0 2944 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1667941163
transform 1 0 4048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_36
timestamp 1667941163
transform 1 0 4416 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_40
timestamp 1667941163
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1667941163
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_87
timestamp 1667941163
transform 1 0 9108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_101
timestamp 1667941163
transform 1 0 10396 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1667941163
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1667941163
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_131
timestamp 1667941163
transform 1 0 13156 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_143
timestamp 1667941163
transform 1 0 14260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_155
timestamp 1667941163
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_177
timestamp 1667941163
transform 1 0 17388 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_203
timestamp 1667941163
transform 1 0 19780 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1667941163
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1667941163
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_257
timestamp 1667941163
transform 1 0 24748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1667941163
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1667941163
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_303
timestamp 1667941163
transform 1 0 28980 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_315
timestamp 1667941163
transform 1 0 30084 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_327
timestamp 1667941163
transform 1 0 31188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_343
timestamp 1667941163
transform 1 0 32660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_364
timestamp 1667941163
transform 1 0 34592 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1667941163
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1667941163
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1667941163
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1667941163
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_105
timestamp 1667941163
transform 1 0 10764 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_114
timestamp 1667941163
transform 1 0 11592 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_122
timestamp 1667941163
transform 1 0 12328 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_126
timestamp 1667941163
transform 1 0 12696 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1667941163
transform 1 0 14812 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_171
timestamp 1667941163
transform 1 0 16836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_183
timestamp 1667941163
transform 1 0 17940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1667941163
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1667941163
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_265
timestamp 1667941163
transform 1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_291
timestamp 1667941163
transform 1 0 27876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1667941163
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1667941163
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_331
timestamp 1667941163
transform 1 0 31556 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_355
timestamp 1667941163
transform 1 0 33764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1667941163
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_390
timestamp 1667941163
transform 1 0 36984 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_398
timestamp 1667941163
transform 1 0 37720 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_402
timestamp 1667941163
transform 1 0 38088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1667941163
transform 1 0 38456 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_47
timestamp 1667941163
transform 1 0 5428 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_62
timestamp 1667941163
transform 1 0 6808 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_74
timestamp 1667941163
transform 1 0 7912 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1667941163
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_104
timestamp 1667941163
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_130
timestamp 1667941163
transform 1 0 13064 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1667941163
transform 1 0 14168 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1667941163
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_192
timestamp 1667941163
transform 1 0 18768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_198
timestamp 1667941163
transform 1 0 19320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_237
timestamp 1667941163
transform 1 0 22908 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_268
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_320
timestamp 1667941163
transform 1 0 30544 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1667941163
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_359
timestamp 1667941163
transform 1 0 34132 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_383
timestamp 1667941163
transform 1 0 36340 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1667941163
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1667941163
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_63
timestamp 1667941163
transform 1 0 6900 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_70
timestamp 1667941163
transform 1 0 7544 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1667941163
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_93
timestamp 1667941163
transform 1 0 9660 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_117
timestamp 1667941163
transform 1 0 11868 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_128
timestamp 1667941163
transform 1 0 12880 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1667941163
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_182
timestamp 1667941163
transform 1 0 17848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_219
timestamp 1667941163
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_231
timestamp 1667941163
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_243
timestamp 1667941163
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1667941163
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1667941163
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1667941163
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_289
timestamp 1667941163
transform 1 0 27692 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1667941163
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_331
timestamp 1667941163
transform 1 0 31556 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_343
timestamp 1667941163
transform 1 0 32660 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1667941163
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_387
timestamp 1667941163
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_399
timestamp 1667941163
transform 1 0 37812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1667941163
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_21
timestamp 1667941163
transform 1 0 3036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_29
timestamp 1667941163
transform 1 0 3772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_33
timestamp 1667941163
transform 1 0 4140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_40
timestamp 1667941163
transform 1 0 4784 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_47
timestamp 1667941163
transform 1 0 5428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1667941163
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_61
timestamp 1667941163
transform 1 0 6716 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_70
timestamp 1667941163
transform 1 0 7544 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_77
timestamp 1667941163
transform 1 0 8188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1667941163
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1667941163
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_117
timestamp 1667941163
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_127
timestamp 1667941163
transform 1 0 12788 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_134
timestamp 1667941163
transform 1 0 13432 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_146
timestamp 1667941163
transform 1 0 14536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1667941163
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1667941163
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1667941163
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1667941163
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_238
timestamp 1667941163
transform 1 0 23000 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_250
timestamp 1667941163
transform 1 0 24104 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_262
timestamp 1667941163
transform 1 0 25208 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1667941163
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_293
timestamp 1667941163
transform 1 0 28060 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_316
timestamp 1667941163
transform 1 0 30176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1667941163
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_349
timestamp 1667941163
transform 1 0 33212 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1667941163
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1667941163
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1667941163
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1667941163
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_49
timestamp 1667941163
transform 1 0 5612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_61
timestamp 1667941163
transform 1 0 6716 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1667941163
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_96
timestamp 1667941163
transform 1 0 9936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_100
timestamp 1667941163
transform 1 0 10304 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_104
timestamp 1667941163
transform 1 0 10672 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_116
timestamp 1667941163
transform 1 0 11776 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_128
timestamp 1667941163
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_150
timestamp 1667941163
transform 1 0 14904 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_179
timestamp 1667941163
transform 1 0 17572 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1667941163
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1667941163
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1667941163
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_221
timestamp 1667941163
transform 1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_227
timestamp 1667941163
transform 1 0 21988 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1667941163
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_282
timestamp 1667941163
transform 1 0 27048 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_294
timestamp 1667941163
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_317
timestamp 1667941163
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_341
timestamp 1667941163
transform 1 0 32476 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_353
timestamp 1667941163
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1667941163
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_387
timestamp 1667941163
transform 1 0 36708 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_394
timestamp 1667941163
transform 1 0 37352 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_400
timestamp 1667941163
transform 1 0 37904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_45
timestamp 1667941163
transform 1 0 5244 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 1667941163
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_72
timestamp 1667941163
transform 1 0 7728 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_80
timestamp 1667941163
transform 1 0 8464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_86
timestamp 1667941163
transform 1 0 9016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1667941163
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_118
timestamp 1667941163
transform 1 0 11960 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_130
timestamp 1667941163
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_136
timestamp 1667941163
transform 1 0 13616 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_140
timestamp 1667941163
transform 1 0 13984 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_152
timestamp 1667941163
transform 1 0 15088 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1667941163
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1667941163
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_193
timestamp 1667941163
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1667941163
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_257
timestamp 1667941163
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1667941163
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1667941163
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_303
timestamp 1667941163
transform 1 0 28980 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1667941163
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1667941163
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_349
timestamp 1667941163
transform 1 0 33212 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_353
timestamp 1667941163
transform 1 0 33580 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_377
timestamp 1667941163
transform 1 0 35788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_389
timestamp 1667941163
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_397
timestamp 1667941163
transform 1 0 37628 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_401
timestamp 1667941163
transform 1 0 37996 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_8
timestamp 1667941163
transform 1 0 1840 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1667941163
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_50
timestamp 1667941163
transform 1 0 5704 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_62
timestamp 1667941163
transform 1 0 6808 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_70
timestamp 1667941163
transform 1 0 7544 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1667941163
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_90
timestamp 1667941163
transform 1 0 9384 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_102
timestamp 1667941163
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1667941163
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1667941163
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_179
timestamp 1667941163
transform 1 0 17572 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1667941163
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1667941163
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_236
timestamp 1667941163
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1667941163
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_265
timestamp 1667941163
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_291
timestamp 1667941163
transform 1 0 27876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_303
timestamp 1667941163
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1667941163
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_321
timestamp 1667941163
transform 1 0 30636 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_329
timestamp 1667941163
transform 1 0 31372 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_350
timestamp 1667941163
transform 1 0 33304 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1667941163
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_378
timestamp 1667941163
transform 1 0 35880 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_390
timestamp 1667941163
transform 1 0 36984 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp 1667941163
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_70
timestamp 1667941163
transform 1 0 7544 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_78
timestamp 1667941163
transform 1 0 8280 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_92
timestamp 1667941163
transform 1 0 9568 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1667941163
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_117
timestamp 1667941163
transform 1 0 11868 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_121
timestamp 1667941163
transform 1 0 12236 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_133
timestamp 1667941163
transform 1 0 13340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_145
timestamp 1667941163
transform 1 0 14444 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1667941163
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_174
timestamp 1667941163
transform 1 0 17112 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_182
timestamp 1667941163
transform 1 0 17848 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_206
timestamp 1667941163
transform 1 0 20056 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_218
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1667941163
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1667941163
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1667941163
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1667941163
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1667941163
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1667941163
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_287
timestamp 1667941163
transform 1 0 27508 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_299
timestamp 1667941163
transform 1 0 28612 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_307
timestamp 1667941163
transform 1 0 29348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_330
timestamp 1667941163
transform 1 0 31464 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_349
timestamp 1667941163
transform 1 0 33212 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_375
timestamp 1667941163
transform 1 0 35604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1667941163
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1667941163
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1667941163
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_9
timestamp 1667941163
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1667941163
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_59
timestamp 1667941163
transform 1 0 6532 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_63
timestamp 1667941163
transform 1 0 6900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_70
timestamp 1667941163
transform 1 0 7544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1667941163
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_120
timestamp 1667941163
transform 1 0 12144 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1667941163
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_146
timestamp 1667941163
transform 1 0 14536 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_179
timestamp 1667941163
transform 1 0 17572 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1667941163
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_219
timestamp 1667941163
transform 1 0 21252 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_223
timestamp 1667941163
transform 1 0 21620 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_235
timestamp 1667941163
transform 1 0 22724 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1667941163
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1667941163
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_277
timestamp 1667941163
transform 1 0 26588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1667941163
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1667941163
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_338
timestamp 1667941163
transform 1 0 32200 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_387
timestamp 1667941163
transform 1 0 36708 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_399
timestamp 1667941163
transform 1 0 37812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_405
timestamp 1667941163
transform 1 0 38364 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_75
timestamp 1667941163
transform 1 0 8004 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_95
timestamp 1667941163
transform 1 0 9844 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_102
timestamp 1667941163
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1667941163
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_118
timestamp 1667941163
transform 1 0 11960 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_126
timestamp 1667941163
transform 1 0 12696 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_140
timestamp 1667941163
transform 1 0 13984 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1667941163
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_204
timestamp 1667941163
transform 1 0 19872 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_216
timestamp 1667941163
transform 1 0 20976 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_250
timestamp 1667941163
transform 1 0 24104 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_262
timestamp 1667941163
transform 1 0 25208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1667941163
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_306
timestamp 1667941163
transform 1 0 29256 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_318
timestamp 1667941163
transform 1 0 30360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1667941163
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_345
timestamp 1667941163
transform 1 0 32844 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_369
timestamp 1667941163
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_381
timestamp 1667941163
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1667941163
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1667941163
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_38
timestamp 1667941163
transform 1 0 4600 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_45
timestamp 1667941163
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_57
timestamp 1667941163
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_61
timestamp 1667941163
transform 1 0 6716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_69
timestamp 1667941163
transform 1 0 7452 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_73
timestamp 1667941163
transform 1 0 7820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1667941163
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_93
timestamp 1667941163
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_105
timestamp 1667941163
transform 1 0 10764 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_112
timestamp 1667941163
transform 1 0 11408 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_131
timestamp 1667941163
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1667941163
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_161
timestamp 1667941163
transform 1 0 15916 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_184
timestamp 1667941163
transform 1 0 18032 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_229
timestamp 1667941163
transform 1 0 22172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_241
timestamp 1667941163
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1667941163
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1667941163
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1667941163
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1667941163
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1667941163
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1667941163
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1667941163
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_333
timestamp 1667941163
transform 1 0 31740 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1667941163
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1667941163
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1667941163
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1667941163
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_42
timestamp 1667941163
transform 1 0 4968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1667941163
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_89
timestamp 1667941163
transform 1 0 9292 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_118
timestamp 1667941163
transform 1 0 11960 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_126
timestamp 1667941163
transform 1 0 12696 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1667941163
transform 1 0 14168 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_182
timestamp 1667941163
transform 1 0 17848 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_186
timestamp 1667941163
transform 1 0 18216 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_207
timestamp 1667941163
transform 1 0 20148 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1667941163
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_230
timestamp 1667941163
transform 1 0 22264 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_242
timestamp 1667941163
transform 1 0 23368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_254
timestamp 1667941163
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_266
timestamp 1667941163
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1667941163
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_304
timestamp 1667941163
transform 1 0 29072 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_316
timestamp 1667941163
transform 1 0 30176 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_328
timestamp 1667941163
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_343
timestamp 1667941163
transform 1 0 32660 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_364
timestamp 1667941163
transform 1 0 34592 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_376
timestamp 1667941163
transform 1 0 35696 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1667941163
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1667941163
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1667941163
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_9
timestamp 1667941163
transform 1 0 1932 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1667941163
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_35
timestamp 1667941163
transform 1 0 4324 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_47
timestamp 1667941163
transform 1 0 5428 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_59
timestamp 1667941163
transform 1 0 6532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_71
timestamp 1667941163
transform 1 0 7636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_108
timestamp 1667941163
transform 1 0 11040 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_115
timestamp 1667941163
transform 1 0 11684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_119
timestamp 1667941163
transform 1 0 12052 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1667941163
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_151
timestamp 1667941163
transform 1 0 14996 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_178
timestamp 1667941163
transform 1 0 17480 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1667941163
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_209
timestamp 1667941163
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_235
timestamp 1667941163
transform 1 0 22724 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1667941163
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1667941163
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_287
timestamp 1667941163
transform 1 0 27508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_299
timestamp 1667941163
transform 1 0 28612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1667941163
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_334
timestamp 1667941163
transform 1 0 31832 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_358
timestamp 1667941163
transform 1 0 34040 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_390
timestamp 1667941163
transform 1 0 36984 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_398
timestamp 1667941163
transform 1 0 37720 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_90
timestamp 1667941163
transform 1 0 9384 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_97
timestamp 1667941163
transform 1 0 10028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1667941163
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_124
timestamp 1667941163
transform 1 0 12512 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_132
timestamp 1667941163
transform 1 0 13248 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_136
timestamp 1667941163
transform 1 0 13616 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_144
timestamp 1667941163
transform 1 0 14352 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1667941163
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1667941163
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_189
timestamp 1667941163
transform 1 0 18492 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_211
timestamp 1667941163
transform 1 0 20516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1667941163
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1667941163
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1667941163
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1667941163
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_293
timestamp 1667941163
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_301
timestamp 1667941163
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_315
timestamp 1667941163
transform 1 0 30084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1667941163
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_361
timestamp 1667941163
transform 1 0 34316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_367
timestamp 1667941163
transform 1 0 34868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1667941163
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_401
timestamp 1667941163
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1667941163
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_89
timestamp 1667941163
transform 1 0 9292 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1667941163
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_116
timestamp 1667941163
transform 1 0 11776 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_123
timestamp 1667941163
transform 1 0 12420 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1667941163
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_146
timestamp 1667941163
transform 1 0 14536 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_152
timestamp 1667941163
transform 1 0 15088 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_176
timestamp 1667941163
transform 1 0 17296 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_182
timestamp 1667941163
transform 1 0 17848 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1667941163
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_221
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1667941163
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_278
timestamp 1667941163
transform 1 0 26680 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_290
timestamp 1667941163
transform 1 0 27784 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1667941163
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_321
timestamp 1667941163
transform 1 0 30636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_345
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1667941163
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 1667941163
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_381
timestamp 1667941163
transform 1 0 36156 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1667941163
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_36
timestamp 1667941163
transform 1 0 4416 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_48
timestamp 1667941163
transform 1 0 5520 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_62
timestamp 1667941163
transform 1 0 6808 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_74
timestamp 1667941163
transform 1 0 7912 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_84
timestamp 1667941163
transform 1 0 8832 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_91
timestamp 1667941163
transform 1 0 9476 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_98
timestamp 1667941163
transform 1 0 10120 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_118
timestamp 1667941163
transform 1 0 11960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_130
timestamp 1667941163
transform 1 0 13064 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_144
timestamp 1667941163
transform 1 0 14352 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_150
timestamp 1667941163
transform 1 0 14904 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_154
timestamp 1667941163
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1667941163
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_189
timestamp 1667941163
transform 1 0 18492 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_211
timestamp 1667941163
transform 1 0 20516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1667941163
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1667941163
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1667941163
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1667941163
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1667941163
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1667941163
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1667941163
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1667941163
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1667941163
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1667941163
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1667941163
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_349
timestamp 1667941163
transform 1 0 33212 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_372
timestamp 1667941163
transform 1 0 35328 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_379
timestamp 1667941163
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1667941163
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1667941163
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_90
timestamp 1667941163
transform 1 0 9384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_105
timestamp 1667941163
transform 1 0 10764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1667941163
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_149
timestamp 1667941163
transform 1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_172
timestamp 1667941163
transform 1 0 16928 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_184
timestamp 1667941163
transform 1 0 18032 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_219
timestamp 1667941163
transform 1 0 21252 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_227
timestamp 1667941163
transform 1 0 21988 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1667941163
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_258
timestamp 1667941163
transform 1 0 24840 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_270
timestamp 1667941163
transform 1 0 25944 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_278
timestamp 1667941163
transform 1 0 26680 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_283
timestamp 1667941163
transform 1 0 27140 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_290
timestamp 1667941163
transform 1 0 27784 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_302
timestamp 1667941163
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_333
timestamp 1667941163
transform 1 0 31740 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1667941163
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_377
timestamp 1667941163
transform 1 0 35788 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_383
timestamp 1667941163
transform 1 0 36340 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_395
timestamp 1667941163
transform 1 0 37444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1667941163
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1667941163
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1667941163
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1667941163
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1667941163
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_74
timestamp 1667941163
transform 1 0 7912 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_86
timestamp 1667941163
transform 1 0 9016 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_98
timestamp 1667941163
transform 1 0 10120 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_102
timestamp 1667941163
transform 1 0 10488 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1667941163
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_118
timestamp 1667941163
transform 1 0 11960 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_133
timestamp 1667941163
transform 1 0 13340 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_139
timestamp 1667941163
transform 1 0 13892 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_151
timestamp 1667941163
transform 1 0 14996 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1667941163
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_191
timestamp 1667941163
transform 1 0 18676 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_199
timestamp 1667941163
transform 1 0 19412 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1667941163
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_250
timestamp 1667941163
transform 1 0 24104 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_256
timestamp 1667941163
transform 1 0 24656 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1667941163
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1667941163
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1667941163
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1667941163
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1667941163
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1667941163
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1667941163
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1667941163
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1667941163
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_401
timestamp 1667941163
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1667941163
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1667941163
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1667941163
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_71
timestamp 1667941163
transform 1 0 7636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_90
timestamp 1667941163
transform 1 0 9384 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_98
timestamp 1667941163
transform 1 0 10120 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_102
timestamp 1667941163
transform 1 0 10488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_116
timestamp 1667941163
transform 1 0 11776 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_124
timestamp 1667941163
transform 1 0 12512 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1667941163
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_152
timestamp 1667941163
transform 1 0 15088 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_164
timestamp 1667941163
transform 1 0 16192 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_176
timestamp 1667941163
transform 1 0 17296 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1667941163
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_213
timestamp 1667941163
transform 1 0 20700 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_234
timestamp 1667941163
transform 1 0 22632 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1667941163
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_262
timestamp 1667941163
transform 1 0 25208 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_273
timestamp 1667941163
transform 1 0 26220 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1667941163
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1667941163
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1667941163
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1667941163
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1667941163
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1667941163
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_389
timestamp 1667941163
transform 1 0 36892 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_48
timestamp 1667941163
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_73
timestamp 1667941163
transform 1 0 7820 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_83
timestamp 1667941163
transform 1 0 8740 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_90
timestamp 1667941163
transform 1 0 9384 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_98
timestamp 1667941163
transform 1 0 10120 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_108
timestamp 1667941163
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_118
timestamp 1667941163
transform 1 0 11960 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_131
timestamp 1667941163
transform 1 0 13156 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_135
timestamp 1667941163
transform 1 0 13524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_141
timestamp 1667941163
transform 1 0 14076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_145
timestamp 1667941163
transform 1 0 14444 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_157
timestamp 1667941163
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1667941163
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_192
timestamp 1667941163
transform 1 0 18768 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_196
timestamp 1667941163
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1667941163
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_293
timestamp 1667941163
transform 1 0 28060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_320
timestamp 1667941163
transform 1 0 30544 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_327
timestamp 1667941163
transform 1 0 31188 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1667941163
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_345
timestamp 1667941163
transform 1 0 32844 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_357
timestamp 1667941163
transform 1 0 33948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_369
timestamp 1667941163
transform 1 0 35052 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_373
timestamp 1667941163
transform 1 0 35420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1667941163
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_12
timestamp 1667941163
transform 1 0 2208 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1667941163
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1667941163
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_102
timestamp 1667941163
transform 1 0 10488 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_110
timestamp 1667941163
transform 1 0 11224 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_114
timestamp 1667941163
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_129
timestamp 1667941163
transform 1 0 12972 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_134
timestamp 1667941163
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_147
timestamp 1667941163
transform 1 0 14628 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_176
timestamp 1667941163
transform 1 0 17296 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_188
timestamp 1667941163
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1667941163
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_261
timestamp 1667941163
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_267
timestamp 1667941163
transform 1 0 25668 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_279
timestamp 1667941163
transform 1 0 26772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_298
timestamp 1667941163
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1667941163
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_316
timestamp 1667941163
transform 1 0 30176 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_328
timestamp 1667941163
transform 1 0 31280 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_349
timestamp 1667941163
transform 1 0 33212 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_357
timestamp 1667941163
transform 1 0 33948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_361
timestamp 1667941163
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_387
timestamp 1667941163
transform 1 0 36708 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_399
timestamp 1667941163
transform 1 0 37812 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1667941163
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_16
timestamp 1667941163
transform 1 0 2576 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_28
timestamp 1667941163
transform 1 0 3680 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_33
timestamp 1667941163
transform 1 0 4140 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_43
timestamp 1667941163
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_80
timestamp 1667941163
transform 1 0 8464 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_88
timestamp 1667941163
transform 1 0 9200 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_102
timestamp 1667941163
transform 1 0 10488 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1667941163
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_118
timestamp 1667941163
transform 1 0 11960 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_126
timestamp 1667941163
transform 1 0 12696 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_138
timestamp 1667941163
transform 1 0 13800 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1667941163
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1667941163
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_213
timestamp 1667941163
transform 1 0 20700 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_253
timestamp 1667941163
transform 1 0 24380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_265
timestamp 1667941163
transform 1 0 25484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1667941163
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_306
timestamp 1667941163
transform 1 0 29256 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_325
timestamp 1667941163
transform 1 0 31004 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1667941163
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_359
timestamp 1667941163
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_371
timestamp 1667941163
transform 1 0 35236 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1667941163
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_8
timestamp 1667941163
transform 1 0 1840 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_38
timestamp 1667941163
transform 1 0 4600 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_50
timestamp 1667941163
transform 1 0 5704 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_61
timestamp 1667941163
transform 1 0 6716 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_73
timestamp 1667941163
transform 1 0 7820 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1667941163
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_122
timestamp 1667941163
transform 1 0 12328 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_128
timestamp 1667941163
transform 1 0 12880 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1667941163
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_146
timestamp 1667941163
transform 1 0 14536 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_154
timestamp 1667941163
transform 1 0 15272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_176
timestamp 1667941163
transform 1 0 17296 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_182
timestamp 1667941163
transform 1 0 17848 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1667941163
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_230
timestamp 1667941163
transform 1 0 22264 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_236
timestamp 1667941163
transform 1 0 22816 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_240
timestamp 1667941163
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_328
timestamp 1667941163
transform 1 0 31280 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_336
timestamp 1667941163
transform 1 0 32016 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1667941163
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_390
timestamp 1667941163
transform 1 0 36984 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_397
timestamp 1667941163
transform 1 0 37628 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_405
timestamp 1667941163
transform 1 0 38364 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1667941163
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_16
timestamp 1667941163
transform 1 0 2576 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_29
timestamp 1667941163
transform 1 0 3772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_41
timestamp 1667941163
transform 1 0 4876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1667941163
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_62
timestamp 1667941163
transform 1 0 6808 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_74
timestamp 1667941163
transform 1 0 7912 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_89
timestamp 1667941163
transform 1 0 9292 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_99
timestamp 1667941163
transform 1 0 10212 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_106
timestamp 1667941163
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_128
timestamp 1667941163
transform 1 0 12880 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1667941163
transform 1 0 13524 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_143
timestamp 1667941163
transform 1 0 14260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_148
timestamp 1667941163
transform 1 0 14720 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_152
timestamp 1667941163
transform 1 0 15088 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1667941163
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_191
timestamp 1667941163
transform 1 0 18676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_197
timestamp 1667941163
transform 1 0 19228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_218
timestamp 1667941163
transform 1 0 21160 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_229
timestamp 1667941163
transform 1 0 22172 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_250
timestamp 1667941163
transform 1 0 24104 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_262
timestamp 1667941163
transform 1 0 25208 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1667941163
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_304
timestamp 1667941163
transform 1 0 29072 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_319
timestamp 1667941163
transform 1 0 30452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_331
timestamp 1667941163
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_369
timestamp 1667941163
transform 1 0 35052 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_378
timestamp 1667941163
transform 1 0 35880 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1667941163
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_34
timestamp 1667941163
transform 1 0 4232 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_46
timestamp 1667941163
transform 1 0 5336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_58
timestamp 1667941163
transform 1 0 6440 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_64
timestamp 1667941163
transform 1 0 6992 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_75
timestamp 1667941163
transform 1 0 8004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1667941163
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 1667941163
transform 1 0 9476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_95
timestamp 1667941163
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_99
timestamp 1667941163
transform 1 0 10212 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_103
timestamp 1667941163
transform 1 0 10580 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_110
timestamp 1667941163
transform 1 0 11224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_117
timestamp 1667941163
transform 1 0 11868 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_125
timestamp 1667941163
transform 1 0 12604 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1667941163
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_157
timestamp 1667941163
transform 1 0 15548 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_184
timestamp 1667941163
transform 1 0 18032 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1667941163
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_257
timestamp 1667941163
transform 1 0 24748 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_278
timestamp 1667941163
transform 1 0 26680 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_285
timestamp 1667941163
transform 1 0 27324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_292
timestamp 1667941163
transform 1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_299
timestamp 1667941163
transform 1 0 28612 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1667941163
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_314
timestamp 1667941163
transform 1 0 29992 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_322
timestamp 1667941163
transform 1 0 30728 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_370
timestamp 1667941163
transform 1 0 35144 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_382
timestamp 1667941163
transform 1 0 36248 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_390
timestamp 1667941163
transform 1 0 36984 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_397
timestamp 1667941163
transform 1 0 37628 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_405
timestamp 1667941163
transform 1 0 38364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_18
timestamp 1667941163
transform 1 0 2760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_25
timestamp 1667941163
transform 1 0 3404 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_34
timestamp 1667941163
transform 1 0 4232 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_43
timestamp 1667941163
transform 1 0 5060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_65
timestamp 1667941163
transform 1 0 7084 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_71
timestamp 1667941163
transform 1 0 7636 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_78
timestamp 1667941163
transform 1 0 8280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_85
timestamp 1667941163
transform 1 0 8924 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_92
timestamp 1667941163
transform 1 0 9568 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1667941163
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_106
timestamp 1667941163
transform 1 0 10856 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_119
timestamp 1667941163
transform 1 0 12052 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_130
timestamp 1667941163
transform 1 0 13064 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_143
timestamp 1667941163
transform 1 0 14260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_150
timestamp 1667941163
transform 1 0 14904 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_158
timestamp 1667941163
transform 1 0 15640 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1667941163
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_177
timestamp 1667941163
transform 1 0 17388 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_200
timestamp 1667941163
transform 1 0 19504 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_212
timestamp 1667941163
transform 1 0 20608 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_253
timestamp 1667941163
transform 1 0 24380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1667941163
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_308
timestamp 1667941163
transform 1 0 29440 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1667941163
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_342
timestamp 1667941163
transform 1 0 32568 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_349
timestamp 1667941163
transform 1 0 33212 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_357
timestamp 1667941163
transform 1 0 33948 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_380
timestamp 1667941163
transform 1 0 36064 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_399
timestamp 1667941163
transform 1 0 37812 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_9
timestamp 1667941163
transform 1 0 1932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1667941163
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1667941163
transform 1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_48
timestamp 1667941163
transform 1 0 5520 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_62
timestamp 1667941163
transform 1 0 6808 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_77
timestamp 1667941163
transform 1 0 8188 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1667941163
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_105
timestamp 1667941163
transform 1 0 10764 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1667941163
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_126
timestamp 1667941163
transform 1 0 12696 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_134
timestamp 1667941163
transform 1 0 13432 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1667941163
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_147
timestamp 1667941163
transform 1 0 14628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_154
timestamp 1667941163
transform 1 0 15272 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_166
timestamp 1667941163
transform 1 0 16376 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1667941163
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_186
timestamp 1667941163
transform 1 0 18216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1667941163
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_210
timestamp 1667941163
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_222
timestamp 1667941163
transform 1 0 21528 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1667941163
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_239
timestamp 1667941163
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1667941163
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1667941163
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_258
timestamp 1667941163
transform 1 0 24840 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_266
timestamp 1667941163
transform 1 0 25576 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_278
timestamp 1667941163
transform 1 0 26680 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_287
timestamp 1667941163
transform 1 0 27508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_294
timestamp 1667941163
transform 1 0 28152 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1667941163
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1667941163
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_313
timestamp 1667941163
transform 1 0 29900 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_343
timestamp 1667941163
transform 1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_351
timestamp 1667941163
transform 1 0 33396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1667941163
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_371
timestamp 1667941163
transform 1 0 35236 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_379
timestamp 1667941163
transform 1 0 35972 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 1667941163
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 1667941163
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0384_
timestamp 1667941163
transform 1 0 28244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0385_
timestamp 1667941163
transform 1 0 22632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0386_
timestamp 1667941163
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0387_
timestamp 1667941163
transform 1 0 22632 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0388_
timestamp 1667941163
transform 1 0 22172 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0389_
timestamp 1667941163
transform 1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0390_
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0391_
timestamp 1667941163
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0392_
timestamp 1667941163
transform 1 0 9384 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0393_
timestamp 1667941163
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0394_
timestamp 1667941163
transform 1 0 13064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0395_
timestamp 1667941163
transform 1 0 35788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0396_
timestamp 1667941163
transform 1 0 13064 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0398_
timestamp 1667941163
transform 1 0 31464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0399_
timestamp 1667941163
transform 1 0 36708 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0400_
timestamp 1667941163
transform 1 0 37720 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0401_
timestamp 1667941163
transform 1 0 30084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1667941163
transform 1 0 20148 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0403_
timestamp 1667941163
transform 1 0 19228 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0404_
timestamp 1667941163
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0405_
timestamp 1667941163
transform 1 0 33856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0406_
timestamp 1667941163
transform 1 0 34868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0407_
timestamp 1667941163
transform 1 0 29532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0408_
timestamp 1667941163
transform 1 0 29716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0409_
timestamp 1667941163
transform 1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0410_
timestamp 1667941163
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0411_
timestamp 1667941163
transform 1 0 32936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0412_
timestamp 1667941163
transform 1 0 33212 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0413_
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0414_
timestamp 1667941163
transform 1 0 9108 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0415_
timestamp 1667941163
transform 1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0416_
timestamp 1667941163
transform 1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0417_
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0418_
timestamp 1667941163
transform 1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0419_
timestamp 1667941163
transform 1 0 5152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0420_
timestamp 1667941163
transform 1 0 5428 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0421_
timestamp 1667941163
transform 1 0 4784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0422_
timestamp 1667941163
transform 1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0423_
timestamp 1667941163
transform 1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0424_
timestamp 1667941163
transform 1 0 4324 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0425_
timestamp 1667941163
transform 1 0 4968 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0426_
timestamp 1667941163
transform 1 0 7268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0427_
timestamp 1667941163
transform 1 0 6624 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0428_
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0429_
timestamp 1667941163
transform 1 0 3864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0430_
timestamp 1667941163
transform 1 0 4508 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0431_
timestamp 1667941163
transform 1 0 27876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0432_
timestamp 1667941163
transform 1 0 32292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0433_
timestamp 1667941163
transform 1 0 32568 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0434_
timestamp 1667941163
transform 1 0 32384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0435_
timestamp 1667941163
transform 1 0 23276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0436_
timestamp 1667941163
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0437_
timestamp 1667941163
transform 1 0 21988 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0438_
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0439_
timestamp 1667941163
transform 1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0440_
timestamp 1667941163
transform 1 0 29440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0441_
timestamp 1667941163
transform 1 0 14536 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0442_
timestamp 1667941163
transform 1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0443_
timestamp 1667941163
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0444_
timestamp 1667941163
transform 1 0 35880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0445_
timestamp 1667941163
transform 1 0 35512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1667941163
transform 1 0 32292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0447_
timestamp 1667941163
transform 1 0 33764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0448_
timestamp 1667941163
transform 1 0 34500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1667941163
transform 1 0 21988 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1667941163
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0451_
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0452_
timestamp 1667941163
transform 1 0 14720 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0453_
timestamp 1667941163
transform 1 0 19688 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0454_
timestamp 1667941163
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1667941163
transform 1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0456_
timestamp 1667941163
transform 1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0457_
timestamp 1667941163
transform 1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1667941163
transform 1 0 22356 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0459_
timestamp 1667941163
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0460_
timestamp 1667941163
transform 1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0461_
timestamp 1667941163
transform 1 0 29256 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0462_
timestamp 1667941163
transform 1 0 12880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0463_
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0464_
timestamp 1667941163
transform 1 0 10580 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0465_
timestamp 1667941163
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0466_
timestamp 1667941163
transform 1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0467_
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0468_
timestamp 1667941163
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0469_
timestamp 1667941163
transform 1 0 23552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0470_
timestamp 1667941163
transform 1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0471_
timestamp 1667941163
transform 1 0 32108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0472_
timestamp 1667941163
transform 1 0 29900 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0473_
timestamp 1667941163
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0474_
timestamp 1667941163
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0475_
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0476_
timestamp 1667941163
transform 1 0 32936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0477_
timestamp 1667941163
transform 1 0 29716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0478_
timestamp 1667941163
transform 1 0 32936 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0479_
timestamp 1667941163
transform 1 0 31280 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0480_
timestamp 1667941163
transform 1 0 24932 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0481_
timestamp 1667941163
transform 1 0 6440 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0482_
timestamp 1667941163
transform 1 0 10212 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0483_
timestamp 1667941163
transform 1 0 11500 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0484_
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0485_
timestamp 1667941163
transform 1 0 25024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0486_
timestamp 1667941163
transform 1 0 23736 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0487_
timestamp 1667941163
transform 1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488_
timestamp 1667941163
transform 1 0 32292 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489_
timestamp 1667941163
transform 1 0 32936 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1667941163
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1667941163
transform 1 0 23184 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1667941163
transform 1 0 15732 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1667941163
transform 1 0 12788 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1667941163
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1667941163
transform 1 0 9752 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496_
timestamp 1667941163
transform 1 0 8372 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497_
timestamp 1667941163
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498_
timestamp 1667941163
transform 1 0 11592 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0499_
timestamp 1667941163
transform 1 0 11684 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0500_
timestamp 1667941163
transform 1 0 16100 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 1667941163
transform 1 0 12328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502_
timestamp 1667941163
transform 1 0 34040 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503_
timestamp 1667941163
transform 1 0 34868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504_
timestamp 1667941163
transform 1 0 13156 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505_
timestamp 1667941163
transform 1 0 3864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1667941163
transform 1 0 9108 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507_
timestamp 1667941163
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508_
timestamp 1667941163
transform 1 0 14720 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509_
timestamp 1667941163
transform 1 0 18676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510_
timestamp 1667941163
transform 1 0 11224 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0511_
timestamp 1667941163
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1667941163
transform 1 0 10212 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0513_
timestamp 1667941163
transform 1 0 9108 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0514_
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1667941163
transform 1 0 7360 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1667941163
transform 1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1667941163
transform 1 0 24104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1667941163
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1667941163
transform 1 0 27140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0520_
timestamp 1667941163
transform 1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1667941163
transform 1 0 26128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1667941163
transform 1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1667941163
transform 1 0 30360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0526_
timestamp 1667941163
transform 1 0 17664 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1667941163
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1667941163
transform 1 0 12144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1667941163
transform 1 0 11684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1667941163
transform 1 0 11684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1667941163
transform 1 0 20516 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1667941163
transform 1 0 13248 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1667941163
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1667941163
transform 1 0 11408 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1667941163
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0538_
timestamp 1667941163
transform 1 0 8280 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539_
timestamp 1667941163
transform 1 0 9844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540_
timestamp 1667941163
transform 1 0 31556 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541_
timestamp 1667941163
transform 1 0 33672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0542_
timestamp 1667941163
transform 1 0 27140 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0543_
timestamp 1667941163
transform 1 0 14628 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0544_
timestamp 1667941163
transform 1 0 23552 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0545_
timestamp 1667941163
transform 1 0 31648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1667941163
transform 1 0 31556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0547_
timestamp 1667941163
transform 1 0 34040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0548_
timestamp 1667941163
transform 1 0 31280 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0549_
timestamp 1667941163
transform 1 0 16652 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1667941163
transform 1 0 4140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0552_
timestamp 1667941163
transform 1 0 32844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1667941163
transform 1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0554_
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0555_
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1667941163
transform 1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0557_
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0558_
timestamp 1667941163
transform 1 0 34040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0559_
timestamp 1667941163
transform 1 0 33580 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0560_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1667941163
transform 1 0 10488 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0562_
timestamp 1667941163
transform 1 0 19228 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0563_
timestamp 1667941163
transform 1 0 11684 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1667941163
transform 1 0 13156 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0565_
timestamp 1667941163
transform 1 0 9384 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1667941163
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0567_
timestamp 1667941163
transform 1 0 14536 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0568_
timestamp 1667941163
transform 1 0 25208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1667941163
transform 1 0 10396 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0570_
timestamp 1667941163
transform 1 0 10396 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1667941163
transform 1 0 16836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0572_
timestamp 1667941163
transform 1 0 2300 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0573_
timestamp 1667941163
transform 1 0 8188 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0574_
timestamp 1667941163
transform 1 0 26864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0575_
timestamp 1667941163
transform 1 0 27324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0576_
timestamp 1667941163
transform 1 0 14260 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0577_
timestamp 1667941163
transform 1 0 34132 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1667941163
transform 1 0 2300 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0579_
timestamp 1667941163
transform 1 0 9752 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0580_
timestamp 1667941163
transform 1 0 8280 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0581_
timestamp 1667941163
transform 1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1667941163
transform 1 0 10212 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0583_
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0584_
timestamp 1667941163
transform 1 0 29256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0585_
timestamp 1667941163
transform 1 0 14628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1667941163
transform 1 0 7360 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1667941163
transform 1 0 25392 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1667941163
transform 1 0 14168 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0589_
timestamp 1667941163
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0590_
timestamp 1667941163
transform 1 0 23000 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0591_
timestamp 1667941163
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0593_
timestamp 1667941163
transform 1 0 7728 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1667941163
transform 1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0595_
timestamp 1667941163
transform 1 0 14996 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1667941163
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0597_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1667941163
transform 1 0 20516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0599_
timestamp 1667941163
transform 1 0 11316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1667941163
transform 1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0601_
timestamp 1667941163
transform 1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0602_
timestamp 1667941163
transform 1 0 23552 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1667941163
transform 1 0 33488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0604_
timestamp 1667941163
transform 1 0 36064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1667941163
transform 1 0 29900 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0606_
timestamp 1667941163
transform 1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1667941163
transform 1 0 35696 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0608_
timestamp 1667941163
transform 1 0 30912 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1667941163
transform 1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0610_
timestamp 1667941163
transform 1 0 33488 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1667941163
transform 1 0 37720 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0612_
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0613_
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1667941163
transform 1 0 8372 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0615_
timestamp 1667941163
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1667941163
transform 1 0 22172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0617_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1667941163
transform 1 0 4784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1667941163
transform 1 0 35144 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1667941163
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1667941163
transform 1 0 35144 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1667941163
transform 1 0 22632 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1667941163
transform 1 0 27048 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1667941163
transform 1 0 9016 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1667941163
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1667941163
transform 1 0 23000 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1667941163
transform 1 0 7728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1667941163
transform 1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0630_
timestamp 1667941163
transform 1 0 34224 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1667941163
transform 1 0 9108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1667941163
transform 1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1667941163
transform 1 0 9108 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1667941163
transform 1 0 36432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1667941163
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1667941163
transform 1 0 27508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1667941163
transform 1 0 29808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1667941163
transform 1 0 23092 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1667941163
transform 1 0 36432 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1667941163
transform 1 0 35880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1667941163
transform 1 0 7636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1667941163
transform 1 0 28336 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1667941163
transform 1 0 27232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1667941163
transform 1 0 36432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1667941163
transform 1 0 37720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1667941163
transform 1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1667941163
transform 1 0 12420 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1667941163
transform 1 0 31924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1667941163
transform 1 0 29348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1667941163
transform 1 0 24472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1667941163
transform 1 0 8004 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1667941163
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1667941163
transform 1 0 6532 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1667941163
transform 1 0 13616 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1667941163
transform 1 0 6716 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1667941163
transform 1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1667941163
transform 1 0 9752 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1667941163
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1667941163
transform 1 0 7268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0660_
timestamp 1667941163
transform 1 0 36708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0661_
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0662_
timestamp 1667941163
transform 1 0 22908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1667941163
transform 1 0 4324 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1667941163
transform 1 0 7544 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1667941163
transform 1 0 20792 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0666_
timestamp 1667941163
transform 1 0 36616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1667941163
transform 1 0 12144 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1667941163
transform 1 0 13524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1667941163
transform 1 0 36064 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1667941163
transform 1 0 22908 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0671_
timestamp 1667941163
transform 1 0 7544 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1667941163
transform 1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1667941163
transform 1 0 29716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1667941163
transform 1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1667941163
transform 1 0 22172 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0678_
timestamp 1667941163
transform 1 0 34684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1667941163
transform 1 0 12788 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 1667941163
transform 1 0 38088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1667941163
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1667941163
transform 1 0 22264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 1667941163
transform 1 0 14260 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1667941163
transform 1 0 30360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1667941163
transform 1 0 5520 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1667941163
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1667941163
transform 1 0 14904 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1667941163
transform 1 0 34132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1667941163
transform 1 0 37628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1667941163
transform 1 0 32292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1667941163
transform 1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1667941163
transform 1 0 6808 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1667941163
transform 1 0 6532 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1667941163
transform 1 0 9108 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1667941163
transform 1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1667941163
transform 1 0 2760 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1667941163
transform 1 0 34868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1667941163
transform 1 0 18676 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1667941163
transform 1 0 34040 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0701_
timestamp 1667941163
transform 1 0 20056 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1667941163
transform 1 0 36708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1667941163
transform 1 0 36708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1667941163
transform 1 0 36248 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1667941163
transform 1 0 9200 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1667941163
transform 1 0 9752 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1667941163
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1667941163
transform 1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0709_
timestamp 1667941163
transform 1 0 23644 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1667941163
transform 1 0 23828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1667941163
transform 1 0 9108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0712_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20516 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0713_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26220 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0714_
timestamp 1667941163
transform 1 0 28428 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1667941163
transform 1 0 37076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1667941163
transform 1 0 36524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1667941163
transform 1 0 37720 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1667941163
transform 1 0 38088 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1667941163
transform 1 0 36708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1667941163
transform 1 0 37076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1667941163
transform 1 0 34960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1667941163
transform 1 0 22632 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1667941163
transform 1 0 25944 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1667941163
transform 1 0 24472 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0725_
timestamp 1667941163
transform 1 0 25116 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1667941163
transform 1 0 13064 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1667941163
transform 1 0 20792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1667941163
transform 1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1667941163
transform 1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1667941163
transform 1 0 11960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1667941163
transform 1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1667941163
transform 1 0 14076 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1667941163
transform 1 0 12880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1667941163
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1667941163
transform 1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0736_
timestamp 1667941163
transform 1 0 22724 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1667941163
transform 1 0 10580 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1667941163
transform 1 0 10580 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1667941163
transform 1 0 29072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1667941163
transform 1 0 28428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1667941163
transform 1 0 10764 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1667941163
transform 1 0 12144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1667941163
transform 1 0 12328 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1667941163
transform 1 0 10948 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1667941163
transform 1 0 9292 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1667941163
transform 1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0747_
timestamp 1667941163
transform 1 0 23552 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1667941163
transform 1 0 24288 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1667941163
transform 1 0 23644 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1667941163
transform 1 0 35236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1667941163
transform 1 0 35604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1667941163
transform 1 0 36064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1667941163
transform 1 0 30360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1667941163
transform 1 0 25116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1667941163
transform 1 0 31280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1667941163
transform 1 0 28612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1667941163
transform 1 0 23644 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0758_
timestamp 1667941163
transform 1 0 24748 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1667941163
transform 1 0 37352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0760_
timestamp 1667941163
transform 1 0 37444 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1667941163
transform 1 0 36432 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1667941163
transform 1 0 31464 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1667941163
transform 1 0 25668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1667941163
transform 1 0 36708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0766_
timestamp 1667941163
transform 1 0 34592 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1667941163
transform 1 0 18032 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1667941163
transform 1 0 18124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0769_
timestamp 1667941163
transform 1 0 20976 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1667941163
transform 1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1667941163
transform 1 0 17296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1667941163
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1667941163
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1667941163
transform 1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1667941163
transform 1 0 32568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1667941163
transform 1 0 36248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1667941163
transform 1 0 30360 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1667941163
transform 1 0 24932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0780_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21344 0 1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1667941163
transform 1 0 25668 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1667941163
transform 1 0 23276 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1667941163
transform 1 0 11684 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1667941163
transform 1 0 11684 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0785_
timestamp 1667941163
transform 1 0 11960 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1667941163
transform 1 0 12328 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1667941163
transform 1 0 11316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1667941163
transform 1 0 32292 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1667941163
transform 1 0 35604 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1667941163
transform 1 0 32936 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0791_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1667941163
transform 1 0 26220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1667941163
transform 1 0 17572 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1667941163
transform 1 0 11684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1667941163
transform 1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1667941163
transform 1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1667941163
transform 1 0 9936 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1667941163
transform 1 0 8648 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1667941163
transform 1 0 10304 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1667941163
transform 1 0 27784 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0802_
timestamp 1667941163
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1667941163
transform 1 0 38088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1667941163
transform 1 0 37444 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1667941163
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1667941163
transform 1 0 25392 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1667941163
transform 1 0 27508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1667941163
transform 1 0 36708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1667941163
transform 1 0 29072 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1667941163
transform 1 0 37352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1667941163
transform 1 0 36248 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1667941163
transform 1 0 36064 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0813_
timestamp 1667941163
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1667941163
transform 1 0 33488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0815_
timestamp 1667941163
transform 1 0 37812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1667941163
transform 1 0 33764 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1667941163
transform 1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1667941163
transform 1 0 34960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1667941163
transform 1 0 26036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1667941163
transform 1 0 37812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1667941163
transform 1 0 33120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1667941163
transform 1 0 27968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0824_
timestamp 1667941163
transform 1 0 21804 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1667941163
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1667941163
transform 1 0 35604 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1667941163
transform 1 0 21988 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1667941163
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1667941163
transform 1 0 18768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1667941163
transform 1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1667941163
transform 1 0 30636 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1667941163
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1667941163
transform 1 0 31004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1667941163
transform 1 0 31924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1667941163
transform 1 0 37168 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1667941163
transform 1 0 36708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1667941163
transform 1 0 32292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1667941163
transform 1 0 33120 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1667941163
transform 1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1667941163
transform 1 0 19412 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1667941163
transform 1 0 18584 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _0843_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32476 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0844_
timestamp 1667941163
transform 1 0 32752 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0845_
timestamp 1667941163
transform 1 0 33488 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0846_
timestamp 1667941163
transform 1 0 34960 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0847_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0848_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30912 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0849_
timestamp 1667941163
transform 1 0 31372 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0850_
timestamp 1667941163
transform 1 0 20700 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0851_
timestamp 1667941163
transform 1 0 24840 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0852_
timestamp 1667941163
transform 1 0 22540 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0853_
timestamp 1667941163
transform 1 0 22264 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0854_
timestamp 1667941163
transform 1 0 22264 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0855_
timestamp 1667941163
transform 1 0 15272 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0856_
timestamp 1667941163
transform 1 0 15640 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0857_
timestamp 1667941163
transform 1 0 15640 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0858_
timestamp 1667941163
transform 1 0 30728 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0859_
timestamp 1667941163
transform 1 0 14536 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0860_
timestamp 1667941163
transform 1 0 14536 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0861_
timestamp 1667941163
transform 1 0 16836 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0862_
timestamp 1667941163
transform 1 0 16836 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0863_
timestamp 1667941163
transform 1 0 15916 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0864_
timestamp 1667941163
transform 1 0 16836 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0865_
timestamp 1667941163
transform 1 0 27508 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0866_
timestamp 1667941163
transform 1 0 24748 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0867_
timestamp 1667941163
transform 1 0 20332 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0868_
timestamp 1667941163
transform 1 0 18308 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0869_
timestamp 1667941163
transform 1 0 18676 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0870_
timestamp 1667941163
transform 1 0 19228 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0871_
timestamp 1667941163
transform 1 0 15364 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0872_
timestamp 1667941163
transform 1 0 23184 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0873_
timestamp 1667941163
transform 1 0 22172 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0874_
timestamp 1667941163
transform 1 0 21804 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0875_
timestamp 1667941163
transform 1 0 31924 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0876_
timestamp 1667941163
transform 1 0 34868 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0877_
timestamp 1667941163
transform 1 0 34868 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0878_
timestamp 1667941163
transform 1 0 26036 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0879_
timestamp 1667941163
transform 1 0 21988 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0880_
timestamp 1667941163
transform 1 0 29716 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0881_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0882_
timestamp 1667941163
transform 1 0 18584 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0883_
timestamp 1667941163
transform 1 0 34500 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0884_
timestamp 1667941163
transform 1 0 34960 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0885_
timestamp 1667941163
transform 1 0 31004 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0886_
timestamp 1667941163
transform 1 0 32200 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0887_
timestamp 1667941163
transform 1 0 24748 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0888_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0889_
timestamp 1667941163
transform 1 0 33304 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0890_
timestamp 1667941163
transform 1 0 32292 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0891_
timestamp 1667941163
transform 1 0 18124 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0892_
timestamp 1667941163
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0893_
timestamp 1667941163
transform 1 0 14536 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0894_
timestamp 1667941163
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0895_
timestamp 1667941163
transform 1 0 16836 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0896_
timestamp 1667941163
transform 1 0 19596 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0897_
timestamp 1667941163
transform 1 0 16192 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0898_
timestamp 1667941163
transform 1 0 26680 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0899_
timestamp 1667941163
transform 1 0 27232 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0900_
timestamp 1667941163
transform 1 0 32752 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0901_
timestamp 1667941163
transform 1 0 29716 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0902_
timestamp 1667941163
transform 1 0 22632 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0903_
timestamp 1667941163
transform 1 0 23644 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0904_
timestamp 1667941163
transform 1 0 20608 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0905_
timestamp 1667941163
transform 1 0 17664 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0906_
timestamp 1667941163
transform 1 0 19320 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0907_
timestamp 1667941163
transform 1 0 20792 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0908_
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0909_
timestamp 1667941163
transform 1 0 15364 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0910_
timestamp 1667941163
transform 1 0 27140 0 -1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0911_
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0912_
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0913_
timestamp 1667941163
transform 1 0 20700 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0914_
timestamp 1667941163
transform 1 0 19596 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0915_
timestamp 1667941163
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0916_
timestamp 1667941163
transform 1 0 15088 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0917_
timestamp 1667941163
transform 1 0 19688 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0918_
timestamp 1667941163
transform 1 0 14536 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0919_
timestamp 1667941163
transform 1 0 19596 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0920_
timestamp 1667941163
transform 1 0 20424 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0921_
timestamp 1667941163
transform 1 0 18492 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0922_
timestamp 1667941163
transform 1 0 22540 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0923_
timestamp 1667941163
transform 1 0 31464 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1667941163
transform 1 0 32568 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1667941163
transform 1 0 25484 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0926_
timestamp 1667941163
transform 1 0 22080 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0927_
timestamp 1667941163
transform 1 0 25116 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0928_
timestamp 1667941163
transform 1 0 34868 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0929_
timestamp 1667941163
transform 1 0 29808 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0930_
timestamp 1667941163
transform 1 0 34132 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0931_
timestamp 1667941163
transform 1 0 32292 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0932_
timestamp 1667941163
transform 1 0 34868 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0933_
timestamp 1667941163
transform 1 0 32016 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0934_
timestamp 1667941163
transform 1 0 33488 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0935_
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0936_
timestamp 1667941163
transform 1 0 28428 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0937_
timestamp 1667941163
transform 1 0 19412 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0938_
timestamp 1667941163
transform 1 0 30084 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0939_
timestamp 1667941163
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0940_
timestamp 1667941163
transform 1 0 34868 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0941_
timestamp 1667941163
transform 1 0 33120 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0942_
timestamp 1667941163
transform 1 0 25760 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0943_
timestamp 1667941163
transform 1 0 28244 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0944_
timestamp 1667941163
transform 1 0 33672 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0945_
timestamp 1667941163
transform 1 0 14536 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0946_
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0947_
timestamp 1667941163
transform 1 0 18124 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _0948_
timestamp 1667941163
transform 1 0 17756 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0949_
timestamp 1667941163
transform 1 0 29348 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1667941163
transform 1 0 22908 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0951_
timestamp 1667941163
transform 1 0 29532 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _0952_
timestamp 1667941163
transform 1 0 30544 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0953_
timestamp 1667941163
transform 1 0 34868 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0954_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _0955_
timestamp 1667941163
transform 1 0 28612 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1667941163
transform 1 0 27140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1667941163
transform 1 0 27140 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0958_
timestamp 1667941163
transform 1 0 17664 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0959_
timestamp 1667941163
transform 1 0 15732 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _0960_
timestamp 1667941163
transform 1 0 19412 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1667941163
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1667941163
transform 1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0987_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1667941163
transform 1 0 13524 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1667941163
transform 1 0 32200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1667941163
transform 1 0 6532 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1667941163
transform 1 0 32752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1667941163
transform 1 0 36708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0994_
timestamp 1667941163
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1667941163
transform 1 0 35788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1667941163
transform 1 0 35972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1667941163
transform 1 0 35512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1667941163
transform 1 0 14352 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1667941163
transform 1 0 37720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1667941163
transform 1 0 29716 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1667941163
transform 1 0 30176 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1667941163
transform 1 0 37352 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1667941163
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1005_
timestamp 1667941163
transform 1 0 3956 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1667941163
transform 1 0 37352 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1667941163
transform 1 0 27876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1008_
timestamp 1667941163
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1667941163
transform 1 0 21160 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1667941163
transform 1 0 26128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1667941163
transform 1 0 1932 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1012_
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1667941163
transform 1 0 32292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1667941163
transform 1 0 37352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1015_
timestamp 1667941163
transform 1 0 19780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1016_
timestamp 1667941163
transform 1 0 22448 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1017_
timestamp 1667941163
transform 1 0 16836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1667941163
transform 1 0 35604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1019_
timestamp 1667941163
transform 1 0 31280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1667941163
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1667941163
transform 1 0 6532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1667941163
transform 1 0 5336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1667941163
transform 1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1025_
timestamp 1667941163
transform 1 0 4784 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1667941163
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1667941163
transform 1 0 37812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1028_
timestamp 1667941163
transform 1 0 13156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1667941163
transform 1 0 37996 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1667941163
transform 1 0 37076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1031_
timestamp 1667941163
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1667941163
transform 1 0 13248 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1667941163
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1667941163
transform 1 0 2300 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1667941163
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1667941163
transform 1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1667941163
transform 1 0 8004 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1667941163
transform 1 0 14628 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1039_
timestamp 1667941163
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1040_
timestamp 1667941163
transform 1 0 36708 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1667941163
transform 1 0 37352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1042_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1043_
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1044_
timestamp 1667941163
transform 1 0 37444 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1044__142 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1045_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27324 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1046_
timestamp 1667941163
transform 1 0 36248 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1047_
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1048_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30084 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1049_
timestamp 1667941163
transform 1 0 37168 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1050_
timestamp 1667941163
transform 1 0 35144 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1051_
timestamp 1667941163
transform 1 0 36248 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _1052_
timestamp 1667941163
transform 1 0 25944 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1053_
timestamp 1667941163
transform 1 0 24564 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1054_
timestamp 1667941163
transform 1 0 13156 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1055_
timestamp 1667941163
transform 1 0 12972 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1056_
timestamp 1667941163
transform 1 0 14352 0 1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1056__143
timestamp 1667941163
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1057_
timestamp 1667941163
transform 1 0 10028 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1058_
timestamp 1667941163
transform 1 0 21436 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1059_
timestamp 1667941163
transform 1 0 21712 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1060_
timestamp 1667941163
transform 1 0 11040 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1061_
timestamp 1667941163
transform 1 0 16836 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1062_
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1063_
timestamp 1667941163
transform 1 0 12604 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1064_
timestamp 1667941163
transform 1 0 11960 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1065_
timestamp 1667941163
transform 1 0 22816 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1066_
timestamp 1667941163
transform 1 0 12604 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1067_
timestamp 1667941163
transform 1 0 8372 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1068__144
timestamp 1667941163
transform 1 0 8372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1068_
timestamp 1667941163
transform 1 0 9016 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1069_
timestamp 1667941163
transform 1 0 27140 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1070_
timestamp 1667941163
transform 1 0 15364 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1071_
timestamp 1667941163
transform 1 0 19412 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1072_
timestamp 1667941163
transform 1 0 10396 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1073_
timestamp 1667941163
transform 1 0 8096 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1074_
timestamp 1667941163
transform 1 0 1564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_4  _1075_
timestamp 1667941163
transform 1 0 12788 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_8  _1076_
timestamp 1667941163
transform 1 0 28520 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1077_
timestamp 1667941163
transform 1 0 34868 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _1078_
timestamp 1667941163
transform 1 0 12880 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1079_
timestamp 1667941163
transform 1 0 6072 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1080__145
timestamp 1667941163
transform 1 0 8740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1080_
timestamp 1667941163
transform 1 0 9108 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1081_
timestamp 1667941163
transform 1 0 26864 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1082_
timestamp 1667941163
transform 1 0 27324 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1083_
timestamp 1667941163
transform 1 0 11684 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1084_
timestamp 1667941163
transform 1 0 22816 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1085_
timestamp 1667941163
transform 1 0 13248 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1086_
timestamp 1667941163
transform 1 0 9200 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1087_
timestamp 1667941163
transform 1 0 11960 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1088_
timestamp 1667941163
transform 1 0 1564 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1089_
timestamp 1667941163
transform 1 0 10028 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1090_
timestamp 1667941163
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1091_
timestamp 1667941163
transform 1 0 35604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1092_
timestamp 1667941163
transform 1 0 36064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1092__146
timestamp 1667941163
transform 1 0 36156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1093_
timestamp 1667941163
transform 1 0 12604 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1094_
timestamp 1667941163
transform 1 0 12144 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1095_
timestamp 1667941163
transform 1 0 10580 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1096_
timestamp 1667941163
transform 1 0 29256 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1097_
timestamp 1667941163
transform 1 0 30636 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1098_
timestamp 1667941163
transform 1 0 15916 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1099_
timestamp 1667941163
transform 1 0 33304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1100_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1101_
timestamp 1667941163
transform 1 0 24564 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1102_
timestamp 1667941163
transform 1 0 34868 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1103_
timestamp 1667941163
transform 1 0 30360 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1104_
timestamp 1667941163
transform 1 0 30636 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1104__147
timestamp 1667941163
transform 1 0 31280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1105_
timestamp 1667941163
transform 1 0 26312 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1106_
timestamp 1667941163
transform 1 0 4324 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1107_
timestamp 1667941163
transform 1 0 15180 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1108_
timestamp 1667941163
transform 1 0 22816 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1109_
timestamp 1667941163
transform 1 0 14536 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1110_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1111_
timestamp 1667941163
transform 1 0 34868 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1112_
timestamp 1667941163
transform 1 0 33212 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1113_
timestamp 1667941163
transform 1 0 33120 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1114_
timestamp 1667941163
transform 1 0 9660 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1115_
timestamp 1667941163
transform 1 0 9568 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1116__148
timestamp 1667941163
transform 1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1116_
timestamp 1667941163
transform 1 0 21988 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1117_
timestamp 1667941163
transform 1 0 8004 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1118_
timestamp 1667941163
transform 1 0 8648 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1119_
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1120_
timestamp 1667941163
transform 1 0 12144 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1121_
timestamp 1667941163
transform 1 0 10212 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1122_
timestamp 1667941163
transform 1 0 9568 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1123_
timestamp 1667941163
transform 1 0 15180 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1124_
timestamp 1667941163
transform 1 0 10396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1125_
timestamp 1667941163
transform 1 0 12052 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1126_
timestamp 1667941163
transform 1 0 31004 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1127_
timestamp 1667941163
transform 1 0 32292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1128_
timestamp 1667941163
transform 1 0 16836 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1129__149
timestamp 1667941163
transform 1 0 21252 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1129_
timestamp 1667941163
transform 1 0 21988 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1130_
timestamp 1667941163
transform 1 0 11684 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1131_
timestamp 1667941163
transform 1 0 10948 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1132_
timestamp 1667941163
transform 1 0 27508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1133_
timestamp 1667941163
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1134_
timestamp 1667941163
transform 1 0 30084 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1135_
timestamp 1667941163
transform 1 0 27600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1136_
timestamp 1667941163
transform 1 0 19872 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1137_
timestamp 1667941163
transform 1 0 24564 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1138_
timestamp 1667941163
transform 1 0 10212 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1139_
timestamp 1667941163
transform 1 0 12972 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1140_
timestamp 1667941163
transform 1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1141__150
timestamp 1667941163
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1141_
timestamp 1667941163
transform 1 0 10304 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1142_
timestamp 1667941163
transform 1 0 7084 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1143_
timestamp 1667941163
transform 1 0 9108 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1144_
timestamp 1667941163
transform 1 0 7360 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1145_
timestamp 1667941163
transform 1 0 7912 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1146_
timestamp 1667941163
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1147_
timestamp 1667941163
transform 1 0 18308 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1148_
timestamp 1667941163
transform 1 0 9384 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1149_
timestamp 1667941163
transform 1 0 2944 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1150_
timestamp 1667941163
transform 1 0 35788 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1151__151
timestamp 1667941163
transform 1 0 35604 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1151_
timestamp 1667941163
transform 1 0 35604 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1152_
timestamp 1667941163
transform 1 0 12880 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1153_
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  _1154_
timestamp 1667941163
transform 1 0 15180 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1155_
timestamp 1667941163
transform 1 0 11316 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1156_
timestamp 1667941163
transform 1 0 11684 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1157__152
timestamp 1667941163
transform 1 0 13248 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1157_
timestamp 1667941163
transform 1 0 12972 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1158_
timestamp 1667941163
transform 1 0 9936 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1159_
timestamp 1667941163
transform 1 0 9200 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1160_
timestamp 1667941163
transform 1 0 13432 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1161_
timestamp 1667941163
transform 1 0 12052 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1162_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23368 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1163_
timestamp 1667941163
transform 1 0 30360 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1164_
timestamp 1667941163
transform 1 0 29992 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1164__153
timestamp 1667941163
transform 1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1165_
timestamp 1667941163
transform 1 0 18124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1166_
timestamp 1667941163
transform 1 0 17664 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1167_
timestamp 1667941163
transform 1 0 29716 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1168_
timestamp 1667941163
transform 1 0 28060 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1169_
timestamp 1667941163
transform 1 0 24840 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1170_
timestamp 1667941163
transform 1 0 12880 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1171_
timestamp 1667941163
transform 1 0 9292 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1172_
timestamp 1667941163
transform 1 0 25484 0 -1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  _1172__154
timestamp 1667941163
transform 1 0 25944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1173_
timestamp 1667941163
transform 1 0 34408 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1174_
timestamp 1667941163
transform 1 0 34868 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1175_
timestamp 1667941163
transform 1 0 9476 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1176_
timestamp 1667941163
transform 1 0 31648 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1177_
timestamp 1667941163
transform 1 0 32568 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1178_
timestamp 1667941163
transform 1 0 29716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1179__155
timestamp 1667941163
transform 1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1179_
timestamp 1667941163
transform 1 0 28888 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1180_
timestamp 1667941163
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1181_
timestamp 1667941163
transform 1 0 30912 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1182_
timestamp 1667941163
transform 1 0 24564 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1183_
timestamp 1667941163
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1184_
timestamp 1667941163
transform 1 0 12696 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1185_
timestamp 1667941163
transform 1 0 9568 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1185__156
timestamp 1667941163
transform 1 0 9568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1186_
timestamp 1667941163
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1187_
timestamp 1667941163
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1188_
timestamp 1667941163
transform 1 0 10212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1189_
timestamp 1667941163
transform 1 0 22448 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1190_
timestamp 1667941163
transform 1 0 20332 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1191__157
timestamp 1667941163
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1191_
timestamp 1667941163
transform 1 0 15732 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1192_
timestamp 1667941163
transform 1 0 14260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1193_
timestamp 1667941163
transform 1 0 21068 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1194_
timestamp 1667941163
transform 1 0 15180 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1195_
timestamp 1667941163
transform 1 0 21988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1196_
timestamp 1667941163
transform 1 0 33580 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1197__158
timestamp 1667941163
transform 1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1197_
timestamp 1667941163
transform 1 0 34132 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1198_
timestamp 1667941163
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1199_
timestamp 1667941163
transform 1 0 28336 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1200_
timestamp 1667941163
transform 1 0 32660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1201_
timestamp 1667941163
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1202_
timestamp 1667941163
transform 1 0 26312 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1203_
timestamp 1667941163
transform 1 0 19964 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1203__159
timestamp 1667941163
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1204_
timestamp 1667941163
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1667941163
transform 1 0 29072 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1206_
timestamp 1667941163
transform 1 0 20792 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1667941163
transform 1 0 31188 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1208_
timestamp 1667941163
transform 1 0 6808 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1209__160
timestamp 1667941163
transform 1 0 5428 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1667941163
transform 1 0 5336 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1667941163
transform 1 0 9108 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1667941163
transform 1 0 7912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1667941163
transform 1 0 6808 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1667941163
transform 1 0 7268 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1214_
timestamp 1667941163
transform 1 0 6532 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1215__161
timestamp 1667941163
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1667941163
transform 1 0 4416 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1216_
timestamp 1667941163
transform 1 0 9108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _1217_
timestamp 1667941163
transform 1 0 9108 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1667941163
transform 1 0 8648 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1220__162
timestamp 1667941163
transform 1 0 36064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1220_
timestamp 1667941163
transform 1 0 34592 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1667941163
transform 1 0 27232 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1222_
timestamp 1667941163
transform 1 0 30176 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1223_
timestamp 1667941163
transform 1 0 28336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1224__163
timestamp 1667941163
transform 1 0 35512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1224_
timestamp 1667941163
transform 1 0 34684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1225_
timestamp 1667941163
transform 1 0 19872 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1226_
timestamp 1667941163
transform 1 0 30452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1227_
timestamp 1667941163
transform 1 0 20700 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1228_
timestamp 1667941163
transform 1 0 37076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _1228__164
timestamp 1667941163
transform 1 0 35788 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _1229_
timestamp 1667941163
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1230_
timestamp 1667941163
transform 1 0 34224 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1231_
timestamp 1667941163
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1232_
timestamp 1667941163
transform 1 0 12420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1232__165
timestamp 1667941163
transform 1 0 12420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _1233_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1234_
timestamp 1667941163
transform 1 0 22448 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1235_
timestamp 1667941163
transform 1 0 10672 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1236_
timestamp 1667941163
transform 1 0 10028 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1237_
timestamp 1667941163
transform 1 0 23460 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_2  _1238_
timestamp 1667941163
transform 1 0 25208 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1239_
timestamp 1667941163
transform 1 0 14260 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _1240_
timestamp 1667941163
transform 1 0 27416 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _1241_
timestamp 1667941163
transform 1 0 17480 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_2  _1242_
timestamp 1667941163
transform 1 0 23276 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25668 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk
timestamp 1667941163
transform 1 0 17664 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1667941163
transform 1 0 16836 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1667941163
transform 1 0 20516 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1667941163
transform 1 0 17940 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1667941163
transform 1 0 17940 0 1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1667941163
transform 1 0 23092 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1667941163
transform 1 0 22908 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1667941163
transform 1 0 28244 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1667941163
transform 1 0 27600 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1667941163
transform 1 0 33396 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1667941163
transform 1 0 29072 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1667941163
transform 1 0 29992 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1667941163
transform 1 0 33396 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1667941163
transform 1 0 32936 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1667941163
transform 1 0 35236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1667941163
transform 1 0 1564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1667941163
transform 1 0 1564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1667941163
transform 1 0 17940 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1667941163
transform 1 0 3956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 12880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1667941163
transform 1 0 25760 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1667941163
transform 1 0 6532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1667941163
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1667941163
transform 1 0 8372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1667941163
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1667941163
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1667941163
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1667941163
transform 1 0 28520 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1667941163
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1667941163
transform 1 0 38088 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1667941163
transform 1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1667941163
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1667941163
transform 1 0 14996 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1667941163
transform 1 0 38088 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1667941163
transform 1 0 32936 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1667941163
transform 1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1667941163
transform 1 0 36616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1667941163
transform 1 0 37444 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1667941163
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1667941163
transform 1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1667941163
transform 1 0 38088 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1667941163
transform 1 0 9108 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1667941163
transform 1 0 11684 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1667941163
transform 1 0 22724 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1667941163
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1667941163
transform 1 0 3128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1667941163
transform 1 0 37996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1667941163
transform 1 0 3956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1667941163
transform 1 0 36708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1667941163
transform 1 0 1564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1667941163
transform 1 0 37444 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1667941163
transform 1 0 1564 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1667941163
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1667941163
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1667941163
transform 1 0 16836 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1667941163
transform 1 0 1564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1667941163
transform 1 0 2024 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1667941163
transform 1 0 1564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1667941163
transform 1 0 3956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1667941163
transform 1 0 37444 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1667941163
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1667941163
transform 1 0 1564 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1667941163
transform 1 0 23184 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1667941163
transform 1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1667941163
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1667941163
transform 1 0 30912 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1667941163
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1667941163
transform 1 0 14904 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1667941163
transform 1 0 37444 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1667941163
transform 1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1667941163
transform 1 0 34132 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1667941163
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1667941163
transform 1 0 1564 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1667941163
transform 1 0 38088 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1667941163
transform 1 0 1564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1667941163
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1667941163
transform 1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1667941163
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1667941163
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1667941163
transform 1 0 38088 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1667941163
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1667941163
transform 1 0 28980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1667941163
transform 1 0 2208 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1667941163
transform 1 0 7176 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1667941163
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output84 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1667941163
transform 1 0 36156 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1667941163
transform 1 0 37996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1667941163
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1667941163
transform 1 0 1564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1667941163
transform 1 0 36616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1667941163
transform 1 0 37996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1667941163
transform 1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1667941163
transform 1 0 18584 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1667941163
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1667941163
transform 1 0 32292 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1667941163
transform 1 0 34868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1667941163
transform 1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1667941163
transform 1 0 16008 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1667941163
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1667941163
transform 1 0 37996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1667941163
transform 1 0 37996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1667941163
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1667941163
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1667941163
transform 1 0 33028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1667941163
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1667941163
transform 1 0 30360 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1667941163
transform 1 0 37996 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1667941163
transform 1 0 27140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1667941163
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1667941163
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1667941163
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1667941163
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1667941163
transform 1 0 1564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1667941163
transform 1 0 37996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1667941163
transform 1 0 37996 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1667941163
transform 1 0 16836 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1667941163
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1667941163
transform 1 0 37996 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1667941163
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1667941163
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1667941163
transform 1 0 37996 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1667941163
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1667941163
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1667941163
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1667941163
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1667941163
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1667941163
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1667941163
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1667941163
transform 1 0 23460 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1667941163
transform 1 0 1564 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1667941163
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1667941163
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1667941163
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1667941163
transform 1 0 21988 0 1 36992
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 19048 800 19168 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 0 nsew signal input
flabel metal3 s 200 7488 800 7608 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 1 nsew signal input
flabel metal2 s 5170 39200 5226 39800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 2 nsew signal input
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 3 nsew signal input
flabel metal2 s 35438 200 35494 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 4 nsew signal input
flabel metal2 s 25778 200 25834 800 0 FreeSans 224 90 0 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 5 nsew signal input
flabel metal3 s 200 22448 800 22568 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 6 nsew signal input
flabel metal3 s 200 6808 800 6928 0 FreeSans 480 0 0 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 7 nsew signal input
flabel metal2 s 18050 39200 18106 39800 0 FreeSans 224 90 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 8 nsew signal input
flabel metal3 s 200 38768 800 38888 0 FreeSans 480 0 0 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 9 nsew signal input
flabel metal2 s 12898 200 12954 800 0 FreeSans 224 90 0 0 ccff_head
port 10 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 ccff_tail
port 11 nsew signal tristate
flabel metal2 s 25778 39200 25834 39800 0 FreeSans 224 90 0 0 chanx_right_in[0]
port 12 nsew signal input
flabel metal2 s 5814 39200 5870 39800 0 FreeSans 224 90 0 0 chanx_right_in[10]
port 13 nsew signal input
flabel metal2 s 24490 200 24546 800 0 FreeSans 224 90 0 0 chanx_right_in[11]
port 14 nsew signal input
flabel metal2 s 9034 39200 9090 39800 0 FreeSans 224 90 0 0 chanx_right_in[12]
port 15 nsew signal input
flabel metal2 s 19982 200 20038 800 0 FreeSans 224 90 0 0 chanx_right_in[13]
port 16 nsew signal input
flabel metal3 s 200 17008 800 17128 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 17 nsew signal input
flabel metal3 s 200 2048 800 2168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 18 nsew signal input
flabel metal2 s 27710 39200 27766 39800 0 FreeSans 224 90 0 0 chanx_right_in[16]
port 19 nsew signal input
flabel metal2 s 11610 200 11666 800 0 FreeSans 224 90 0 0 chanx_right_in[17]
port 20 nsew signal input
flabel metal3 s 39200 31968 39800 32088 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 21 nsew signal input
flabel metal3 s 39200 27208 39800 27328 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 22 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 chanx_right_in[2]
port 23 nsew signal input
flabel metal3 s 200 688 800 808 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 24 nsew signal input
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 25 nsew signal input
flabel metal2 s 14830 39200 14886 39800 0 FreeSans 224 90 0 0 chanx_right_in[5]
port 26 nsew signal input
flabel metal3 s 39200 30608 39800 30728 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 27 nsew signal input
flabel metal3 s 39200 28568 39800 28688 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 28 nsew signal input
flabel metal2 s 32218 39200 32274 39800 0 FreeSans 224 90 0 0 chanx_right_in[8]
port 29 nsew signal input
flabel metal2 s 18050 200 18106 800 0 FreeSans 224 90 0 0 chanx_right_in[9]
port 30 nsew signal input
flabel metal2 s 36082 39200 36138 39800 0 FreeSans 224 90 0 0 chanx_right_out[0]
port 31 nsew signal tristate
flabel metal3 s 39200 12248 39800 12368 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 32 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 chanx_right_out[11]
port 33 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 34 nsew signal tristate
flabel metal3 s 200 15648 800 15768 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 35 nsew signal tristate
flabel metal3 s 39200 2048 39800 2168 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 36 nsew signal tristate
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 chanx_right_out[15]
port 37 nsew signal tristate
flabel metal3 s 39200 35368 39800 35488 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 38 nsew signal tristate
flabel metal3 s 39200 8 39800 128 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 39 nsew signal tristate
flabel metal2 s 19338 39200 19394 39800 0 FreeSans 224 90 0 0 chanx_right_out[18]
port 40 nsew signal tristate
flabel metal2 s 34150 200 34206 800 0 FreeSans 224 90 0 0 chanx_right_out[1]
port 41 nsew signal tristate
flabel metal2 s 30930 39200 30986 39800 0 FreeSans 224 90 0 0 chanx_right_out[2]
port 42 nsew signal tristate
flabel metal2 s 34150 39200 34206 39800 0 FreeSans 224 90 0 0 chanx_right_out[3]
port 43 nsew signal tristate
flabel metal3 s 39200 37408 39800 37528 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 44 nsew signal tristate
flabel metal2 s 16118 39200 16174 39800 0 FreeSans 224 90 0 0 chanx_right_out[5]
port 45 nsew signal tristate
flabel metal3 s 39200 10888 39800 11008 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 46 nsew signal tristate
flabel metal3 s 39200 13608 39800 13728 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 47 nsew signal tristate
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 48 nsew signal tristate
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 chanx_right_out[9]
port 49 nsew signal tristate
flabel metal3 s 39200 38768 39800 38888 0 FreeSans 480 0 0 0 chany_bottom_in[0]
port 50 nsew signal input
flabel metal3 s 39200 32648 39800 32768 0 FreeSans 480 0 0 0 chany_bottom_in[10]
port 51 nsew signal input
flabel metal2 s 24490 39200 24546 39800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 52 nsew signal input
flabel metal2 s 12254 39200 12310 39800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 53 nsew signal input
flabel metal3 s 39200 23808 39800 23928 0 FreeSans 480 0 0 0 chany_bottom_in[13]
port 54 nsew signal input
flabel metal2 s 8390 39200 8446 39800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 55 nsew signal input
flabel metal2 s 11610 39200 11666 39800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 56 nsew signal input
flabel metal2 s 22558 39200 22614 39800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 57 nsew signal input
flabel metal2 s 10322 200 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 58 nsew signal input
flabel metal2 s 2594 39200 2650 39800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 59 nsew signal input
flabel metal3 s 39200 14968 39800 15088 0 FreeSans 480 0 0 0 chany_bottom_in[1]
port 60 nsew signal input
flabel metal2 s 3882 39200 3938 39800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 61 nsew signal input
flabel metal3 s 39200 688 39800 808 0 FreeSans 480 0 0 0 chany_bottom_in[3]
port 62 nsew signal input
flabel metal3 s 200 14288 800 14408 0 FreeSans 480 0 0 0 chany_bottom_in[4]
port 63 nsew signal input
flabel metal3 s 39200 7488 39800 7608 0 FreeSans 480 0 0 0 chany_bottom_in[5]
port 64 nsew signal input
flabel metal3 s 200 28568 800 28688 0 FreeSans 480 0 0 0 chany_bottom_in[6]
port 65 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 66 nsew signal input
flabel metal3 s 200 21088 800 21208 0 FreeSans 480 0 0 0 chany_bottom_in[8]
port 67 nsew signal input
flabel metal2 s 16118 200 16174 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 68 nsew signal input
flabel metal3 s 200 24488 800 24608 0 FreeSans 480 0 0 0 chany_bottom_out[0]
port 69 nsew signal tristate
flabel metal2 s 32862 39200 32918 39800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 70 nsew signal tristate
flabel metal3 s 200 32648 800 32768 0 FreeSans 480 0 0 0 chany_bottom_out[11]
port 71 nsew signal tristate
flabel metal2 s 30286 200 30342 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 72 nsew signal tristate
flabel metal3 s 39200 25168 39800 25288 0 FreeSans 480 0 0 0 chany_bottom_out[13]
port 73 nsew signal tristate
flabel metal3 s 39200 5448 39800 5568 0 FreeSans 480 0 0 0 chany_bottom_out[14]
port 74 nsew signal tristate
flabel metal2 s 26422 39200 26478 39800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 75 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 76 nsew signal tristate
flabel metal2 s 37370 39200 37426 39800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 77 nsew signal tristate
flabel metal2 s 662 200 718 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 78 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 79 nsew signal tristate
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 80 nsew signal tristate
flabel metal3 s 200 13608 800 13728 0 FreeSans 480 0 0 0 chany_bottom_out[3]
port 81 nsew signal tristate
flabel metal3 s 39200 21768 39800 21888 0 FreeSans 480 0 0 0 chany_bottom_out[4]
port 82 nsew signal tristate
flabel metal3 s 39200 15648 39800 15768 0 FreeSans 480 0 0 0 chany_bottom_out[5]
port 83 nsew signal tristate
flabel metal2 s 16762 39200 16818 39800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 84 nsew signal tristate
flabel metal2 s 3238 200 3294 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 85 nsew signal tristate
flabel metal3 s 39200 3408 39800 3528 0 FreeSans 480 0 0 0 chany_bottom_out[8]
port 86 nsew signal tristate
flabel metal3 s 39200 17008 39800 17128 0 FreeSans 480 0 0 0 chany_bottom_out[9]
port 87 nsew signal tristate
flabel metal3 s 200 27208 800 27328 0 FreeSans 480 0 0 0 chany_top_in[0]
port 88 nsew signal input
flabel metal2 s 1950 39200 2006 39800 0 FreeSans 224 90 0 0 chany_top_in[10]
port 89 nsew signal input
flabel metal3 s 200 25848 800 25968 0 FreeSans 480 0 0 0 chany_top_in[11]
port 90 nsew signal input
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 chany_top_in[12]
port 91 nsew signal input
flabel metal3 s 200 39448 800 39568 0 FreeSans 480 0 0 0 chany_top_in[13]
port 92 nsew signal input
flabel metal2 s 38658 39200 38714 39800 0 FreeSans 224 90 0 0 chany_top_in[14]
port 93 nsew signal input
flabel metal2 s 8390 200 8446 800 0 FreeSans 224 90 0 0 chany_top_in[15]
port 94 nsew signal input
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 chany_top_in[16]
port 95 nsew signal input
flabel metal2 s 23202 200 23258 800 0 FreeSans 224 90 0 0 chany_top_in[17]
port 96 nsew signal input
flabel metal2 s 37370 200 37426 800 0 FreeSans 224 90 0 0 chany_top_in[18]
port 97 nsew signal input
flabel metal2 s 13542 39200 13598 39800 0 FreeSans 224 90 0 0 chany_top_in[1]
port 98 nsew signal input
flabel metal2 s 30930 200 30986 800 0 FreeSans 224 90 0 0 chany_top_in[2]
port 99 nsew signal input
flabel metal2 s 3882 200 3938 800 0 FreeSans 224 90 0 0 chany_top_in[3]
port 100 nsew signal input
flabel metal2 s 14830 200 14886 800 0 FreeSans 224 90 0 0 chany_top_in[4]
port 101 nsew signal input
flabel metal3 s 39200 4088 39800 4208 0 FreeSans 480 0 0 0 chany_top_in[5]
port 102 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 chany_top_in[6]
port 103 nsew signal input
flabel metal3 s 39200 20408 39800 20528 0 FreeSans 480 0 0 0 chany_top_in[7]
port 104 nsew signal input
flabel metal2 s 32218 200 32274 800 0 FreeSans 224 90 0 0 chany_top_in[8]
port 105 nsew signal input
flabel metal3 s 200 23808 800 23928 0 FreeSans 480 0 0 0 chany_top_in[9]
port 106 nsew signal input
flabel metal3 s 39200 10208 39800 10328 0 FreeSans 480 0 0 0 chany_top_out[0]
port 107 nsew signal tristate
flabel metal3 s 200 31968 800 32088 0 FreeSans 480 0 0 0 chany_top_out[10]
port 108 nsew signal tristate
flabel metal3 s 39200 22448 39800 22568 0 FreeSans 480 0 0 0 chany_top_out[11]
port 109 nsew signal tristate
flabel metal3 s 39200 34008 39800 34128 0 FreeSans 480 0 0 0 chany_top_out[12]
port 110 nsew signal tristate
flabel metal2 s 36726 200 36782 800 0 FreeSans 224 90 0 0 chany_top_out[13]
port 111 nsew signal tristate
flabel metal3 s 39200 36048 39800 36168 0 FreeSans 480 0 0 0 chany_top_out[14]
port 112 nsew signal tristate
flabel metal3 s 200 12248 800 12368 0 FreeSans 480 0 0 0 chany_top_out[15]
port 113 nsew signal tristate
flabel metal3 s 200 34008 800 34128 0 FreeSans 480 0 0 0 chany_top_out[16]
port 114 nsew signal tristate
flabel metal3 s 200 3408 800 3528 0 FreeSans 480 0 0 0 chany_top_out[17]
port 115 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 chany_top_out[18]
port 116 nsew signal tristate
flabel metal3 s 200 4088 800 4208 0 FreeSans 480 0 0 0 chany_top_out[1]
port 117 nsew signal tristate
flabel metal3 s 200 37408 800 37528 0 FreeSans 480 0 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 23202 39200 23258 39800 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6458 200 6514 800 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 1950 200 2006 800 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal3 s 200 8848 800 8968 0 FreeSans 480 0 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 21270 39200 21326 39800 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 pReset
port 126 nsew signal input
flabel metal2 s 35438 39200 35494 39800 0 FreeSans 224 90 0 0 prog_clk
port 127 nsew signal input
flabel metal3 s 39200 6808 39800 6928 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 128 nsew signal input
flabel metal3 s 200 36048 800 36168 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 129 nsew signal input
flabel metal3 s 200 10888 800 11008 0 FreeSans 480 0 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
port 130 nsew signal input
flabel metal2 s 7102 200 7158 800 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
port 131 nsew signal input
flabel metal2 s 13542 200 13598 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal2 s 21270 200 21326 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 39200 25848 39800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal2 s 22558 200 22614 800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
port 136 nsew signal input
flabel metal2 s 28998 39200 29054 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
port 137 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
port 138 nsew signal input
flabel metal2 s 7102 39200 7158 39800 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
port 139 nsew signal input
flabel metal2 s 27066 200 27122 800 0 FreeSans 224 90 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
port 140 nsew signal input
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
port 141 nsew signal input
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 142 nsew signal bidirectional
flabel metal3 s 39200 18368 39800 18488 0 FreeSans 480 0 0 0 vssd1
port 143 nsew signal bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 143 nsew signal bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal1 36662 22202 36662 22202 0 _0000_
rlabel metal1 34546 19482 34546 19482 0 _0001_
rlabel metal1 18768 21114 18768 21114 0 _0002_
rlabel metal1 19550 20298 19550 20298 0 _0003_
rlabel metal1 17020 21590 17020 21590 0 _0004_
rlabel metal1 16981 23018 16981 23018 0 _0005_
rlabel metal1 17894 20570 17894 20570 0 _0006_
rlabel metal1 19044 19482 19044 19482 0 _0007_
rlabel metal1 18446 18938 18446 18938 0 _0008_
rlabel metal1 29072 21114 29072 21114 0 _0009_
rlabel metal2 28336 19958 28336 19958 0 _0010_
rlabel metal1 36248 20570 36248 20570 0 _0011_
rlabel metal1 30544 21658 30544 21658 0 _0012_
rlabel metal1 24932 21658 24932 21658 0 _0013_
rlabel metal1 25760 20570 25760 20570 0 _0014_
rlabel metal2 21160 25806 21160 25806 0 _0015_
rlabel metal1 11914 33626 11914 33626 0 _0016_
rlabel metal2 20102 35462 20102 35462 0 _0017_
rlabel metal2 12098 33745 12098 33745 0 _0018_
rlabel metal1 12880 33422 12880 33422 0 _0019_
rlabel metal1 14720 29478 14720 29478 0 _0020_
rlabel via2 31970 20485 31970 20485 0 _0021_
rlabel metal3 35719 34612 35719 34612 0 _0022_
rlabel metal1 32844 20570 32844 20570 0 _0023_
rlabel via2 26358 18955 26358 18955 0 _0024_
rlabel metal1 17756 19482 17756 19482 0 _0025_
rlabel metal2 14950 32776 14950 32776 0 _0026_
rlabel metal1 12466 32776 12466 32776 0 _0027_
rlabel metal2 21114 32198 21114 32198 0 _0028_
rlabel via2 10994 34731 10994 34731 0 _0029_
rlabel metal1 19734 33864 19734 33864 0 _0030_
rlabel metal1 17250 36312 17250 36312 0 _0031_
rlabel metal1 19918 34537 19918 34537 0 _0032_
rlabel metal1 27186 19482 27186 19482 0 _0033_
rlabel metal1 37996 20570 37996 20570 0 _0034_
rlabel metal1 37444 20570 37444 20570 0 _0035_
rlabel metal1 27876 19958 27876 19958 0 _0036_
rlabel metal1 25254 19482 25254 19482 0 _0037_
rlabel metal1 27600 20026 27600 20026 0 _0038_
rlabel metal1 36623 34986 36623 34986 0 _0039_
rlabel via2 29210 17323 29210 17323 0 _0040_
rlabel metal1 36117 36822 36117 36822 0 _0041_
rlabel metal1 35466 34680 35466 34680 0 _0042_
rlabel metal2 35972 33524 35972 33524 0 _0043_
rlabel metal1 33541 31790 33541 31790 0 _0044_
rlabel metal1 38272 17850 38272 17850 0 _0045_
rlabel metal1 32752 19414 32752 19414 0 _0046_
rlabel via2 28658 17867 28658 17867 0 _0047_
rlabel metal1 23598 18802 23598 18802 0 _0048_
rlabel metal1 33764 18598 33764 18598 0 _0049_
rlabel metal1 26082 19482 26082 19482 0 _0050_
rlabel metal1 37904 18394 37904 18394 0 _0051_
rlabel metal1 33948 18870 33948 18870 0 _0052_
rlabel metal1 27600 18326 27600 18326 0 _0053_
rlabel metal1 29769 24786 29769 24786 0 _0054_
rlabel metal1 35473 25942 35473 25942 0 _0055_
rlabel metal1 19642 29036 19642 29036 0 _0056_
rlabel metal1 21351 23018 21351 23018 0 _0057_
rlabel metal2 18906 23800 18906 23800 0 _0058_
rlabel metal1 20976 27098 20976 27098 0 _0059_
rlabel metal2 30774 23494 30774 23494 0 _0060_
rlabel metal1 25576 20502 25576 20502 0 _0061_
rlabel metal2 31142 21325 31142 21325 0 _0062_
rlabel metal1 31970 21114 31970 21114 0 _0063_
rlabel metal1 38456 17782 38456 17782 0 _0064_
rlabel metal1 36938 18394 36938 18394 0 _0065_
rlabel metal1 31372 19482 31372 19482 0 _0066_
rlabel metal2 33258 19584 33258 19584 0 _0067_
rlabel metal1 28060 17850 28060 17850 0 _0068_
rlabel metal1 19504 21114 19504 21114 0 _0069_
rlabel metal2 18722 22610 18722 22610 0 _0070_
rlabel metal2 20746 22916 20746 22916 0 _0071_
rlabel metal1 35512 21046 35512 21046 0 _0072_
rlabel metal1 36248 21658 36248 21658 0 _0073_
rlabel metal1 37628 21114 37628 21114 0 _0074_
rlabel metal1 37306 21590 37306 21590 0 _0075_
rlabel metal1 36800 20026 36800 20026 0 _0076_
rlabel metal1 33863 36074 33863 36074 0 _0077_
rlabel metal1 34270 18326 34270 18326 0 _0078_
rlabel metal1 22678 20026 22678 20026 0 _0079_
rlabel via2 26082 18411 26082 18411 0 _0080_
rlabel metal1 24387 36822 24387 36822 0 _0081_
rlabel metal1 19826 22474 19826 22474 0 _0082_
rlabel metal1 21436 31790 21436 31790 0 _0083_
rlabel metal1 17066 21318 17066 21318 0 _0084_
rlabel metal1 14766 20026 14766 20026 0 _0085_
rlabel metal1 15870 27336 15870 27336 0 _0086_
rlabel metal1 29256 20502 29256 20502 0 _0087_
rlabel metal1 14759 27030 14759 27030 0 _0088_
rlabel metal1 14122 22746 14122 22746 0 _0089_
rlabel metal1 17020 22202 17020 22202 0 _0090_
rlabel metal1 17250 19482 17250 19482 0 _0091_
rlabel metal2 16698 35802 16698 35802 0 _0092_
rlabel metal2 13110 33796 13110 33796 0 _0093_
rlabel metal1 28704 20570 28704 20570 0 _0094_
rlabel metal2 28566 20553 28566 20553 0 _0095_
rlabel metal1 14950 29784 14950 29784 0 _0096_
rlabel metal2 12834 30464 12834 30464 0 _0097_
rlabel metal2 16146 30736 16146 30736 0 _0098_
rlabel metal1 16238 34408 16238 34408 0 _0099_
rlabel metal2 9062 34816 9062 34816 0 _0100_
rlabel via2 28934 20043 28934 20043 0 _0101_
rlabel metal1 24065 33898 24065 33898 0 _0102_
rlabel metal2 21942 24446 21942 24446 0 _0103_
rlabel metal1 34822 19414 34822 19414 0 _0104_
rlabel metal1 35834 20570 35834 20570 0 _0105_
rlabel metal2 36202 22610 36202 22610 0 _0106_
rlabel metal1 30038 18938 30038 18938 0 _0107_
rlabel metal2 21344 21284 21344 21284 0 _0108_
rlabel metal1 31333 29546 31333 29546 0 _0109_
rlabel metal1 28711 28118 28711 28118 0 _0110_
rlabel metal2 20608 28220 20608 28220 0 _0111_
rlabel metal1 36761 23766 36761 23766 0 _0112_
rlabel metal1 37037 22678 37037 22678 0 _0113_
rlabel metal1 35696 21114 35696 21114 0 _0114_
rlabel metal2 32338 20502 32338 20502 0 _0115_
rlabel metal1 26726 17306 26726 17306 0 _0116_
rlabel metal1 25530 17850 25530 17850 0 _0117_
rlabel metal1 35650 20332 35650 20332 0 _0118_
rlabel metal1 18170 20400 18170 20400 0 _0119_
rlabel metal1 18446 21522 18446 21522 0 _0120_
rlabel metal1 33028 20434 33028 20434 0 _0121_
rlabel metal1 19826 20536 19826 20536 0 _0122_
rlabel metal1 36110 18734 36110 18734 0 _0123_
rlabel metal2 37858 17952 37858 17952 0 _0124_
rlabel metal2 31970 21114 31970 21114 0 _0125_
rlabel metal2 31050 15878 31050 15878 0 _0126_
rlabel metal2 37950 9996 37950 9996 0 _0127_
rlabel metal2 19642 17850 19642 17850 0 _0128_
rlabel metal1 34224 12410 34224 12410 0 _0129_
rlabel metal1 27646 15130 27646 15130 0 _0130_
rlabel metal2 32982 12036 32982 12036 0 _0131_
rlabel metal2 7590 11322 7590 11322 0 _0132_
rlabel metal1 7176 19482 7176 19482 0 _0133_
rlabel metal1 5244 21522 5244 21522 0 _0134_
rlabel metal1 5198 28492 5198 28492 0 _0135_
rlabel metal1 7084 27438 7084 27438 0 _0136_
rlabel metal1 4738 24752 4738 24752 0 _0137_
rlabel metal2 32614 13430 32614 13430 0 _0138_
rlabel metal1 24794 13328 24794 13328 0 _0139_
rlabel metal1 19826 12410 19826 12410 0 _0140_
rlabel metal2 16330 15164 16330 15164 0 _0141_
rlabel metal2 35926 15300 35926 15300 0 _0142_
rlabel metal1 34730 13940 34730 13940 0 _0143_
rlabel metal2 14858 12988 14858 12988 0 _0144_
rlabel metal2 20378 9146 20378 9146 0 _0145_
rlabel metal1 15318 9520 15318 9520 0 _0146_
rlabel metal1 28612 12954 28612 12954 0 _0147_
rlabel metal1 12006 19822 12006 19822 0 _0148_
rlabel metal1 9246 18224 9246 18224 0 _0149_
rlabel metal2 24794 6970 24794 6970 0 _0150_
rlabel metal1 30130 11084 30130 11084 0 _0151_
rlabel metal2 28934 9078 28934 9078 0 _0152_
rlabel metal2 22724 16524 22724 16524 0 _0153_
rlabel metal1 32752 19346 32752 19346 0 _0154_
rlabel metal1 36662 19822 36662 19822 0 _0155_
rlabel metal1 20884 19346 20884 19346 0 _0156_
rlabel metal1 28474 20366 28474 20366 0 _0157_
rlabel metal2 37674 15674 37674 15674 0 _0158_
rlabel metal2 37122 14552 37122 14552 0 _0159_
rlabel metal1 36340 14518 36340 14518 0 _0160_
rlabel metal1 27600 32946 27600 32946 0 _0161_
rlabel metal2 36478 30940 36478 30940 0 _0162_
rlabel via2 15410 20995 15410 20995 0 _0163_
rlabel metal1 30176 34170 30176 34170 0 _0164_
rlabel metal1 36800 16150 36800 16150 0 _0165_
rlabel metal2 35374 17374 35374 17374 0 _0166_
rlabel metal1 36478 15368 36478 15368 0 _0167_
rlabel metal1 25806 16490 25806 16490 0 _0168_
rlabel metal1 24242 12070 24242 12070 0 _0169_
rlabel metal1 13892 31382 13892 31382 0 _0170_
rlabel metal1 14076 32742 14076 32742 0 _0171_
rlabel metal1 13662 36040 13662 36040 0 _0172_
rlabel metal1 10626 19414 10626 19414 0 _0173_
rlabel metal2 21666 14824 21666 14824 0 _0174_
rlabel metal2 22126 18904 22126 18904 0 _0175_
rlabel metal2 11270 30226 11270 30226 0 _0176_
rlabel metal1 16652 11866 16652 11866 0 _0177_
rlabel metal2 25346 17102 25346 17102 0 _0178_
rlabel metal1 13110 32810 13110 32810 0 _0179_
rlabel metal1 12190 28424 12190 28424 0 _0180_
rlabel metal1 23460 15334 23460 15334 0 _0181_
rlabel metal2 13846 26112 13846 26112 0 _0182_
rlabel metal1 9476 27030 9476 27030 0 _0183_
rlabel metal1 12282 20570 12282 20570 0 _0184_
rlabel metal1 26450 34170 26450 34170 0 _0185_
rlabel metal1 13018 34952 13018 34952 0 _0186_
rlabel metal1 17204 18666 17204 18666 0 _0187_
rlabel metal1 10350 35122 10350 35122 0 _0188_
rlabel metal2 8326 23902 8326 23902 0 _0189_
rlabel metal1 2116 35802 2116 35802 0 _0190_
rlabel metal2 14398 27846 14398 27846 0 _0191_
rlabel metal1 29164 18394 29164 18394 0 _0192_
rlabel metal1 34684 17578 34684 17578 0 _0193_
rlabel metal1 15042 27098 15042 27098 0 _0194_
rlabel metal1 8418 23834 8418 23834 0 _0195_
rlabel metal1 9338 25160 9338 25160 0 _0196_
rlabel metal2 27462 18530 27462 18530 0 _0197_
rlabel metal1 27278 31994 27278 31994 0 _0198_
rlabel metal2 8326 35190 8326 35190 0 _0199_
rlabel metal1 23460 17238 23460 17238 0 _0200_
rlabel metal1 14030 20502 14030 20502 0 _0201_
rlabel metal2 9430 22814 9430 22814 0 _0202_
rlabel metal1 12742 24786 12742 24786 0 _0203_
rlabel metal1 2024 36822 2024 36822 0 _0204_
rlabel metal1 10120 24854 10120 24854 0 _0205_
rlabel via1 35098 19771 35098 19771 0 _0206_
rlabel metal1 35006 13498 35006 13498 0 _0207_
rlabel metal1 36294 12920 36294 12920 0 _0208_
rlabel metal2 12834 31586 12834 31586 0 _0209_
rlabel metal1 19320 17306 19320 17306 0 _0210_
rlabel metal2 10810 30872 10810 30872 0 _0211_
rlabel metal2 29486 16286 29486 16286 0 _0212_
rlabel metal1 30682 15062 30682 15062 0 _0213_
rlabel metal1 15732 14314 15732 14314 0 _0214_
rlabel metal2 33534 17374 33534 17374 0 _0215_
rlabel metal1 27416 14994 27416 14994 0 _0216_
rlabel metal2 24794 14110 24794 14110 0 _0217_
rlabel metal1 34454 18938 34454 18938 0 _0218_
rlabel metal1 31280 14246 31280 14246 0 _0219_
rlabel metal2 31050 14348 31050 14348 0 _0220_
rlabel metal1 26910 17578 26910 17578 0 _0221_
rlabel metal1 4600 33558 4600 33558 0 _0222_
rlabel metal2 16790 20264 16790 20264 0 _0223_
rlabel metal1 23644 18938 23644 18938 0 _0224_
rlabel metal2 14766 23528 14766 23528 0 _0225_
rlabel metal2 29946 20264 29946 20264 0 _0226_
rlabel metal2 35098 21794 35098 21794 0 _0227_
rlabel metal2 32890 17000 32890 17000 0 _0228_
rlabel metal1 33580 20026 33580 20026 0 _0229_
rlabel metal1 11178 20808 11178 20808 0 _0230_
rlabel metal2 9798 23154 9798 23154 0 _0231_
rlabel metal2 22218 15232 22218 15232 0 _0232_
rlabel metal1 9108 31382 9108 31382 0 _0233_
rlabel metal2 8878 17374 8878 17374 0 _0234_
rlabel metal2 8786 19822 8786 19822 0 _0235_
rlabel metal1 12098 29274 12098 29274 0 _0236_
rlabel metal2 10442 16728 10442 16728 0 _0237_
rlabel metal1 11776 26010 11776 26010 0 _0238_
rlabel metal2 15410 19550 15410 19550 0 _0239_
rlabel metal2 11546 30056 11546 30056 0 _0240_
rlabel metal2 12282 19720 12282 19720 0 _0241_
rlabel metal2 31234 19278 31234 19278 0 _0242_
rlabel metal2 31326 18734 31326 18734 0 _0243_
rlabel metal2 17066 9758 17066 9758 0 _0244_
rlabel metal2 22218 9214 22218 9214 0 _0245_
rlabel metal2 11914 14110 11914 14110 0 _0246_
rlabel metal2 11178 17442 11178 17442 0 _0247_
rlabel metal2 27738 8670 27738 8670 0 _0248_
rlabel metal2 27370 11118 27370 11118 0 _0249_
rlabel metal1 30636 16218 30636 16218 0 _0250_
rlabel metal1 27048 15674 27048 15674 0 _0251_
rlabel metal2 20102 11934 20102 11934 0 _0252_
rlabel metal2 24794 9656 24794 9656 0 _0253_
rlabel metal1 10396 32538 10396 32538 0 _0254_
rlabel metal2 14858 30226 14858 30226 0 _0255_
rlabel metal2 14398 16286 14398 16286 0 _0256_
rlabel metal1 10580 18666 10580 18666 0 _0257_
rlabel metal2 7314 32606 7314 32606 0 _0258_
rlabel metal1 9522 21930 9522 21930 0 _0259_
rlabel metal2 7590 21352 7590 21352 0 _0260_
rlabel metal2 9246 33320 9246 33320 0 _0261_
rlabel metal1 13248 34170 13248 34170 0 _0262_
rlabel metal2 18538 16830 18538 16830 0 _0263_
rlabel metal1 9430 30362 9430 30362 0 _0264_
rlabel metal2 4002 35190 4002 35190 0 _0265_
rlabel metal1 35282 36006 35282 36006 0 _0266_
rlabel metal1 34960 34170 34960 34170 0 _0267_
rlabel metal2 13110 19822 13110 19822 0 _0268_
rlabel metal1 12742 21930 12742 21930 0 _0269_
rlabel metal2 12098 35870 12098 35870 0 _0270_
rlabel metal2 11546 27608 11546 27608 0 _0271_
rlabel metal1 12696 30294 12696 30294 0 _0272_
rlabel metal2 12834 34782 12834 34782 0 _0273_
rlabel metal2 9982 30124 9982 30124 0 _0274_
rlabel metal1 9568 34986 9568 34986 0 _0275_
rlabel metal1 14214 36822 14214 36822 0 _0276_
rlabel metal2 12282 23970 12282 23970 0 _0277_
rlabel metal2 23598 15708 23598 15708 0 _0278_
rlabel metal1 31234 14824 31234 14824 0 _0279_
rlabel metal1 30820 14586 30820 14586 0 _0280_
rlabel metal1 18676 12886 18676 12886 0 _0281_
rlabel metal2 21298 15232 21298 15232 0 _0282_
rlabel metal1 29716 13362 29716 13362 0 _0283_
rlabel metal1 28060 13974 28060 13974 0 _0284_
rlabel metal2 25070 13838 25070 13838 0 _0285_
rlabel metal1 12006 32878 12006 32878 0 _0286_
rlabel metal1 8050 34646 8050 34646 0 _0287_
rlabel metal2 25070 33286 25070 33286 0 _0288_
rlabel metal2 33166 20774 33166 20774 0 _0289_
rlabel metal2 35098 12223 35098 12223 0 _0290_
rlabel metal2 10350 34340 10350 34340 0 _0291_
rlabel metal1 33074 15504 33074 15504 0 _0292_
rlabel metal1 31970 20808 31970 20808 0 _0293_
rlabel metal1 29808 11322 29808 11322 0 _0294_
rlabel metal1 29164 9690 29164 9690 0 _0295_
rlabel metal1 24104 6766 24104 6766 0 _0296_
rlabel metal1 30958 11322 30958 11322 0 _0297_
rlabel metal2 24978 9826 24978 9826 0 _0298_
rlabel metal1 26358 7378 26358 7378 0 _0299_
rlabel metal2 11178 19550 11178 19550 0 _0300_
rlabel metal1 9430 18394 9430 18394 0 _0301_
rlabel metal1 29026 13362 29026 13362 0 _0302_
rlabel metal1 23000 18394 23000 18394 0 _0303_
rlabel metal1 10580 20434 10580 20434 0 _0304_
rlabel metal2 22678 15946 22678 15946 0 _0305_
rlabel metal1 20378 9146 20378 9146 0 _0306_
rlabel metal1 15548 9418 15548 9418 0 _0307_
rlabel metal1 14628 13498 14628 13498 0 _0308_
rlabel metal2 21298 11356 21298 11356 0 _0309_
rlabel metal1 15686 10642 15686 10642 0 _0310_
rlabel metal1 22678 12818 22678 12818 0 _0311_
rlabel metal1 33810 15368 33810 15368 0 _0312_
rlabel metal2 34546 14484 34546 14484 0 _0313_
rlabel metal1 16606 15130 16606 15130 0 _0314_
rlabel metal1 29302 15130 29302 15130 0 _0315_
rlabel metal1 32660 14450 32660 14450 0 _0316_
rlabel metal1 13202 17544 13202 17544 0 _0317_
rlabel metal1 26542 13396 26542 13396 0 _0318_
rlabel metal1 19964 12682 19964 12682 0 _0319_
rlabel metal1 32085 14042 32085 14042 0 _0320_
rlabel metal1 29164 12818 29164 12818 0 _0321_
rlabel metal2 21022 16490 21022 16490 0 _0322_
rlabel metal1 31924 13362 31924 13362 0 _0323_
rlabel metal2 7038 27132 7038 27132 0 _0324_
rlabel metal1 5060 24650 5060 24650 0 _0325_
rlabel metal1 7176 27982 7176 27982 0 _0326_
rlabel metal1 8004 27506 8004 27506 0 _0327_
rlabel metal1 7314 24786 7314 24786 0 _0328_
rlabel metal1 7912 25262 7912 25262 0 _0329_
rlabel metal2 6670 20264 6670 20264 0 _0330_
rlabel metal2 4830 21828 4830 21828 0 _0331_
rlabel metal1 9338 11220 9338 11220 0 _0332_
rlabel metal2 9338 18088 9338 18088 0 _0333_
rlabel metal1 5198 24922 5198 24922 0 _0334_
rlabel metal2 8878 14076 8878 14076 0 _0335_
rlabel metal1 34040 11730 34040 11730 0 _0336_
rlabel metal2 28198 15402 28198 15402 0 _0337_
rlabel metal1 30038 11866 30038 11866 0 _0338_
rlabel metal1 29210 14586 29210 14586 0 _0339_
rlabel metal2 34914 13022 34914 13022 0 _0340_
rlabel metal2 20102 17374 20102 17374 0 _0341_
rlabel metal2 30222 15640 30222 15640 0 _0342_
rlabel metal2 20286 19584 20286 19584 0 _0343_
rlabel metal1 37536 9418 37536 9418 0 _0344_
rlabel metal1 32131 16150 32131 16150 0 _0345_
rlabel metal1 35190 11730 35190 11730 0 _0346_
rlabel metal2 11914 22848 11914 22848 0 _0347_
rlabel metal1 12926 9690 12926 9690 0 _0348_
rlabel metal1 24978 20842 24978 20842 0 _0349_
rlabel metal2 22678 10200 22678 10200 0 _0350_
rlabel metal1 10764 12886 10764 12886 0 _0351_
rlabel metal1 9890 25942 9890 25942 0 _0352_
rlabel metal1 23230 12886 23230 12886 0 _0353_
rlabel metal1 25070 15334 25070 15334 0 _0354_
rlabel metal1 14582 9010 14582 9010 0 _0355_
rlabel metal2 27646 15368 27646 15368 0 _0356_
rlabel metal1 17342 11798 17342 11798 0 _0357_
rlabel metal2 23506 10574 23506 10574 0 _0358_
rlabel metal3 1234 19108 1234 19108 0 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 1234 7548 1234 7548 0 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 5336 37230 5336 37230 0 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1234 5508 1234 5508 0 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 35466 1894 35466 1894 0 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal2 25806 1588 25806 1588 0 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal3 1234 22508 1234 22508 0 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal3 1234 6868 1234 6868 0 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal1 18170 37196 18170 37196 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 2898 38573 2898 38573 0 bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 12926 1588 12926 1588 0 ccff_head
rlabel metal2 29026 1520 29026 1520 0 ccff_tail
rlabel metal2 25806 38260 25806 38260 0 chanx_right_in[0]
rlabel metal1 6302 37230 6302 37230 0 chanx_right_in[10]
rlabel metal2 24518 1588 24518 1588 0 chanx_right_in[11]
rlabel metal1 8832 37230 8832 37230 0 chanx_right_in[12]
rlabel metal2 20010 1588 20010 1588 0 chanx_right_in[13]
rlabel metal3 1234 17068 1234 17068 0 chanx_right_in[14]
rlabel metal3 1740 2108 1740 2108 0 chanx_right_in[15]
rlabel metal1 28520 37230 28520 37230 0 chanx_right_in[16]
rlabel metal2 11638 1588 11638 1588 0 chanx_right_in[17]
rlabel metal2 38318 32215 38318 32215 0 chanx_right_in[18]
rlabel metal2 38318 27353 38318 27353 0 chanx_right_in[1]
rlabel metal2 9706 1588 9706 1588 0 chanx_right_in[2]
rlabel metal3 1786 748 1786 748 0 chanx_right_in[3]
rlabel metal2 38318 8687 38318 8687 0 chanx_right_in[4]
rlabel metal2 15180 37230 15180 37230 0 chanx_right_in[5]
rlabel metal2 38318 30447 38318 30447 0 chanx_right_in[6]
rlabel metal2 38318 28883 38318 28883 0 chanx_right_in[7]
rlabel metal1 33166 36788 33166 36788 0 chanx_right_in[8]
rlabel metal2 18078 1588 18078 1588 0 chanx_right_in[9]
rlabel metal1 36248 37094 36248 37094 0 chanx_right_out[0]
rlabel metal3 38740 12308 38740 12308 0 chanx_right_out[10]
rlabel metal2 33534 1520 33534 1520 0 chanx_right_out[11]
rlabel metal3 1234 30668 1234 30668 0 chanx_right_out[12]
rlabel metal3 1234 15708 1234 15708 0 chanx_right_out[13]
rlabel metal2 36846 2193 36846 2193 0 chanx_right_out[14]
rlabel metal1 20148 37094 20148 37094 0 chanx_right_out[15]
rlabel via2 38226 35445 38226 35445 0 chanx_right_out[16]
rlabel metal1 36110 2312 36110 2312 0 chanx_right_out[17]
rlabel metal1 19090 37094 19090 37094 0 chanx_right_out[18]
rlabel metal2 34178 1520 34178 1520 0 chanx_right_out[1]
rlabel metal2 30958 38328 30958 38328 0 chanx_right_out[2]
rlabel metal1 34822 37094 34822 37094 0 chanx_right_out[3]
rlabel metal1 36202 36278 36202 36278 0 chanx_right_out[4]
rlabel metal1 16192 37094 16192 37094 0 chanx_right_out[5]
rlabel metal2 38226 10863 38226 10863 0 chanx_right_out[6]
rlabel via2 38226 13685 38226 13685 0 chanx_right_out[7]
rlabel via2 38226 19125 38226 19125 0 chanx_right_out[8]
rlabel metal2 27738 1520 27738 1520 0 chanx_right_out[9]
rlabel metal2 36754 37825 36754 37825 0 chany_bottom_in[0]
rlabel metal2 37490 32793 37490 32793 0 chany_bottom_in[10]
rlabel metal1 24656 37230 24656 37230 0 chany_bottom_in[11]
rlabel metal2 12282 38226 12282 38226 0 chany_bottom_in[12]
rlabel metal2 38318 24021 38318 24021 0 chany_bottom_in[13]
rlabel metal1 8786 37298 8786 37298 0 chany_bottom_in[14]
rlabel metal1 11730 36822 11730 36822 0 chany_bottom_in[15]
rlabel metal1 22724 37230 22724 37230 0 chany_bottom_in[16]
rlabel metal2 10350 1588 10350 1588 0 chany_bottom_in[17]
rlabel metal2 2622 37988 2622 37988 0 chany_bottom_in[18]
rlabel via2 38134 15011 38134 15011 0 chany_bottom_in[1]
rlabel metal2 4048 36754 4048 36754 0 chany_bottom_in[2]
rlabel metal1 36938 3536 36938 3536 0 chany_bottom_in[3]
rlabel metal3 1234 14348 1234 14348 0 chany_bottom_in[4]
rlabel metal2 37490 7701 37490 7701 0 chany_bottom_in[5]
rlabel metal3 1142 28628 1142 28628 0 chany_bottom_in[6]
rlabel metal2 16790 1894 16790 1894 0 chany_bottom_in[7]
rlabel metal3 1188 21148 1188 21148 0 chany_bottom_in[8]
rlabel metal2 16146 1588 16146 1588 0 chany_bottom_in[9]
rlabel metal3 1234 24548 1234 24548 0 chany_bottom_out[0]
rlabel metal1 33212 37094 33212 37094 0 chany_bottom_out[10]
rlabel metal3 1234 32708 1234 32708 0 chany_bottom_out[11]
rlabel metal1 30452 2822 30452 2822 0 chany_bottom_out[12]
rlabel metal2 38226 25177 38226 25177 0 chany_bottom_out[13]
rlabel via2 38226 5525 38226 5525 0 chany_bottom_out[14]
rlabel metal1 26910 37094 26910 37094 0 chany_bottom_out[15]
rlabel metal1 38778 35258 38778 35258 0 chany_bottom_out[16]
rlabel metal1 37536 36890 37536 36890 0 chany_bottom_out[17]
rlabel metal2 690 1792 690 1792 0 chany_bottom_out[18]
rlabel metal2 5198 1520 5198 1520 0 chany_bottom_out[1]
rlabel metal2 38686 1792 38686 1792 0 chany_bottom_out[2]
rlabel metal3 1234 13668 1234 13668 0 chany_bottom_out[3]
rlabel via2 38226 21845 38226 21845 0 chany_bottom_out[4]
rlabel metal2 38226 15793 38226 15793 0 chany_bottom_out[5]
rlabel metal1 16928 37094 16928 37094 0 chany_bottom_out[6]
rlabel metal2 3266 1520 3266 1520 0 chany_bottom_out[7]
rlabel metal2 38226 3417 38226 3417 0 chany_bottom_out[8]
rlabel via2 38226 17051 38226 17051 0 chany_bottom_out[9]
rlabel metal3 1188 27268 1188 27268 0 chany_top_in[0]
rlabel metal1 2024 37298 2024 37298 0 chany_top_in[10]
rlabel metal3 1234 25908 1234 25908 0 chany_top_in[11]
rlabel metal3 1188 20468 1188 20468 0 chany_top_in[12]
rlabel metal2 3450 38369 3450 38369 0 chany_top_in[13]
rlabel metal1 38088 37298 38088 37298 0 chany_top_in[14]
rlabel metal2 8418 1588 8418 1588 0 chany_top_in[15]
rlabel metal3 1142 17748 1142 17748 0 chany_top_in[16]
rlabel metal2 23230 1588 23230 1588 0 chany_top_in[17]
rlabel metal2 37398 1894 37398 1894 0 chany_top_in[18]
rlabel metal1 14122 37230 14122 37230 0 chany_top_in[1]
rlabel metal2 30958 1588 30958 1588 0 chany_top_in[2]
rlabel metal2 3910 1894 3910 1894 0 chany_top_in[3]
rlabel metal2 14858 1588 14858 1588 0 chany_top_in[4]
rlabel metal2 37490 4369 37490 4369 0 chany_top_in[5]
rlabel metal2 38134 29427 38134 29427 0 chany_top_in[6]
rlabel metal1 34500 20910 34500 20910 0 chany_top_in[7]
rlabel metal2 32246 1588 32246 1588 0 chany_top_in[8]
rlabel metal3 1142 23868 1142 23868 0 chany_top_in[9]
rlabel via2 38226 10251 38226 10251 0 chany_top_out[0]
rlabel metal3 1234 32028 1234 32028 0 chany_top_out[10]
rlabel via2 38226 22491 38226 22491 0 chany_top_out[11]
rlabel metal2 38226 34221 38226 34221 0 chany_top_out[12]
rlabel metal2 36754 823 36754 823 0 chany_top_out[13]
rlabel metal2 38226 36057 38226 36057 0 chany_top_out[14]
rlabel metal3 1234 12308 1234 12308 0 chany_top_out[15]
rlabel metal3 1234 34068 1234 34068 0 chany_top_out[16]
rlabel metal3 1234 3468 1234 3468 0 chany_top_out[17]
rlabel metal2 46 1656 46 1656 0 chany_top_out[18]
rlabel metal3 1234 4148 1234 4148 0 chany_top_out[1]
rlabel metal2 2898 36499 2898 36499 0 chany_top_out[2]
rlabel metal1 10488 37094 10488 37094 0 chany_top_out[3]
rlabel metal1 23460 37094 23460 37094 0 chany_top_out[4]
rlabel metal3 1234 29308 1234 29308 0 chany_top_out[5]
rlabel metal2 6486 1520 6486 1520 0 chany_top_out[6]
rlabel metal2 1978 1520 1978 1520 0 chany_top_out[7]
rlabel metal3 1234 8908 1234 8908 0 chany_top_out[8]
rlabel metal2 21298 38158 21298 38158 0 chany_top_out[9]
rlabel metal1 32982 33524 32982 33524 0 clknet_0_prog_clk
rlabel metal2 18170 24990 18170 24990 0 clknet_4_0_0_prog_clk
rlabel metal1 32384 22610 32384 22610 0 clknet_4_10_0_prog_clk
rlabel metal1 34684 27438 34684 27438 0 clknet_4_11_0_prog_clk
rlabel metal1 31234 31790 31234 31790 0 clknet_4_12_0_prog_clk
rlabel metal2 27186 35632 27186 35632 0 clknet_4_13_0_prog_clk
rlabel metal2 32246 30226 32246 30226 0 clknet_4_14_0_prog_clk
rlabel metal1 33166 36652 33166 36652 0 clknet_4_15_0_prog_clk
rlabel metal2 17802 27744 17802 27744 0 clknet_4_1_0_prog_clk
rlabel metal2 19458 24480 19458 24480 0 clknet_4_2_0_prog_clk
rlabel metal1 18262 29070 18262 29070 0 clknet_4_3_0_prog_clk
rlabel metal1 16790 32402 16790 32402 0 clknet_4_4_0_prog_clk
rlabel metal2 16882 36176 16882 36176 0 clknet_4_5_0_prog_clk
rlabel metal2 20838 33116 20838 33116 0 clknet_4_6_0_prog_clk
rlabel metal2 19366 35360 19366 35360 0 clknet_4_7_0_prog_clk
rlabel metal1 25668 22066 25668 22066 0 clknet_4_8_0_prog_clk
rlabel metal1 26266 26418 26266 26418 0 clknet_4_9_0_prog_clk
rlabel metal1 19366 26758 19366 26758 0 mem_bottom_track_1.DFFR_0_.D
rlabel metal2 2346 34255 2346 34255 0 mem_bottom_track_1.DFFR_0_.Q
rlabel metal1 25024 18734 25024 18734 0 mem_bottom_track_1.DFFR_1_.Q
rlabel metal1 15824 33898 15824 33898 0 mem_bottom_track_1.DFFR_2_.Q
rlabel via2 17158 33813 17158 33813 0 mem_bottom_track_1.DFFR_3_.Q
rlabel metal1 20056 33626 20056 33626 0 mem_bottom_track_1.DFFR_4_.Q
rlabel metal1 18298 28934 18298 28934 0 mem_bottom_track_1.DFFR_5_.Q
rlabel metal2 20102 26792 20102 26792 0 mem_bottom_track_1.DFFR_6_.Q
rlabel metal1 19090 31246 19090 31246 0 mem_bottom_track_1.DFFR_7_.Q
rlabel metal2 33672 17476 33672 17476 0 mem_bottom_track_17.DFFR_0_.D
rlabel metal1 33580 19822 33580 19822 0 mem_bottom_track_17.DFFR_0_.Q
rlabel metal1 35374 24650 35374 24650 0 mem_bottom_track_17.DFFR_1_.Q
rlabel metal1 25668 32334 25668 32334 0 mem_bottom_track_17.DFFR_2_.Q
rlabel metal2 19182 20638 19182 20638 0 mem_bottom_track_17.DFFR_3_.Q
rlabel metal1 31280 21930 31280 21930 0 mem_bottom_track_17.DFFR_4_.Q
rlabel metal1 32844 21862 32844 21862 0 mem_bottom_track_17.DFFR_5_.Q
rlabel metal1 32982 14484 32982 14484 0 mem_bottom_track_17.DFFR_6_.Q
rlabel metal1 34500 23494 34500 23494 0 mem_bottom_track_17.DFFR_7_.Q
rlabel metal2 16514 28322 16514 28322 0 mem_bottom_track_25.DFFR_0_.Q
rlabel metal1 17158 28390 17158 28390 0 mem_bottom_track_25.DFFR_1_.Q
rlabel metal1 17657 23494 17657 23494 0 mem_bottom_track_25.DFFR_2_.Q
rlabel metal1 7958 20434 7958 20434 0 mem_bottom_track_25.DFFR_3_.Q
rlabel metal1 16330 19822 16330 19822 0 mem_bottom_track_25.DFFR_4_.Q
rlabel metal1 13984 20910 13984 20910 0 mem_bottom_track_25.DFFR_5_.Q
rlabel metal1 17020 24718 17020 24718 0 mem_bottom_track_25.DFFR_6_.Q
rlabel metal1 20378 16626 20378 16626 0 mem_bottom_track_25.DFFR_7_.Q
rlabel metal1 16882 11662 16882 11662 0 mem_bottom_track_33.DFFR_0_.Q
rlabel metal1 15640 13158 15640 13158 0 mem_bottom_track_33.DFFR_1_.Q
rlabel metal1 20010 22678 20010 22678 0 mem_bottom_track_33.DFFR_2_.Q
rlabel metal2 27324 19516 27324 19516 0 mem_bottom_track_33.DFFR_3_.Q
rlabel metal1 27278 21590 27278 21590 0 mem_bottom_track_33.DFFR_4_.Q
rlabel metal1 27048 14994 27048 14994 0 mem_bottom_track_9.DFFR_0_.Q
rlabel metal2 29164 19346 29164 19346 0 mem_bottom_track_9.DFFR_1_.Q
rlabel metal2 19274 16966 19274 16966 0 mem_bottom_track_9.DFFR_2_.Q
rlabel metal1 15594 19822 15594 19822 0 mem_bottom_track_9.DFFR_3_.Q
rlabel metal1 35236 21318 35236 21318 0 mem_bottom_track_9.DFFR_4_.Q
rlabel metal1 34500 20366 34500 20366 0 mem_bottom_track_9.DFFR_5_.Q
rlabel metal2 33304 19788 33304 19788 0 mem_bottom_track_9.DFFR_6_.Q
rlabel metal1 16652 31858 16652 31858 0 mem_right_track_0.DFFR_0_.D
rlabel metal1 18216 31926 18216 31926 0 mem_right_track_0.DFFR_0_.Q
rlabel metal1 20654 31858 20654 31858 0 mem_right_track_0.DFFR_1_.Q
rlabel metal2 21022 33907 21022 33907 0 mem_right_track_0.DFFR_2_.Q
rlabel metal1 15870 36142 15870 36142 0 mem_right_track_0.DFFR_3_.Q
rlabel metal1 33304 37162 33304 37162 0 mem_right_track_0.DFFR_4_.Q
rlabel metal1 34960 34986 34960 34986 0 mem_right_track_0.DFFR_5_.Q
rlabel metal1 32338 12172 32338 12172 0 mem_right_track_10.DFFR_0_.D
rlabel metal3 21367 21012 21367 21012 0 mem_right_track_10.DFFR_0_.Q
rlabel metal1 17894 21352 17894 21352 0 mem_right_track_10.DFFR_1_.Q
rlabel metal2 26634 14756 26634 14756 0 mem_right_track_12.DFFR_0_.Q
rlabel metal1 32798 11730 32798 11730 0 mem_right_track_12.DFFR_1_.Q
rlabel metal1 20378 19346 20378 19346 0 mem_right_track_14.DFFR_0_.Q
rlabel metal2 32246 11866 32246 11866 0 mem_right_track_14.DFFR_1_.Q
rlabel metal2 21482 24633 21482 24633 0 mem_right_track_16.DFFR_0_.Q
rlabel metal1 36938 10676 36938 10676 0 mem_right_track_16.DFFR_1_.Q
rlabel metal2 15870 10370 15870 10370 0 mem_right_track_18.DFFR_0_.Q
rlabel metal1 22034 11764 22034 11764 0 mem_right_track_18.DFFR_1_.Q
rlabel metal1 36938 34952 36938 34952 0 mem_right_track_2.DFFR_0_.Q
rlabel metal1 18906 13974 18906 13974 0 mem_right_track_2.DFFR_1_.Q
rlabel metal1 24702 16218 24702 16218 0 mem_right_track_2.DFFR_2_.Q
rlabel metal1 27048 21862 27048 21862 0 mem_right_track_2.DFFR_3_.Q
rlabel metal1 32614 15062 32614 15062 0 mem_right_track_2.DFFR_4_.Q
rlabel metal3 32407 17884 32407 17884 0 mem_right_track_2.DFFR_5_.Q
rlabel metal1 31786 15504 31786 15504 0 mem_right_track_20.DFFR_0_.Q
rlabel metal1 33948 25942 33948 25942 0 mem_right_track_20.DFFR_1_.Q
rlabel metal2 32338 13056 32338 13056 0 mem_right_track_22.DFFR_0_.Q
rlabel metal2 20102 22746 20102 22746 0 mem_right_track_22.DFFR_1_.Q
rlabel metal2 14858 27778 14858 27778 0 mem_right_track_24.DFFR_0_.Q
rlabel metal1 17986 27982 17986 27982 0 mem_right_track_24.DFFR_1_.Q
rlabel metal1 8004 11730 8004 11730 0 mem_right_track_26.DFFR_0_.Q
rlabel metal2 32338 32419 32338 32419 0 mem_right_track_4.DFFR_0_.Q
rlabel metal2 34086 32436 34086 32436 0 mem_right_track_4.DFFR_1_.Q
rlabel metal1 32653 34374 32653 34374 0 mem_right_track_4.DFFR_2_.Q
rlabel metal1 34270 36822 34270 36822 0 mem_right_track_4.DFFR_3_.Q
rlabel metal2 35926 36448 35926 36448 0 mem_right_track_4.DFFR_4_.Q
rlabel metal1 24794 32878 24794 32878 0 mem_right_track_4.DFFR_5_.Q
rlabel metal1 20930 34544 20930 34544 0 mem_right_track_6.DFFR_0_.Q
rlabel metal1 19918 34714 19918 34714 0 mem_right_track_6.DFFR_1_.Q
rlabel metal1 19826 34034 19826 34034 0 mem_right_track_6.DFFR_2_.Q
rlabel via1 19642 33915 19642 33915 0 mem_right_track_6.DFFR_3_.Q
rlabel metal2 16330 33745 16330 33745 0 mem_right_track_6.DFFR_4_.Q
rlabel metal2 21482 32368 21482 32368 0 mem_right_track_6.DFFR_5_.Q
rlabel metal1 30222 33422 30222 33422 0 mem_right_track_8.DFFR_0_.Q
rlabel metal1 25346 16592 25346 16592 0 mem_top_track_0.DFFR_0_.Q
rlabel metal1 31050 33490 31050 33490 0 mem_top_track_0.DFFR_1_.Q
rlabel metal1 32660 36006 32660 36006 0 mem_top_track_0.DFFR_2_.Q
rlabel metal1 34500 34986 34500 34986 0 mem_top_track_0.DFFR_3_.Q
rlabel metal1 35788 15538 35788 15538 0 mem_top_track_0.DFFR_4_.Q
rlabel metal1 35558 16082 35558 16082 0 mem_top_track_0.DFFR_5_.Q
rlabel metal2 32752 19142 32752 19142 0 mem_top_track_0.DFFR_6_.Q
rlabel metal3 34017 16524 34017 16524 0 mem_top_track_0.DFFR_7_.Q
rlabel metal2 13018 36380 13018 36380 0 mem_top_track_16.DFFR_0_.D
rlabel metal2 34178 17748 34178 17748 0 mem_top_track_16.DFFR_0_.Q
rlabel metal1 16790 33422 16790 33422 0 mem_top_track_16.DFFR_1_.Q
rlabel metal2 16238 36227 16238 36227 0 mem_top_track_16.DFFR_2_.Q
rlabel metal2 2346 35615 2346 35615 0 mem_top_track_16.DFFR_3_.Q
rlabel metal1 17204 32470 17204 32470 0 mem_top_track_16.DFFR_4_.Q
rlabel metal1 16744 30158 16744 30158 0 mem_top_track_16.DFFR_5_.Q
rlabel metal1 15594 26894 15594 26894 0 mem_top_track_16.DFFR_6_.Q
rlabel metal1 12466 20502 12466 20502 0 mem_top_track_16.DFFR_7_.Q
rlabel metal2 26174 15572 26174 15572 0 mem_top_track_24.DFFR_0_.Q
rlabel metal2 17802 10268 17802 10268 0 mem_top_track_24.DFFR_1_.Q
rlabel metal1 17710 17102 17710 17102 0 mem_top_track_24.DFFR_2_.Q
rlabel metal2 31648 19108 31648 19108 0 mem_top_track_24.DFFR_3_.Q
rlabel metal2 33166 22321 33166 22321 0 mem_top_track_24.DFFR_4_.Q
rlabel metal1 30084 19414 30084 19414 0 mem_top_track_24.DFFR_5_.Q
rlabel metal1 17204 17646 17204 17646 0 mem_top_track_32.DFFR_0_.Q
rlabel metal1 15272 30634 15272 30634 0 mem_top_track_32.DFFR_1_.Q
rlabel metal1 17112 31790 17112 31790 0 mem_top_track_32.DFFR_2_.Q
rlabel metal2 19642 35428 19642 35428 0 mem_top_track_32.DFFR_3_.Q
rlabel metal1 18032 36822 18032 36822 0 mem_top_track_32.DFFR_4_.Q
rlabel metal2 13570 28084 13570 28084 0 mem_top_track_8.DFFR_0_.Q
rlabel metal1 16698 26418 16698 26418 0 mem_top_track_8.DFFR_1_.Q
rlabel metal1 16468 11730 16468 11730 0 mem_top_track_8.DFFR_2_.Q
rlabel metal1 21850 19346 21850 19346 0 mem_top_track_8.DFFR_3_.Q
rlabel metal1 19826 34408 19826 34408 0 mem_top_track_8.DFFR_4_.Q
rlabel metal1 15042 31382 15042 31382 0 mem_top_track_8.DFFR_5_.Q
rlabel metal2 20286 34748 20286 34748 0 mem_top_track_8.DFFR_6_.Q
rlabel metal1 10212 24718 10212 24718 0 mux_bottom_track_1.INVTX1_0_.out
rlabel metal1 22724 17238 22724 17238 0 mux_bottom_track_1.INVTX1_1_.out
rlabel metal2 13478 19924 13478 19924 0 mux_bottom_track_1.INVTX1_2_.out
rlabel metal1 9062 10778 9062 10778 0 mux_bottom_track_1.INVTX1_3_.out
rlabel via2 1610 36227 1610 36227 0 mux_bottom_track_1.INVTX1_4_.out
rlabel metal2 27002 16507 27002 16507 0 mux_bottom_track_1.INVTX1_5_.out
rlabel metal2 27462 33762 27462 33762 0 mux_bottom_track_1.INVTX1_6_.out
rlabel metal1 11730 35598 11730 35598 0 mux_bottom_track_1.INVTX1_7_.out
rlabel metal1 5566 24106 5566 24106 0 mux_bottom_track_1.INVTX1_8_.out
rlabel metal2 20470 18632 20470 18632 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 12880 35598 12880 35598 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 12926 24650 12926 24650 0 mux_bottom_track_1.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 6762 24140 6762 24140 0 mux_bottom_track_1.out
rlabel metal2 32706 20434 32706 20434 0 mux_bottom_track_17.INVTX1_0_.out
rlabel metal1 20930 19890 20930 19890 0 mux_bottom_track_17.INVTX1_1_.out
rlabel via2 12558 21845 12558 21845 0 mux_bottom_track_17.INVTX1_2_.out
rlabel metal1 37904 16558 37904 16558 0 mux_bottom_track_17.INVTX1_3_.out
rlabel metal1 35328 17102 35328 17102 0 mux_bottom_track_17.INVTX1_4_.out
rlabel metal1 26174 16626 26174 16626 0 mux_bottom_track_17.INVTX1_5_.out
rlabel metal2 5106 33184 5106 33184 0 mux_bottom_track_17.INVTX1_6_.out
rlabel metal2 12282 21250 12282 21250 0 mux_bottom_track_17.INVTX1_7_.out
rlabel metal1 29992 5338 29992 5338 0 mux_bottom_track_17.INVTX1_8_.out
rlabel metal1 33534 21420 33534 21420 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel via1 34362 16507 34362 16507 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 35926 2992 35926 2992 0 mux_bottom_track_17.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 36018 3230 36018 3230 0 mux_bottom_track_17.out
rlabel metal1 14306 18700 14306 18700 0 mux_bottom_track_25.INVTX1_0_.out
rlabel metal2 12282 29631 12282 29631 0 mux_bottom_track_25.INVTX1_1_.out
rlabel metal1 10580 11322 10580 11322 0 mux_bottom_track_25.INVTX1_2_.out
rlabel metal2 8050 34782 8050 34782 0 mux_bottom_track_25.INVTX1_3_.out
rlabel metal1 9522 30804 9522 30804 0 mux_bottom_track_25.INVTX1_4_.out
rlabel metal1 8142 31416 8142 31416 0 mux_bottom_track_25.INVTX1_5_.out
rlabel metal1 7590 11186 7590 11186 0 mux_bottom_track_25.INVTX1_6_.out
rlabel metal2 8142 17238 8142 17238 0 mux_bottom_track_25.INVTX1_7_.out
rlabel metal1 9614 23154 9614 23154 0 mux_bottom_track_25.INVTX1_8_.out
rlabel metal2 13202 17102 13202 17102 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 9154 18190 9154 18190 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 18538 19414 18538 19414 0 mux_bottom_track_25.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 26358 5882 26358 5882 0 mux_bottom_track_25.out
rlabel metal2 25990 8432 25990 8432 0 mux_bottom_track_33.INVTX1_0_.out
rlabel metal2 23598 13498 23598 13498 0 mux_bottom_track_33.INVTX1_1_.out
rlabel metal2 27278 11118 27278 11118 0 mux_bottom_track_33.INVTX1_2_.out
rlabel metal1 18630 11254 18630 11254 0 mux_bottom_track_33.INVTX1_3_.out
rlabel metal2 10810 14076 10810 14076 0 mux_bottom_track_33.INVTX1_4_.out
rlabel metal1 9936 25806 9936 25806 0 mux_bottom_track_33.INVTX1_5_.out
rlabel metal1 10856 6834 10856 6834 0 mux_bottom_track_33.INVTX1_6_.out
rlabel metal2 14950 9928 14950 9928 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 24518 12886 24518 12886 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal2 18630 12070 18630 12070 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 35558 35666 35558 35666 0 mux_bottom_track_33.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 37582 35258 37582 35258 0 mux_bottom_track_33.out
rlabel metal2 24702 14858 24702 14858 0 mux_bottom_track_9.INVTX1_0_.out
rlabel metal1 29670 16014 29670 16014 0 mux_bottom_track_9.INVTX1_1_.out
rlabel metal1 28934 14960 28934 14960 0 mux_bottom_track_9.INVTX1_2_.out
rlabel metal1 15686 12410 15686 12410 0 mux_bottom_track_9.INVTX1_3_.out
rlabel metal1 34454 16456 34454 16456 0 mux_bottom_track_9.INVTX1_4_.out
rlabel metal1 12742 31926 12742 31926 0 mux_bottom_track_9.INVTX1_5_.out
rlabel metal2 12650 18666 12650 18666 0 mux_bottom_track_9.INVTX1_6_.out
rlabel metal1 9430 33286 9430 33286 0 mux_bottom_track_9.INVTX1_7_.out
rlabel metal1 36156 11866 36156 11866 0 mux_bottom_track_9.INVTX1_8_.out
rlabel metal1 19550 14314 19550 14314 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 13294 17969 13294 17969 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 35972 13838 35972 13838 0 mux_bottom_track_9.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 34776 18054 34776 18054 0 mux_bottom_track_9.out
rlabel metal1 13340 15130 13340 15130 0 mux_right_track_0.INVTX1_1_.out
rlabel metal2 17802 14926 17802 14926 0 mux_right_track_0.INVTX1_2_.out
rlabel metal1 36064 31994 36064 31994 0 mux_right_track_0.INVTX1_3_.out
rlabel metal1 13064 35666 13064 35666 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 36432 36142 36432 36142 0 mux_right_track_0.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 37260 36142 37260 36142 0 mux_right_track_0.out
rlabel metal1 29532 13226 29532 13226 0 mux_right_track_10.INVTX1_1_.out
rlabel metal1 10258 20468 10258 20468 0 mux_right_track_10.INVTX1_2_.out
rlabel metal2 23414 19537 23414 19537 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 12650 20332 12650 20332 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 14950 19210 14950 19210 0 mux_right_track_10.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal2 14582 34442 14582 34442 0 mux_right_track_10.out
rlabel metal1 21712 18802 21712 18802 0 mux_right_track_12.INVTX1_1_.out
rlabel metal1 29164 14994 29164 14994 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 34040 11594 34040 11594 0 mux_right_track_12.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35374 11118 35374 11118 0 mux_right_track_12.out
rlabel metal2 20010 16116 20010 16116 0 mux_right_track_14.INVTX1_1_.out
rlabel metal2 21390 17510 21390 17510 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 34086 12852 34086 12852 0 mux_right_track_14.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 35190 12614 35190 12614 0 mux_right_track_14.out
rlabel metal1 32430 15980 32430 15980 0 mux_right_track_16.INVTX1_1_.out
rlabel metal1 33718 16014 33718 16014 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 36754 15266 36754 15266 0 mux_right_track_16.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 36432 16218 36432 16218 0 mux_right_track_16.out
rlabel metal1 15134 14382 15134 14382 0 mux_right_track_18.INVTX1_2_.out
rlabel metal1 21252 11118 21252 11118 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 17894 9860 17894 9860 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 21022 10438 21022 10438 0 mux_right_track_18.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 22632 7854 22632 7854 0 mux_right_track_18.out
rlabel metal1 13938 8602 13938 8602 0 mux_right_track_2.INVTX1_1_.out
rlabel metal1 36455 12274 36455 12274 0 mux_right_track_2.INVTX1_3_.out
rlabel metal2 21574 14688 21574 14688 0 mux_right_track_2.INVTX1_4_.out
rlabel metal1 29578 14314 29578 14314 0 mux_right_track_2.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 19596 12750 19596 12750 0 mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 30958 14314 30958 14314 0 mux_right_track_2.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 30176 6290 30176 6290 0 mux_right_track_2.out
rlabel metal1 37398 12410 37398 12410 0 mux_right_track_20.INVTX1_2_.out
rlabel metal1 16330 15946 16330 15946 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 33718 14994 33718 14994 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 33718 15538 33718 15538 0 mux_right_track_20.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 35604 14586 35604 14586 0 mux_right_track_20.out
rlabel metal2 12466 16881 12466 16881 0 mux_right_track_22.INVTX1_2_.out
rlabel metal1 31372 13702 31372 13702 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 20930 13974 20930 13974 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 28244 12614 28244 12614 0 mux_right_track_22.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 32706 8942 32706 8942 0 mux_right_track_22.out
rlabel metal1 9476 35598 9476 35598 0 mux_right_track_24.INVTX1_1_.out
rlabel metal1 7682 27030 7682 27030 0 mux_right_track_24.INVTX1_2_.out
rlabel metal2 7958 27642 7958 27642 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal2 6026 25160 6026 25160 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 7222 27676 7222 27676 0 mux_right_track_24.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6900 28730 6900 28730 0 mux_right_track_24.out
rlabel metal1 16767 9486 16767 9486 0 mux_right_track_26.INVTX1_1_.out
rlabel metal1 3910 25330 3910 25330 0 mux_right_track_26.INVTX1_2_.out
rlabel metal1 9430 11322 9430 11322 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 5382 21862 5382 21862 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal1 8510 17714 8510 17714 0 mux_right_track_26.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 6762 16048 6762 16048 0 mux_right_track_26.out
rlabel metal2 34546 20910 34546 20910 0 mux_right_track_4.INVTX1_1_.out
rlabel metal1 13064 36210 13064 36210 0 mux_right_track_4.INVTX1_4_.out
rlabel via2 10166 35445 10166 35445 0 mux_right_track_4.mux_2level_tapbuf_basis_input2_mem2_0_out
rlabel metal1 31786 16660 31786 16660 0 mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel via2 32798 16507 32798 16507 0 mux_right_track_4.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal2 31510 35190 31510 35190 0 mux_right_track_4.out
rlabel metal1 8878 28594 8878 28594 0 mux_right_track_6.INVTX1_1_.out
rlabel metal1 8648 19686 8648 19686 0 mux_right_track_6.INVTX1_3_.out
rlabel metal1 11086 34986 11086 34986 0 mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 14076 34646 14076 34646 0 mux_right_track_6.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 23276 35122 23276 35122 0 mux_right_track_6.out
rlabel metal2 23414 6426 23414 6426 0 mux_right_track_8.INVTX1_1_.out
rlabel metal1 20746 16048 20746 16048 0 mux_right_track_8.INVTX1_2_.out
rlabel metal2 26634 9792 26634 9792 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_0_out
rlabel metal1 29716 10778 29716 10778 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_1_out
rlabel metal2 34730 12342 34730 12342 0 mux_right_track_8.mux_2level_tapbuf_basis_input2_mem1_2_out
rlabel metal1 38456 13498 38456 13498 0 mux_right_track_8.out
rlabel metal2 24702 11458 24702 11458 0 mux_top_track_0.INVTX1_0_.out
rlabel metal1 29670 35122 29670 35122 0 mux_top_track_0.INVTX1_1_.out
rlabel metal2 36110 17629 36110 17629 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal2 17066 19720 17066 19720 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 37674 11730 37674 11730 0 mux_top_track_0.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal1 37720 10030 37720 10030 0 mux_top_track_0.out
rlabel metal1 35052 16762 35052 16762 0 mux_top_track_16.INVTX1_0_.out
rlabel metal1 10212 35054 10212 35054 0 mux_top_track_16.INVTX1_1_.out
rlabel metal2 35926 17459 35926 17459 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 17388 35054 17388 35054 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 6210 10030 6210 10030 0 mux_top_track_16.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 2070 9724 2070 9724 0 mux_top_track_16.out
rlabel metal1 23966 8874 23966 8874 0 mux_top_track_24.INVTX1_0_.out
rlabel metal2 27738 8194 27738 8194 0 mux_top_track_24.INVTX1_1_.out
rlabel metal1 29302 16694 29302 16694 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 20976 11798 20976 11798 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 28428 16150 28428 16150 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal1 33028 18122 33028 18122 0 mux_top_track_24.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal1 37168 17238 37168 17238 0 mux_top_track_24.out
rlabel metal2 20930 35173 20930 35173 0 mux_top_track_32.INVTX1_0_.out
rlabel metal1 7590 18394 7590 18394 0 mux_top_track_32.INVTX1_1_.out
rlabel metal1 8326 20978 8326 20978 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_0_out
rlabel metal1 10258 22066 10258 22066 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_1_out
rlabel metal1 14996 15062 14996 15062 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_2_out
rlabel metal2 13202 33422 13202 33422 0 mux_top_track_32.mux_2level_tapbuf_basis_input3_mem3_3_out
rlabel metal2 5014 34748 5014 34748 0 mux_top_track_32.out
rlabel metal2 22310 11730 22310 11730 0 mux_top_track_8.INVTX1_0_.out
rlabel metal2 11178 32844 11178 32844 0 mux_top_track_8.INVTX1_1_.out
rlabel metal2 17250 14382 17250 14382 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_0_out
rlabel metal1 13294 19176 13294 19176 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_1_out
rlabel metal1 14306 36210 14306 36210 0 mux_top_track_8.mux_2level_tapbuf_basis_input4_mem4_2_out
rlabel metal2 8510 36550 8510 36550 0 mux_top_track_8.out
rlabel metal1 1610 19448 1610 19448 0 net1
rlabel metal1 9154 33456 9154 33456 0 net10
rlabel metal2 38042 10948 38042 10948 0 net100
rlabel metal1 36202 10778 36202 10778 0 net101
rlabel metal1 35696 16422 35696 16422 0 net102
rlabel metal1 25530 7718 25530 7718 0 net103
rlabel metal1 5290 23562 5290 23562 0 net104
rlabel metal1 33028 37230 33028 37230 0 net105
rlabel metal2 1610 33354 1610 33354 0 net106
rlabel metal1 29670 3026 29670 3026 0 net107
rlabel via2 21206 21131 21206 21131 0 net108
rlabel metal1 38042 5644 38042 5644 0 net109
rlabel metal1 19550 2584 19550 2584 0 net11
rlabel metal1 27324 37230 27324 37230 0 net110
rlabel metal1 38042 35088 38042 35088 0 net111
rlabel metal2 37536 32980 37536 32980 0 net112
rlabel metal1 1610 2992 1610 2992 0 net113
rlabel metal1 4692 2414 4692 2414 0 net114
rlabel metal1 38042 3060 38042 3060 0 net115
rlabel metal2 1610 13430 1610 13430 0 net116
rlabel metal1 36846 18122 36846 18122 0 net117
rlabel metal2 26910 14654 26910 14654 0 net118
rlabel metal2 18676 19142 18676 19142 0 net119
rlabel via2 6762 36125 6762 36125 0 net12
rlabel metal2 4002 6732 4002 6732 0 net120
rlabel metal1 38042 3468 38042 3468 0 net121
rlabel metal1 38042 17238 38042 17238 0 net122
rlabel metal1 38042 9996 38042 9996 0 net123
rlabel metal1 1840 32402 1840 32402 0 net124
rlabel metal1 37398 16422 37398 16422 0 net125
rlabel metal1 37996 34578 37996 34578 0 net126
rlabel metal1 21206 2414 21206 2414 0 net127
rlabel metal1 37950 36142 37950 36142 0 net128
rlabel metal1 1610 12852 1610 12852 0 net129
rlabel metal1 6624 37094 6624 37094 0 net13
rlabel metal1 1610 34612 1610 34612 0 net130
rlabel metal1 1748 3502 1748 3502 0 net131
rlabel metal1 2806 2448 2806 2448 0 net132
rlabel metal1 1932 4590 1932 4590 0 net133
rlabel metal1 1564 35666 1564 35666 0 net134
rlabel metal1 14674 36652 14674 36652 0 net135
rlabel via2 8050 36635 8050 36635 0 net136
rlabel metal1 1840 20570 1840 20570 0 net137
rlabel metal2 6578 4828 6578 4828 0 net138
rlabel metal1 2024 2414 2024 2414 0 net139
rlabel metal1 24656 2618 24656 2618 0 net14
rlabel metal2 1610 9146 1610 9146 0 net140
rlabel metal2 13294 33337 13294 33337 0 net141
rlabel metal2 37582 10030 37582 10030 0 net142
rlabel metal2 14490 35938 14490 35938 0 net143
rlabel metal1 8786 21454 8786 21454 0 net144
rlabel metal2 9246 25568 9246 25568 0 net145
rlabel metal2 36202 13022 36202 13022 0 net146
rlabel metal2 31326 11424 31326 11424 0 net147
rlabel metal1 21712 13838 21712 13838 0 net148
rlabel metal1 21712 8398 21712 8398 0 net149
rlabel metal2 9154 34442 9154 34442 0 net15
rlabel metal1 10258 18802 10258 18802 0 net150
rlabel metal1 35650 34646 35650 34646 0 net151
rlabel metal2 13110 35054 13110 35054 0 net152
rlabel metal2 30130 8738 30130 8738 0 net153
rlabel metal1 25806 32946 25806 32946 0 net154
rlabel metal2 28934 10812 28934 10812 0 net155
rlabel metal2 9614 19312 9614 19312 0 net156
rlabel metal2 15778 9860 15778 9860 0 net157
rlabel metal1 34730 14994 34730 14994 0 net158
rlabel metal2 20010 13600 20010 13600 0 net159
rlabel metal1 21390 2550 21390 2550 0 net16
rlabel metal1 5428 25874 5428 25874 0 net160
rlabel metal1 4554 22134 4554 22134 0 net161
rlabel metal2 34638 11866 34638 11866 0 net162
rlabel metal1 35190 12750 35190 12750 0 net163
rlabel metal1 36524 14314 36524 14314 0 net164
rlabel metal2 12466 9860 12466 9860 0 net165
rlabel metal2 9798 15980 9798 15980 0 net17
rlabel metal1 2898 3162 2898 3162 0 net18
rlabel metal1 28286 36152 28286 36152 0 net19
rlabel metal1 4830 8058 4830 8058 0 net2
rlabel metal1 12144 2618 12144 2618 0 net20
rlabel metal2 38134 32946 38134 32946 0 net21
rlabel metal1 38548 16626 38548 16626 0 net22
rlabel metal1 11224 2550 11224 2550 0 net23
rlabel metal1 6026 2890 6026 2890 0 net24
rlabel metal2 38134 9588 38134 9588 0 net25
rlabel metal1 14306 32402 14306 32402 0 net26
rlabel metal1 37490 18190 37490 18190 0 net27
rlabel metal1 37306 16694 37306 16694 0 net28
rlabel metal2 32430 36448 32430 36448 0 net29
rlabel metal1 5842 37094 5842 37094 0 net3
rlabel metal1 18262 11118 18262 11118 0 net30
rlabel metal1 36478 36550 36478 36550 0 net31
rlabel metal1 38272 32878 38272 32878 0 net32
rlabel metal1 24610 37128 24610 37128 0 net33
rlabel metal1 14122 11118 14122 11118 0 net34
rlabel metal1 38364 12206 38364 12206 0 net35
rlabel metal1 9016 19822 9016 19822 0 net36
rlabel metal2 32430 7956 32430 7956 0 net37
rlabel metal2 8832 19278 8832 19278 0 net38
rlabel metal2 8234 2822 8234 2822 0 net39
rlabel metal1 1564 5882 1564 5882 0 net4
rlabel metal2 2806 35258 2806 35258 0 net40
rlabel metal2 20194 15708 20194 15708 0 net41
rlabel metal1 12834 36822 12834 36822 0 net42
rlabel metal2 36754 3910 36754 3910 0 net43
rlabel metal1 1932 20434 1932 20434 0 net44
rlabel metal2 23230 7650 23230 7650 0 net45
rlabel metal1 2254 21522 2254 21522 0 net46
rlabel metal1 19481 2890 19481 2890 0 net47
rlabel metal1 13616 33490 13616 33490 0 net48
rlabel metal2 17618 14654 17618 14654 0 net49
rlabel metal2 36478 7446 36478 7446 0 net5
rlabel metal1 4508 12818 4508 12818 0 net50
rlabel metal1 2254 37230 2254 37230 0 net51
rlabel metal2 7590 27540 7590 27540 0 net52
rlabel metal1 20470 20910 20470 20910 0 net53
rlabel metal2 8050 20060 8050 20060 0 net54
rlabel metal1 37766 37196 37766 37196 0 net55
rlabel metal1 10810 2278 10810 2278 0 net56
rlabel metal1 4922 18190 4922 18190 0 net57
rlabel metal1 23506 2346 23506 2346 0 net58
rlabel metal2 30406 6460 30406 6460 0 net59
rlabel metal1 26772 2278 26772 2278 0 net6
rlabel metal1 18584 37366 18584 37366 0 net60
rlabel metal1 31464 12818 31464 12818 0 net61
rlabel metal1 4324 3162 4324 3162 0 net62
rlabel metal1 15962 2482 15962 2482 0 net63
rlabel metal2 37766 4896 37766 4896 0 net64
rlabel metal2 38226 28169 38226 28169 0 net65
rlabel metal2 34178 21318 34178 21318 0 net66
rlabel metal1 32338 2482 32338 2482 0 net67
rlabel metal1 2323 24242 2323 24242 0 net68
rlabel metal1 20056 14450 20056 14450 0 net69
rlabel metal2 7314 23460 7314 23460 0 net7
rlabel metal1 37950 7514 37950 7514 0 net70
rlabel metal2 6578 35462 6578 35462 0 net71
rlabel metal1 11316 11526 11316 11526 0 net72
rlabel metal1 7314 2516 7314 2516 0 net73
rlabel metal1 18285 10642 18285 10642 0 net74
rlabel metal1 22080 2618 22080 2618 0 net75
rlabel metal1 37904 16762 37904 16762 0 net76
rlabel metal1 22816 3162 22816 3162 0 net77
rlabel metal2 32338 35904 32338 35904 0 net78
rlabel metal2 28658 36057 28658 36057 0 net79
rlabel metal1 5382 7174 5382 7174 0 net8
rlabel metal2 6946 34578 6946 34578 0 net80
rlabel metal1 6026 36754 6026 36754 0 net81
rlabel metal1 27462 7854 27462 7854 0 net82
rlabel metal1 3128 10778 3128 10778 0 net83
rlabel metal3 30107 9860 30107 9860 0 net84
rlabel metal1 36800 36346 36800 36346 0 net85
rlabel metal1 37076 10234 37076 10234 0 net86
rlabel metal1 33212 8806 33212 8806 0 net87
rlabel metal2 4738 29988 4738 29988 0 net88
rlabel metal1 2185 16082 2185 16082 0 net89
rlabel metal2 14950 36992 14950 36992 0 net9
rlabel metal1 36662 2448 36662 2448 0 net90
rlabel metal1 19711 37230 19711 37230 0 net91
rlabel metal1 38226 35666 38226 35666 0 net92
rlabel metal2 35926 3162 35926 3162 0 net93
rlabel metal1 16790 36822 16790 36822 0 net94
rlabel metal1 34914 2380 34914 2380 0 net95
rlabel metal1 30912 35802 30912 35802 0 net96
rlabel metal2 33718 36720 33718 36720 0 net97
rlabel metal1 36846 36074 36846 36074 0 net98
rlabel metal1 14812 34170 14812 34170 0 net99
rlabel metal2 19366 1588 19366 1588 0 pReset
rlabel metal1 33810 29512 33810 29512 0 prog_clk
rlabel metal3 38786 6868 38786 6868 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal3 1050 36108 1050 36108 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal3 1188 10948 1188 10948 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 7130 1588 7130 1588 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 13570 1588 13570 1588 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 21298 1588 21298 1588 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 38318 26129 38318 26129 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 22724 3026 22724 3026 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 31418 36822 31418 36822 0 top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_
rlabel metal1 29118 36142 29118 36142 0 top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_
rlabel metal1 1564 35122 1564 35122 0 top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_
rlabel metal1 7268 37230 7268 37230 0 top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_
rlabel metal2 27094 1588 27094 1588 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_
rlabel metal3 1234 10268 1234 10268 0 top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
